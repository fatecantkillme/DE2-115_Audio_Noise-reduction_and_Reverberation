��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<��魁�7��4Ix`#=�*���8��svFƱ�U]aVF}�S&��Z7��bsPq���p�pay����J�b{#��])	��h��3Y�0,��U�~sIN��7d�Ywy����B^;V�NŒF��me��ñ�n&��{]�¾��p���b�7���𢕥q~ʡ2:�6xE8h�.��G��S��-��Y� ���/��*�C61��g8��ժ[�X�/�������������u�
l),AaP�
Kw�ˡ(@��W_���d������(̇ꏸ���6�7�4r����䎢߯T�V@����wR.�?��7�.Z����ls���Y�7�E[@��W�H�*$6�
X�g��#��.�;D���t�+�[�sz����� 3o�&��Yȃ5;F��������ċ����C��P��+�c��E(U�kF �?fs]�߸[��(8,��KW-�q��
?,a�����Y��������=���m9����9����?#�j{��4
�@ȵ�q ������т̵ �.-㯀S`2_��_O����H��'%�;�8�
�2��}	�gQd�f�x볗Md�Ф,�|ڷ�M�Ll�I�o��!<��p����������Z����<~���2�3�Uv�TX|�A�ˮR�r��k��xJ�W+���\��̀[�uȭ�L޾m��g.4�OQ��b;����S�W_��\�8P�����O�cc�\���;���Cޕ�s��f���Ʌ9���xs%Uw�jb��Ȩu�{�5[�t�Ҟ��&�Y0q�Ia�1�t�I���k���}R;�9�4��@Z��/~Z���7nfm�V*��Z6���jT0�Ԡ&}?�T��4���>��*���h�儘��d�
+/�W��g7[��>*���iv<��D-����l�z�N5��ŀC�|�`�)v�
�
�-*�O>��ɬح)Ac�p��w:�'렛�a�x�|V��<��ȉ��h���w�+w�99�w���B������օ3�!CH����Pf{�s��XA��ނ�j�a�n��{��ܤF�L��`�t$�&��vʽU��66��i�xDm~�V:o�,�2Ĺ�9�M���:�?�Zd(��+�=ź��p��Z4���Ny����MǦ���7���R����Im���{��)=e������S�<�)I��-��*��q�c���"���Q7R8T��c_XQ���>��W,`�O�&���L�%�o4.1��p�TKB�E���x���nu�����j�w~���n_	�P�����q����L�T�u�@�JGK�B+�%���1PI�^ʚGc���7���ޟ�(%|&�Ab����#� �jѫ)0��y����;3����Qw�e�Z��Lq����VUDJj^Q���fF&��U���B$�_���ֹjm�?����Ow�!���L󾠪�˾:}�u�-愞:�!�!�̰��_����k-�Yd(x�/G�S��W,��k,�w�������1`�|Qa��e�Il�s����	Mg�y9����3