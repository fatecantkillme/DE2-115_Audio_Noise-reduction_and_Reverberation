��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<ꊃ���7���+�q�j%�q�A������*h�x;&�ͺ|�Gqc���a���y�+�C4��@��Tռ�C���Et�̽]�_��K�bYo��N�!U��~c|(S酹ȺO!�m��p�����#k ��n�a�ݯ�~�1��h?���U6#�u�U%*E���zY��Z(BI"@���*�s+��ju�!MCzCq��"?,yl�YL4�~��s���&��_5�N�M�c�*�R�?�V����=��S0!}�Ĭ���y$�(���8�>���q�����M���1a��[ =���S��GT}xD�| �y{��il����^;K��H�m��V[��ߟ�-��e:^��O����9� E�ɛZ%BY�,{�:����Ѭβ_�4�C+O��x.�G@�=nZ���Ͼ� C[�8u�rm5��2R�81��:���I>l��x6l�4�vǡ8\?��� ���e���F�8��Py�ߊ|�^\�.B�_�6g�	e9��2�3��Nόz5t���Z��p��k#�%�{��YseTu#U^�|;���̚�G�J��u����aH��z7M�3�^�+#V7�<��3i��f�{w7~W���l?1/�Q��vY���RW��6��[W@�%�$���ȭ������s$լ�}L{���IPu�7�$-���q0�F�۴��:Sc��ַq	ط8�����d���I�{v��p3�ت@j�=D].���!�gi1C>�!�("�5)Zy��ʉ3�����
iE�jY�^�X�T}�@�ᶕ�#��OV��@T��Ƅ�S�8�?��T�w��DA&�Ҩ�X��ła���қ#�O��3�ty89��?�m���q���R��j�,�u�ҟ��Wm��8��;���4��Ꭼ2>$�`e�z�g�CѪ�.�]N���M�[{�q0�m��tK^�����,e���=з-�pmˬuS��
�H���l���\u�gǾ{ᕞ!����<� �1Ձ��9�mx��Jo̒�L�0�o~�Ɗ� �"���̉`P3;����+	擢�`���6n�،ԉ�A8��o�X�3�M���;M �P!yc��l����l���p�g�y����?�HU�ml�L+hj�9s��y�D%����A���I�h���Z��K\_���6�=����;G\4��c�B�9Q��ۻt��"�|<'W���<΄U�6BP@,�`���eLcSP7_�q��kDz�G��J��>��{����
���-.�����J5`<�2��2����I�s�H�땗��D����'��� i͖`<���(T������5��m�*����)�Z����?H�]�t�� �#��?�{����w��
�ȝê��^R��l�(z����v�o�dE���=N��HDE%�Nw|��f�1[0�����M����<�ʀ��������������j:/r�T4b�A�MB��iӠ��jH�Ǥ(K��B��H;7�5!d�V�Þt$�ϙ6�'@��>iU��证^���ռP3.�
�#1&�. O���5��K)8�ކ�r��E3�?N�C�ra�k�3���9���M��}�_����_�0��񛝭1=���ҡ����E(8
�xu��*K�h��X["�w�P���=�9������t^��� LTR>o���f��6a�޳�@�2�M�%p��cn���(}-a8�ߥ>����0w���<�t�$��Qn�A�X$eڍ��szs|!1��� Z���v�; f�@�#�d����2�$=�4t6�o�O�nj�n�r`�f��H�О���ѵ��KmC�(��n���n��4`���?t9�.�iѱnC6�_�UL�s��{�e�Ƥ�u��(�`�YM�|���	���|(��(�{K��L��L% �L�zJ�\��"z�\�a�khcq��{@3UGf,�6��Y�R���>��\I�pY���;��a�/L�&dH��{�+O�������Т���i�
�lQ���UB�6�����k�� W ���?	��	1x�s�N^{�E�����������?6R���9��m�v0	:�a�M�0�{
T]�� D��(����WWl�^��U����!L���q��۠��Xm���rHC)]fQy�9�o#T�G�b9{��oVYDb�����?cN
��;���{��BFW�Nc�
��;���XF:s%3�q܍�b�g@ni�U��6��@�1.��pL�J�?�-�����eJ��\ԫ�p�$��Q���M��[����:I~��,��wb���E%	��ħNw�M�'B�������P;��Q�Bw��5��W�'��-�g���� �VC��t��|���/7�d}I�5莆N�ݪ(ѩ8i��ѰeNR�%tF֚
�����b��)���N[>r��j3�~!nn���i���_D��;9��-˙��ɑ�,�����!�B�8�A�d��b����%ao�UX ��tǍ�aM^���+��"�'N�[C��x�˙��f_V�L�J�N��@��d���ƥC���O����"���V am�Yx)��$�.�m�D Ku���?E���f�֧$����IP�퉞*��h��I�)C}ˁ.�����Z����kB��6Ͷ�U����*�j�P���� ������X�Dg����aiʥڟ�ܖ�!�q�uD_8Ԫ�BO��5�f�ο��Ǧ�F�� �k�*祲mY���ϣ'��ګ po-��)���S�	��T�t_��Z?H$:mm��U�U����ԅ��Z�� ��F�~#t��B���!n'�i��샱�iS��1E(4������q,��Lq��ٳ�V�z}@r��aq��6�50��y�2�������H�cN���8���/~�`��1W���m��$�J���ʹ�!�vT�4po
���s2�&�ٍ�K��IU��#/"�����6Q�~�f��
p*�t7�T�G�!Wˣi;]:$"�f@�]���y��FBؗ��*�?��jl���E�t���󕔶��@��u�i��s5kr��VM�8|�S2�y�J�q{��۴��ޢU�]�s����vc�)m�M��"���Ǫ;4B4��BhW�;�	�!�J�&��h��M�	S��[~�?v�O1�M�і'!�I�/{�woL���e�1�<�F|��0X�P���F$L#��6<Ƒ����y�.%P����S����5;�i�d3���D�E ȥ9 Gݖ>�z��c��,.K��^`,�*fo�{w6s%w����cV.���ۘ�t%�x1�{oz ��߼�rh�BL|����OM#��14I}�P=ʼ�ie/�e�W�{��@���0`>�� �l�/� f*��E����r
@=֍]��Gg�7^�"G`�[-v�a&ߋ{�3H��[���:�����P	gZWl�3�j�k�e��Xș�	K9=nk���	����^�x������e�r��5c8�������_s�|e2ܫс��Ǳ4
��L����>�ގ�#ǿT�݃ZV��#��T�ç��t�� �I����}��� w��4��Ҥ���m4���PCB�:��e�]�~ľP�;m���x��{ƕ
��U�>+~��x
h0Ϙ3��8�sL�װKM;!�L� �-��gY�����𯚁oP˴��ʁ��F�d-x_'#r�:vy<Ϭ�O��ܬ�����/�*P�1t�_>���Q�P�*q�N����ŷ�aڵ���D� ��6oG6T\Gj�X�͞^�"\�|ʝ�sz���M=�f��S�9;�Wz��_��N���N��E���t|"HF��R�"��S�z��9��5�tu<��#� �Xؕ6(~<�'7�{�`�����ڼ�KWٗ���ߌK�I���Hgh����56VY�c�?^T�v���� �dW��$?��"�?�Zt��q�[wc��LPX~"pp�\�N��v-�eZ���6Ϯ��B���?ŜWa�5�
6]��Od���B�\�����6 u}Bb��'���=1�<���^]̇���ϛj/� {�!��lqWj5i�vٕZ�f�뉑�՜������Q�WA{�D��)I�G�j����ö�\��y!�k�4]�[��P;�a���y����ތ�b����49cM�P���2_��G��"^���v"B@=�9�ɢ%g��C�ĉ
'm9��U�c��}���m5m�_G�?Y����Ty��F��u\4�ߑ�V������^�|Q:� s��� ��',UB�{pCf�rg"N��y� �7�J�< &�I���f������N_��ޟv0!�Nk��'�����YD�����q𽴑D�,�sy�$�fJI��f����9IkF��x,O'�؞�� )��)8�t6;Nk���x���R�����b+a������/Ƴ(l�,*����"/mڮ��Vh�Bge��ԧ��е�2	��-O{�ܽ󭠏 3)mz�!����!��u!�:���L*�I���	��;*�u/�fԤĢ�$Fz"~(dL���q�����78/ݐ��o��v}~��Ϻc�ˋ��!�1�Z� >Bٴ.~y�槵�e3�;K��be:2�����f��Q�b���5����Uh�3�3Z�Q�1,\�\���6n �� �7сd\,D��<�-�1d(� ��<�zt��(ˣƳO����Vm�&Sd��D�u�+tHftWLل����p���i��Zw�O4e�Ƕ�y���*�[��z�n/o��o&� ]U�AcE�v�Q4=-�'Y��aM�iS�8Â����t��6�q��)Tvh�IQ-��y��!��;��5U�E�� ���w�ۺf�� ��Sv�/S�&������!P��&��3U��z�J���Ip�\/1��B�1�����a�Ls�V�M��e�51F�̭�i�S��>-ܭ{�g��eۜ7*X��q
N���Ţ�IaO��b�N�d@���oh�P\>�T>b�L�y��r�&!�[�����{5�.�!�H49��i���>�Y���2�����c�1;�&���X(O�XW�[���Ci(���nqٓ�1<�]4�.���H2�5cҢ�S8����L��P��0R���y��&������������^��WJfoSN��/DU�Id�ǋg�3�����{/I�ߒ�lGyl����T��X��l��ۚ|����B-˓� � �73r�O���H�f�$�'�:/���&E=U���J������+A�2n
���:j��R�1��,��:bM�������I0us����j��m�Fu",L�[lW�l�f�_v�hZ��$O���w4�a�<�8|�Yy[�J�����K���u����?r4�ޖ��x��s�t��cf0� `�����e�<$��(Cz�X��EO��+&�|-~��$)��s@瓎�8����ɀ����#r+��=eᖚ�$
Y�ȯ��̪���z��-�������/�wɨ�u6�H�`�������n�n��w�M��yd�uD'������]��3��'�-��Ǌ�f*�V|�wU�s�
m�kqm�3>B�3VmO��i���VqP�}0� )��]�z��Û�$�.�3GN� GH�*?�ʯ�pK�{]�?�?��P����M2���ToP1�@��j3\�>a���~a�����	��H-�����xDϜ�69�/TٗJ���l�؂J(xӋK�k�sZ�~&���d��~�z�"/̔I�	��ڴ	�}�T��h?1�s�X
" 9��F6��~ȠL:���Q�,�-I�{1�I��
�r[�C8`E fj�K�^HR�ݹP��á�e�6���� �:��O@�Q��C�Hc��0s!���Q�k5�2�D�:šUK�*�a�/em��*�k��<<�]�u�����$��-��bk�u� �?2����	�J4�H�N��c�L?� ܚ�9d�C�t���O,������(˴ly��;��j�ܾ!�� �e�w�3�%�#^t�"�S|[�#b���Ŵ6��?l�dm�ɟ���9��h�~���P�/�`��b�|�ic���I������)J'L�-�Z��-�^#����K�.POGp���Ϳ+�~H��(�t���!'�������,ġS�t���ʾ�V���Q,�c�bt;��XG�3a���dq�!�tR��̫�0+a�¾�\��a��3.�6�,�s���I��(���	d�qcG"oӘ�g����`4�4�+�^\XE�ග��?�9|ZϜ���&�C�lO�U�����.���ч)!x(c���������>tru�3�!]�[�Y(���r���5bN���u������n�oc��[E���i�=c1ٯ��ŕ�%o*�=���Xd�h@{MP$��*疎��c�֬Z��O�Ut�e7�����b��)�fZ:��U�
N�j7�:��^�RW��2´S���n��t.@�-���ز-�4���l~�W�e]�vJ5�S����H����?��+���� �I�?*F!�˛RU�.����tF7~�F�����;��"��"і2��EuT�CB�>w�*�hi��VC�Y:�^X�ד�]�~7�~>�z]K�`�|j�>o�B�h��9'�;hDJ���&Z�,�s�h�"�I�O�ƴF�ׯBߢVK�m�w��YKb��bH����K.)�"5H@J�3O��D��i(ǋ��Q(r���Z������ɛ+b���X�
<��A�ݫ�ٸ�o�W��t(
�˧B���a%�e�����7�ӏ?�3a��گ��ʦj��Jʊ����K������72��M� ���9(��W78�=N���Mc@��V]�23��v��!O�O���d��w)�z��,�NN|O�H���gLA\���(ۯ�_qUkA��*"Ё7K�ĽJ:����o���;�����@q�(�z����yl�xݰ�|�b����8R+��A�}(�C�b��"Ed�<V�R���ߠ�B�M�\$�_�	��Qsa�����ŔMKG+g��	�U��K�\F=9ǵA���ͨ6�� �V�_����ӽ�^42��-|��Ih����L� B�쟜|:��*4��,�7�C�)/�S��h���DNV�gR&k.E5��a�O0��]w����X�����y��·��1���ݦs�=�6�Jeϊ+� �w��`B��W&�\LD��e>�|�F��/d�an��]v��+c�@Fv��sW���.�ZS���cz�~"i��L��"]�j�C'�Ɠ�u�]�#FV��	�����HrV�ۂ�օ8G"�h!�3�ũ��@F.�q2 ��Rқ�8%^<�5B�U(���כ3����Zjm��v����RP*�i�3S��7~ٜX��ac���^���v�6d����n������vx~.n��,�Z�E����)�0f�ǕO�8dNM����8�=�c/*�V�.&H\���[Bl�|��U���J{^Rص��� ��Ք�tG��;cD��eNDǬ��g<v���A�<w�ν`J�L��+XA��<Oʵa��"�o���ti'2�PF,�I��X�<�I�[�mq��Ciy�Ef���ȣ�WXUG�/X5�R��0����(߉-�Gv�����j��
8r��-4��a]irG�ҍgŀ
����	�?U�����$L9ͅ�:n��}S��4�p1�m���U�?z���V��*�W��'4���t4�ESWU}��/KB������bt��ī��PN��]�_S�ZR�} ��*W�.PLAȇ�ǂ�k�*���å�u�jCō����}������۫��*j��$�4Q��wCGb�S���s��o顥;�C�,ԍ��+�0��h�bL.���r������̧]��hVZȱO��|v�� �^6ў�[W]�a�y��Z	��]_qW���(�6Wш��}Dv8KZ��Jv%�Ӻ_��[� b��,���- ���P�3Z���8�T���!����8�o�Gڽ˽�Yw�9��1W8�\F+�+��H���8��F����/9U G�}zqQ���P7��&`���q�4��)� &Xr2��5��rҐ��p7��xx���Qy�|sc�����������)Q=Lހ�TQ)#[���E�ke1-��ب�7�����41�vi�X5��a@̳�Y��r�T�9c|3$�G�/̡���pRld^3�,�u�8�0�_Sb��э ?:\����iC6aL�Gj_���ߧ]7�\��49�5�O
�C�,|��BD�e�쵁|�ǈ�eS�d��Oz~���ͪ��i[5�]���Sq�sy1��6�I@vC��h����*��*�WB�h���W����"HG!+ڸ��Skl�c�l���U#�Ɩ����RI��m��!x=�~:�Z5'K�w����ސ��!x�fߞ����ᶛ��h��'�
�B?�'r�g�;��o��T.��_w�Uj'��g؞�iFS[�;<��������57��5^8\��&����1g�k�N�)Ւ�X�Cd1%QN_�%�a���^�CĐq���ܰOKl��,Y��?�1��@��9���cbzK+�ޙ\"Q�M�t[�{�O���'�t(�`�!���뺑��{ё(����mHo�-��E�I'��& ��
^:��������ο�'}����p�9�O*���֝P�h�B�qob��|�-5�՜ۿ���^��*�1��&� G�8�p������?�7��T�2ytr���@��-k��� b�.�w$���b���Ȳ;#S��)'�Ϩ�n��M`"�a�r5?P\L��T�OC�������ar����ԥ�Ls�tD��I�}8"�/��jϗIMVQT�M��Қ�iؕ�/W��_zU�?A����_s��c͵=�q��#�tzB�_�[�0�����b��+6W��0R
�a��I�u�ւ<x�U�8Jq�G�3��+��b�#ܨ�}��rV�j��yjyĒ`3�p\Y����S ��q�"< T
[:�	}H�����O(Ũ&����&������n�.��"ֈ��`PV^�m�$�jo�����²��d��O��*��1��iG�Y-����XuZ�i
g7�	�-S�,������X�[`߄G�/���s�7t�S����`��M���)~Z����}����2�TWu\yo�r�=�H����n,�u�l�xa}{��gA��d2m�QӜ�����Н�q��k���-��T4��������Li��6����v���"Q�e\�^�M�iŖ <���4�a�K?s��sתq�>'����5��Ggi�G�����CQ���K��Eۄ
Ѯ�N�����e+/���A2��H��m�A��X�Q���ju˜l��Lܓ���Ԏ�3�ԅj���h��dAQ�V�ߧ�I�k�����T��/� �w�)�9��Y�)-1�g����~F&���\ O�4����R������}����φ����t�����"|"�����E�=�_�C�®Э�\�h�:���&q�uf����8P޵W)K6�,?ں���ւ{�UB��q*�cg�
��]J�P�2C���I5��y���J�� Q`��K�e�J��s��VZ�w��/1�K�+��o�ܠ�['WnT��1�tV�.\5�$��)�#n��f=��ɔ�8�>([E2� �C,����N�u��s母�5	���
i}ܡ�%���ɶ���I�b|����H��bj�$,�!	��!�w``a����?eJ����2k����f����}W64RC;���T�L#q�}$O���5,�Y���T�A���1n��'1>,����T�a�Œ�ꈆ�鿙��F��5��@�BY[0��SxKW[^�f�^����������O�]0���L�t6O���o����2�4��y�v/�#���iT�sj�K{0LŗOvK��(��Ԛ��?��׳�ט���ҫ�\G���Ɨ�w�>&<~K�&�ږ�;�)˹��^��A��Co�yC�M�����-�W���9�}�w��{%��`B��$�Y��5�Ǿ�#N�`���aO�_���� �/����i{'�N��C�h(ۂv����p)���"_ծo�B`M*p�
ӏ4U�N��4lC�R�ھ���]��詶5��Xl�i�G0� ��~�|O'8��4��wh�T�A^�pm��»�n0��;�����U1e.o�֞� NR��ԧ�� ,-U�<��5)рV�*�9��P��dE��R��E����6�&2 ��}���\�4{��͖�b��V��B}XD��������P�
gή�*3��2�3�J�P���$���(m�}��͞PK�<�@		G�k�
�
�!�r�]=�H��y�T�ou�vy ����6-�%��sf��o���S��.���N�&U*I��KS�X��[hh����I�Ǽ�aA�r�R�{j�a�{(hpy:\�:t����S�s��' �L�\O���i�WL�xn2��:"�0�I�dbz1�gfũ�&�'��' ��iN(���p2��6jٴ����N},g���"; �By����!�����z����"� �������[��"������w�-3a��_�n�*��v�������ӆ��n[둂�'�>^���~aĊ:n�1��G%I���
��*���e���O�P����W�����5��.
�hG�ڱ�_��rd�|�3�eT���%_C_���F�_�n__(��>{�]�	Y�س8X���TS����@c�kuZ��}��>K����C��q��~��!�e�N���,4��[��5��H�����L�j��e�4H+:�?�:��Cᣝ"����`Hm<gU�~��b�Abw]L��Y���y(ޟ��#T�J)��K�=Ę��_h�-���6�(�-������A#*|�E�,%���-YNr*'�H\#�����[l��>E �	���r�\S�7t�p�^ڭsDz"��v&��:$�rp��
7�[+���//��Q�R�WI#3M���s>Dۉ w�4XT��$�ц��A!�y��-���;���!uiʺ����]���(����'�tX$����(�e�*�fI�-�%��k���N�c6Y�'�vg�g_m���(���/�;/:������o���#%Wr����f��G��Ņ�������5��B���]%��l�g��hX���i�}̢&n�Cl�����坻\�TF��SM���a.��*��-1N=���>�Կʚ�A�Jjtz)P1�Tn��Jb��hB-�����>k7�\�d�����9�&(�B�cQ5j���ѦopV^�X�0���[����s�����;�K��8/X��e��T/ZƸ�]t��Ȳ���Ln�:����2��m���41���J��y0=E��? ���c=���d��n�����_�n�3Tڼ�겡?q.��-����K���b啋й&�������XS����cD�*w͞"�m�t*�"