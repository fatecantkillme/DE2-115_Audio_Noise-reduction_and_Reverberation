��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�8k�)9�k���J�f ۘEN�R��>�Ug:�&�1�a4ⳉ=���Hpsx��I̡����3������u��,���=�
�D�ܱ|��+)��5��Nm��ݕ�9#���|�Q�����J��E<v�)q��yGV��c� �nVA"��B3����%��ـ/3�������` �hH�T����(�+��t��M��hP5;�R#	��$�����.;��
�q]ue4�K���rC@�*Mn�຀��y�A�h���M�l��}IS��вw�̬!�*߸!(1��X%W�)��xc��Ql�nR��s_2�'e鏑�5-�!������e���a�Q2	���<�6�_��_��$*��"��V1�l�k��L�����g
���isI�D�jv��s)��C��;I˝+��F��%�Nl� �i�a�	��&���DkL�>��T���U&ꮳf{�"������`Ǯ�ӭ�B�(H=�7U�@p
Y����������7g�LWar�2��ft�F舫E,>f�� 5�w��(�v��Z"tB�l�͋8�,ζ+T1�k�oN�ئ�p�!��m	���֢���;�t"�J��$=HXAE|��t@<{��y��N���'G�p���	�Y��,p�._�|�`�7b~� ���C�����:�Q�����G!,W�=.�<�7���ǉ����G��j��=��Pf��;��T�����9�J��9��I�!		�\t�|[]$��Z���ٵ��c�YAT�>sͯB8���{�G�JLg�Z��7�Q��a��	3�jƭ+;51�PݶNy�Ӕ;
�})8F���b��b�9�����RA�\h��$5F���!��9�`��R��yz�EÇ1�s����73���u��_t7'�8,��Q+N�g;�s���njZl��01�;W&�#r@���AJE�I2�v�����C��_e~�[�TFA�������.�_4�_�����x�	��;��C�eb��>��?9:����w7!n¼ρ::ArR� �s�6�-ƍ ���D�	%�]XWu6ioȾh�q�3S>@d�y���_Z
��̈���mJ��w��E�k��A���A�RL�G�QC�·��3���c����"_����]^�9ӷο�a2�q�A�]���M�{�䬠�W�?��u�?p�w��V���%5H&Z#�e���UH����X��u��5����l�Ml�[�x2)�3�������!���Y=Է-�Y���X�D�Vג�I.�D����]*,R�^ؑa����n��Z̯�f���F~i�x��x��\�,������"�>.,n)��Q�����M+2ÆaO���v����zf�±���{Zn�v7H;� vOM~po��
�k�����D*��-1�S>��\@M��ϜwrP`3Dt]^�[� �v��/��Oǌu?͔6#2?�k���uxQxJ��/jH�2�X�.�3���(2xZ��f��aJ�=P=жӽ�g�q�ޭ���[�����z�p���PL����&U�/H����ϋ-M�-�����t~�~�|`8����c��+&���à[�wm�vۻ\Q��X���%�q;z&!����#�2�sl����(���:ʪ����t��P�/���ʈ6�����)4�@@�e�����A�@�LK����8	l���&i~�<m5��u�V��af�(S��8 -�ֲ�g�b@ �<z4��q�*|O��v��y��^��Y�p�"���8�!k#1�h&:�D��N_*udO�� �F���.���#���{�����֋`a*��j��C����3Ѱ
3E@�տb+tW���)Mo� �e�T���< ���t.�DO:%���m+�Ǎ�=ip��^u����<�^"�[�|�}m�,T���v����P���@*:�_�?��~��ۏܥ����_kug.��fT��E�AN�%���a�=u���ZE�ĥ�h�mW�	k;<�k�GA)��~��RA�J��yK�RO�PI?�J
��� ��y���V�u2���s3n���3�}˔��2|�hd1FWQ`�My����PRa��#�����#$���Za�f�X-ܸY�!��Tͬӕ�0�m`P�Bk��7��+gc�Ä�s#��)/in�����R�*ou�|NTB���q~��:1�,��40 $�k�l$�[�'��{�����	"/�0̤�v��@�R�`���q�;����d���o��5:v�����ɒ/�_,֖.��bK6�Z2TI�H[��=i����W�����O���6=��|��,Uy�*��b�ز�$TF��m9�|�^S2�N}p�-<�@����@������]}��8KU5$k�_�E{�� ���auz�7�Yd��j��~�G�7;X�������Y/�3`�}����z%yP��5��j'��fM*������y�2�g$ӕ�0�9P� �!8ݑ��	z%�m/l�� n��1���dI:����p�4R���2V���ϣ&5X� M�N��Sd8�:7{cP p��W��Q�.&�0!�^W댑�6�}F�`��x�L��K[4s���1�ꭁ��ug�a,݁����z^
,.��J����*�$
Q#����(0i/��C��Tl�gw��9\�+[rn�a6�i�[��/rDӽ̢tY�B-ܒ�N�A��{��&l5G!��C@��o�N�	h'!n:�����=
�*��o@D� -x�m����@�mpT]�΃�����Ｄ��?%��m�Q��q��ϲ*d��*A����Jegy#����D9B�&(A���1�dz�p�����9H�����zFzo��Ѐ�{�_q�-�j$�_�{��ݪ�7�=l����J��WR'�	�����iGR������&��M[�[��oG���Rb�t�ؤk%mu䞭M�b��6&���aMz�����@[V�5��
���6ӡu2�+�u۫O��XYX�J���}FV�D5���]2�&W�+U�/�}q���W¥�zU�Ȉ�%��Ő����R���/�@�"����LP�����vMҡ$��X#�y������j]$@�}2:Y,��ε�ަ�_�^⬢�zlJtW�0+��sr�g��=�E�
P�?]d����wd��<WLU;{č��?���.zG鮟��z ��S�{�C������6x9+����Ic��	,���uSx�]�-U=����u�+�S ��H��T
/�w�I���P����?�5D�C�rê��L��su���8���[��Y�)/~��gE�����j�@�n��Ƣv"	g�

�[����мRr�=�&��;�	~E.WB@��Ԋ4��[;������	 A��*1n��������
w!--��co���d���w	[6��é�2�~.H[�[F��7ŎN1����E�w�o�;l^�Хp@!��T���>իx1���J1ۛ�h�)��K���%4�ۙOv��ʰ$λ�]�8���BPW���!���\�3�=H	�ΏBON��c�*������^x��5=a�o�*X_&�$�.�mA��m�rk"Y��С'��xb��u�35 ߖps#�0-��֬�홰���'b�S�ޔ>�BMa^����@h��I_�pO���C�[s�ߚ�&1�L|+8����Ey���R��@W�b,DF?��X~�ʊ;N�)��l>�HbE%�uR��ᄣ�y�@bZ�"H�ʩ���룎��dA;�
9�r�|��߲�Xki��4�I��YJd�'�5J�f�U��fw�:T����cH�� �B��z_\G8x�$)����`�U���ER`#dL	b���%�ߤ �>��,�B��8�B��]�;$��3��!_���r��S�U7f�Z�q�hQXc=���2��v�j����;�J
�[	� +�5N壸Y]���b�ڬ�L��@�[!K-���9� �wH�/�m]?��o������u(l5eF���dC����/����&%���|�-��ˎE�K��,�N��[s����I��ξs�o��Z&�h���>nt�v{�"�]����hf'�C�	ѣ���[̄W�.��,�d��G��#G�Jz���l3���b�g��f�!��?���`jȟn�BR�=�s�5�k��&'e�녨��?P�n���M�y�Q��Ĳ����q�-_"�VߎS�|?y��u��P:}�ĉA���`��%�)n�ۅ�X b���d��rЍ�cN}����U�7V�	�ٞ��T�����B�����������o<�2�(�,�ї'�*����F����h���d� }�a�s68���ޠn�I�\���c��Xl��閨/�\��[֌���̽a�*[��i������U�����x<H4��a���C�g-%���j|���.��P�+��%3�qZ�Vv+1�P�7?"�����ɗus���q�$x���`�m���?���?�,�4)�5���6����_#���Z��F��aǀ�%Tsv���g[�(ZiylJw�)�5��MtR�E�Eiy�?[����dw퐿����m���I&�zM��c
��Ԙ�ڷ����P�	���y���s�����}u%���fj�c�g�v�%�@b��ϯ��}��]؄�ɧ�H��&QSע@�u�y�P��9��؅��vBF �n�0�Qq8��ml�zP�~IbKd���X�T�����ڪ��vȉ�u`钜��,�5m'x��MW��$�/��n{/��<_yV�0���
a��+?��@�$��q���	��p�'�XD�CVvB7�*�����4>��ꗃ��|��R_6���'�:�^~.�Х�4 r��6X�����Ÿ��r@Y��6F6]��AӞ���� 6Z�}jFG3�E��ү���NS{��p"-+r�
x��!9�$�}(�����#D�{s��xx!�16�x����bDv��:}<R��5�vMZ�h`4-V;�^K�F-h&w\���cI&�Ƙ�,6�8t����Ѐd���"���\C[a�:�x�5��c�
��4�v�� �{M&�M�#_(ޥ������7)H;���D��hZ��ƚ��~pA�=~�1v7�ן2�#��P�8��b�i�ZO�N�bw1����
���Zh�� �)|���a��S�F}��c*���O��*����u�'�xf��~Pn���Ue�)�r�������W���J����}|�st�=��H�¤
.�1ʶ��@`�X��5�@��j��0��	h8O��~�`�C�0D܅� �a.��ͨ޿1����0����x��=��`>fo>BC*l�O3Z�~'c-�T~�~��lox[�`>��n�J*�MG���i{�$�%Ф�r��(Nr�����y��9�!�w�OI�G!6tԔ_9���yl�Nܒ�P@֒������& �y�Z':�$�� ��B�W�F�42�G�Km�(�F��M���ϥS���o�ZF���N�˳�yM�Y��yaϢ�P�%�o0�l֝.�-v.�"��� C�c�z���/]2��H�!|���֐q%�t�l�
�V$�!�ӑj�l ��!����؞S��0�x=^��v�ԺA`}DiXyt��'��&b4X���e�xI�ME)�$�tN�z�������<�U��������I��S��QE�!(ۃ��ɹQ~���|�1���=�SY�y�}�'�u6u6$=H��9�o�F���D���GR�XZe�銼�������]��49���� B+.	�q7��N�z�s�f�F|W�:����
uN7R�T�,�>���ė��Ux�s)���m���c=���2р��#�}L��ob���`���E��������� ��Un:�V'�{4DS������0��Q0F�h�~K%j�K�`Fh�s�\�X=����:�����ɹ^�f�H��{M�L�;�t�>O����{�w»��1���pxp����ey]-3�_@2n�`��g��{\uP�9��׻k�`��ؘ:V����7��)�P��a^%��Jy�m@�6���@���
�)�Y�5��yu�Y{�F�a�3���RF���ܜ}��U0-Ik3}�����e1�9�I��f�T/�����t���l�o�7��Ӿll~�F��!̽���˓KV{C���[�<�i�� �6D!U�ݗ�Wl=� X�I����*S����m�J����{��V���	������N��vcL:P�K������|=7[������k���4\B8�KQ��nW#��=�G]�@�f+ӯsp��?�^���[� �!�^+ό�b�0@ݽ�3z[�!�nW��c��J؜z3[��ߚ?_?��t�6�rn.�y7�a������sGW's�fI���n��Q�����T��ZZǭ��N!1S[@��l����Q��,?���� %ϭ?�G���4,��p<#�YkR��2�N@��U{\,��T�R�휂�D3L�4��e���ݫaÏ��.W7�d��B�%:��A�T�a�;��?��'瘄��-��f�X]n���<�/_���A�[Р��罬g��"�ϰ
}��u&V�.�¢
R<��ͅ"�&�2! ]�jϧ:�P�O���QM��Q��*B{�d�A�q�V�J����a�w��Y��]a�`��ӳ���k0�$Dx�J� �lU
���C*/!1����	�M��������������L0+l�K�T7����d��XWZso�����:�F|�����H�Ѵ�oi�|���r��`̯�H�iT�[x=a!b$��}�B��>�y������Q�|v*�j�a�׷��H��;l�z��;_�ĬZ�P�
]kFB���M��;N,�m�=�"\�EHW��9UA?�(��nJ꽗�L�B>#��OO��nC�b�����;�����ǜ���B�l��2�b#�ۤ>H����0ڬ�&D:7V5��ȈEd����CMƳ����Y����+�E^vw���ۆ�68tڶ�I��7��?�� ��c}��ς�m4IW$��{<���6�,�`����a]�U��B�r{*�P1?�J�S�S)�=����f���J�;x�U���R C;�iXcS���/6--+�򜸺"�np1��I[U/�K���Q��4�OF���%K����a��gi�>����C����|��Tu�?��0m��Z?�U��
�����ŊS���5"ϛ��<�4׾�v�T�}�jY -99�L�xFj�oC1�IFT�ZT���,��GZ*
�[P����ln	���g ��w�Y�X�v����5�gMq�e��{����u�J�o�Z�Y���{o�<Ў�ٵl�I�h0����9�ڙ��F�۲q�&���S<��9��Q�#�%&�75% ��%O����,�.���V*�Ϗ�1��`;/m�}>�/+��"d"M-��i�(Y�|c*���z*�捭�k��q�����5Ȳ�9	$�"�^�bT�
��LZ����q��Y�v/�j�KF8s��{b8QUˌ	d��P���V�ף�f����N�`�����oc����ikNӾ�+B8���ݑ�Q�B2�3�1E��B��ʡ[a7���������K��͗L��:���kw����At���Rrop�
��$�����;�x*�	�&g�d{i���s��"��h3Q�#�2E궇���Q�Ȱ�r)(��d������]ጲ�	�d!^[� �,�h^�=�@% ���\i���V�}�ɟp���q�o�Q��=�n!`DQF��cDg�U�<���,��c�'����0��i\Q��_c���1�KǴ6�p<����14���/Uқ%Wt�ef=͇{����Og����"�7����2?�_�nPD�68�DA�&bt�v��ټ�˵�y���2lP;�\Q�q	:&)��,:{�$T�"�q��\�h�����s�\`���^�R�.
8h�%�����4�=4�ȶ�'�)���b���(s�ݖ��	�N���֡�H�"ై�O
pfX���J��F�M5��[Y�s���W�������m�7�[����TkO�.�o�����GCV,�N�6S�_g�Y�m4� {�M:J���nY��5L�����a�Ӈq��[wy��Uu����wT�X>Bućj��K6��CM�	q�߈�#k�ݢ�`%���*�����%S9��f)LoĪ�.Iv��ER�mwxt}cv@��C뀏�ڭ4��n��Z�$��yR}���FřjP�7w�wp,�9ɠ/7x$8=��W�;�*�@��ue
(�M�dѻd̗�X]��$UnɆg��VIλ�:@�ΰ����%4��iJ� {�9U�.>_5��G�̗��7����a�0��Cw�k��}��Q��)_S����g�F���W5f�+�%m#bc��-/wGt�lz3T) }5��69�kP�.��R �1��6o����)G�h�!*��Oje���ڰub����\]^�p����#�@h��W��JI�*ᮈt}J�<�#�V��o�oz �������d�~�-���z�
��i'iI��N�3�9|>���9�a�}Յ��Mk5W���cq�
����n;ŗ8|%�L���a�D���[��ݳkBQO)��|I�ܡ]ݸK{�T*I3g��`�La��O��W��AJi0mx��Vl�����	3.T�/.��3��#���H��e8�ޒ��+V={���G΃�-�x� S��%��[�����E��`�ǋ�,P	7.a.�	�[:l<NU�\1a��HM�u��ьWW�.��5�RԢVD��,^��l�/_��@�a'0�эa=�L�qhe�<^��E�(��բ�H���O�:�^9}Ts��%.��J��}N�8��[�S��i�l��Ɋ����P;�"�--�]�_�ćg����vH�����(�϶!;_ ���?F?�"+����T�͟'iV!^��I2(�6v����Ӯ�$/[���>�]-��2�S�>�{�O�=��.�YU���b�tz���ɿ���wU/fuy�l}:�(���0�̝��#�/+4	�<)�V��C��#��
�6����^�Opn��h���ޭ���'o���)aӎ60����G���Pc/=go�#!�	o[���bK����״x��ܴ�^}����ڿ��m�=�,#�у6` Z��gH�<Rx;��<����̔�v����X,W���"v9�J�̿���� 0m��F"�ï3}`����1��������ę�W���rYN	s�m�U_��~)�h]=l�Zz�b�b6t�\X挫����:2~ԋ����1 ]O��m,O��b3�|J �'A����) �y�b��|<���c`�����������x�-g����<-t=��m����Z9�H[�_M=p%fin>幺vUҷ��,�����f��~�g��3BǢ��'��H%�u:rr�}��`�^&�T֥�c���d2{��d8?����p���&=��t�E�H��C�B�J{�!P`콒yn�Y{����l�^����)�t�} �\�c����jpr��V|������U̹�eZ��C>E�w�$�uU��(o�Ր��N��Ia	�LM�3��vf"�>�-(B/ic�$���YNq���]J��|�0���yޓD]e4-�l	�4��mLn�D�4M��5�_>@�~dȏ�� K����'jd��<5�e˯P�`�=U��4�	�%�T�@��L���(���
=h�u�N������f�;�R6~{A%)�6��M�B��ZI���HeZ�!��fAܝ�4Ho���ZcH%��y)C��tk�KڥF�x�襕ݞh���P:6ߑp�}�v7��Ei��PR�jH���Z��aP�]�ff�).����e޾�w(iIe:shI��,�@�B�RIkKRE| �F�����v',E
K�n�-7�	|<�Ɲ6p[����E~$�����_:l���Z�DT�و��dT�Ir,j8���4+�ܓs�0!����9Q�jn�60���(:G��O�&�及[�UzS1B ��Ia���T >�4��XGj�N��'<�NH�q�K���$K<�g<��Ĥ�1"c���=��mBm�$ ��%�4��Ύ�C��p���4g��ʌ�J��Z�NTX}<�f�{����H�Z�Çt�^?}<��L�U&Ӯ`X����M5���ԑ�j���w�.��uM����ܡ�c�����>^�`n�&e:5%&���lN�r�66�ؠ2z i^ Tv�j��:{���-�TW�͖~e��')%j�����s��k �x)�$MR�0�{L�K8*��ib��h��)�������,r��2�+V�f�n��ݍ��E�*f�,�7e3hy<%;q=к��I��ɠ*�9�|VJ����% !�nC��-��SZ��
�s�$�.Vt#=c�Y�f���5��cVmY��&�yi��Ȇ&L(P��F�%#�g�:�fs����1��E[fX�s�)>�F�x�H�8)	$ߜ]��:6r!��3�#��VG�<�@4H�{sC��9�Γ���r\���M;aɥ���H�a�S1=��U6�-u�{z��4����p�>�M���Kl�uN@�DX�;�b�t�I�r�Q��Pwڄ���АI(f����`��}P1�g�0�C�����[�1D*�� |F�+t�I�����ý�
��j��#�w��a!~h��s�튶>��0� ��y�Cn8&��(a1$�(����S�[މ��c,Y	�J�b����2(,h���)'	Q�e�9`�:ZŞ��&tǝ��"�҇��	$N�0`�[�T2uu�n����������朮W-)��q�{������`�,Lqk ��ɞ!����I� H믏�>��������Pq`���H�NY|vpc�j��Nm���Y�h*4��³��~Le�p��U���<���ǢL!�M��P �B�ʉXfKuj���e���%{��.��-����(<���!ePPo|�t�V��zkW*�g�ʶA\�٪�O�1�GiU����JY1��wF�/'K�|��C�2]����H�)����촅��g�5�+o�g�b�����>� O��Ojۯ���6H]&�R�J�p-�����Q�Ma#ʓG�����~"\L�.���rn79\2�xM;��u��V�K���׬٫E:�|M����tN��>��ml$�Q3�;�$��قѥR�=�z����l�[�"�r�B<ݎF.����=r�Aq6Ac|�=h�� �_i�X�.;]�Q�����iK\�U�
s�XeC����P3�? �4�h�7?X���¨s��r����Y����_$ܽ�J[u�������}WGNjӦ��?ύq�N�Z�.��#`��5!}
��|_+[vK�qCݒ��W�C�'�`2	5���R!47�{��==����Xy=r�&b��)!H�m�6�-�{�|~�rYH�sf��(��"��|t�I'h-��c<�����g\ؾ��M��/���Vl��`~Ť?�TǇ�w�ŷ�O��*0ǈ��h
��v�	�x��<M��=�8�BD���9`�3D� ��:	;h�+Jb~d�+���[�_l|�CB�[���b�๺��ri�A�NlĮq��^F0���L�I�P��l�8�A�ږ�ܰERRPB��	Ų[��3ި�_�Py9��b�X�I�e����7Cm���+�K�����$���&�3�w���&�7�u��k��*�641������}�	
rϳ=��ڶL����G�Ζh�+6Ƕk �`����%+9�=:Q�;�A�p[�E��E靖��F�M�y�T},���q�t�(ߝp1���)�B(�O����+�.?����H��w+��>/~+C��]���O��U��T�K�0!Q�v��_D��U�X��ɚѵs�vp�Gx$ς��&zG+�sR�o��.�6���
��HUy$�FU������Ŝ�"y��dc�[�=�	�!� �^RO�WJ��rk���9�D����Q�>�:.��3d����m(F@�/l�}��]��*�l�6�7�O]�+z��XcW��6؈������JG�7�y����������;�^�։}����i���׏�w�/��6�����_rϴ`��d��h�bI���
ŝ����ڤ��r���F �ںQK�>��\��<���y�⇊����
r~	[�hҞ�:�ݨC\V�6�������dÓ�����/��$��V
<�f*��a,���{��gx�A���dD�H_O?���d$��a-)���K B���;��pRs8��s>��F:�pY��K���A
V��y��d+���-!�����/�H��/j8�`p���7;��~vBx��o"��Y�J��}��]�a �&/Ů6,����t{s�GF����us�z��,MM�;Sf�eD����`���!�y�}@0nHa��d7�� �Rn��i#L�Zj<�6�VHeQ�dS�r���d�!n��U&�}c��#��aDq@b��=����|�f�h%�KV�`�g�OW���OL�J�Ӱ�kH���PM~��2�A0���Z�.���Z0�oZ���Gbθ���z+�Xa��
~�S�<�3��] �-�c��72�VޜΚLҷ�@iߖc�1w�U����$��`#� )��&�z��J�gһX6b��U��(x]~���C�`[��D�
��'��<������*��CE��6�D}�������a� ���@���gg:: �p�Rkf��g����>��7�A�sw�f�3$�M��ڞ$9�x��{�Eq\LQJ[?拢5��
m�_�:e�����<z1*�K|i$>��|�~B�gFO�0i�3�� I>:�f�H��dE4+��_�dK8W��u��#;y��6+"|F���T�μوȺ�K�0�؊�#�VRm�(����1V[���\��!�&�4Ѓ����)p����Ҝ��e�C��28�ӷ��ʖ��5��*�"�N������S��_VPo]�d��LKf��F���y���J�6��+����]��?�s�%���8�N~X3u��;\ �����T����aJG
�6voW�<���V;/�0��$�y
J��o�g�Եxy���utϳ��D�P �����Tu 76��T����ŵ8t��g�ޓ��Ho-#p���D\۠W9��8(����-�k m��B�nP��	JT�=s��J��C�LH,[�]P�Jj���X�d�Z޴�k�|H2 [n���r�0v5�D[5��ը񀊨f�t����)ԩ�#-$�=z�����f�wζ}��J��[�ž��9b�x��s����3�T��o#zg���<'��{�7(��~��y�t}w�n�v��;�8~��!)-\|4(�#��Pk^��Gw�xD��m��B���v&xE�y!�_��Iuć�\J}����J|~;9�BY݋zڠ�i�8���l]��)��d�)[��,|����l�1��J��(�G�J���aii�'A<ƈ����<���H���HQ&R���U7U3E�jf��oT��3j�灂�(U�� ��(��\1G�`/��Xo�����ڴhv�VY!%Y�N2��"M=49H�7W�r*���M�s��N�/����H���lCKFs���ڭMI7��tIy�o�5��)��򓿊v��S�����ؖ�+N��a�U:�oR����}Q������*�<u?��<��ˠ:�s��n��`�c�r���;��O�����f)�--�`.M�������2Gcl��W%ٰ��W��V��
���#l�k8�e1; G��0Ɯ�,K�N	y���U�3)�Z^%}\��p{Y2&"��j*^�Sݐ������MX�$ÞΕ���-F�=�#���Ң��*�?*����i�VӆOl��B��tT*:i1k��'v��d6ZjI���"��;�0<�����M�&��+:�7E;��m_��B]ò[+�/mC�_�W,����ŹUt�\b��(ZOD�e'ExL�
%9�׮O���77Z�n!�ۛE1Ͼ����L~��r�,�ht9G6ͷ�&� 3�%�[���g?.�D�8p���s��֥cK�.�m�>�!iU�b6�� �R������-,5�2����P�E��[Z/�E�~
�$�܏i���]� Z%9��i8՚\"+���o�T������Ӽ?���k2v�b�ppὺVu�3<PHa*
�l��䏸�,JU2?�g�KNcQ�Oq��ٷ����Ǻ�@7��� �X;eZVQV
0���EL��[H��ARx6OH]Jɣk���t=6�?��E8@w3��ai�sE���?������J�؂��4R҅�M�`|��;.{����>4C�#���E��m���8es`?��K���<� 	��n81D���
�y�JO-w��fN��l�wN�2�R�#M^z����������}�!���:Q{���up����������;��w`��\�h��5�?�r*�r�ݐ�V>t�_�<N2�mj�>/��{>�UnǸǍ�M������k,�$�n���m���}�)�"t�l����`hˤD����k��[6�y4|�z�szǭA-%��<��}��]m�A��)�7^��n8a��W�)�WvYU4$<�6𝷈.��_���]�͸�,�5����]?΂Z��u7�Я�ܙ+�	��mĭ=��<��Q�o��$1,�]�e�����.9fS�d���$	Z��2�Y7���q�P1�RŚ�rOi�&�~@��4��ٴ��v42��59� ���r��̎���c�<�_g��׾f�� ^> ��m�	��4��it�}$;7P�><��)@o]��P�&<7��:�{�a�%��>�G�$�c�m��w����0W>1� x�6C�Ԭ�Z[U䤷/HE�/�FJńN�4��*�aK� �M~b�KpoJ�YvO�Ȋ��b�O	c��66[w$f "�c,�k��nC�R���]��=��6^�R�g���h#or�Q�(����ئ����,w̮/�nEQ�x�}�4�3kV?cB�N�������)`VB=<�n��Lc�L�'��k��M�4.��_	0#�$������6ܐ�d#���.0�S�"=�	&3
����J��i�yLۀ�RoTv�P�Kf�ߒ?�34�5x�J�5��ǵ�p��ԗ ���]�� �����!b�����|{�7,�4��wS��> ]a�c� ��oe���Q�_��&��@��S�̦�$����N7r�m01��mkjSp���5��wH�.�nL;oF:HĽ@���N�f�� $��d�"����G3���h���,� �ʂ5k֖C��0-LJR�x{v{4�Z�c�U�dqƕZ�-@-�Y�Ѫ$��;�W�9Z\�S����hp��0��>�E�؅��>ɷlo�$s�q*%�F��C�/� �KS���i,�D\�c�䑥�e���}����IN�K���~[�މ�`�)1Y��V��z��oub���4���B�<����Y^iXQ?c��+�k��'ݰ�b╲�k���S���	Ln,$3��AI>mZ��fw���-�3&U���	����x��"��ˋ+A���!tG�*�a�T��R�89b�e�����¿��\��N�3y׫�E@�R-�r��}��n*n�"Y�i`,��R�EUzn�d�$yٙ\����Q�)���Ym���8tG��C 1�<��I�>v�bre<��5-�a�.��Vbi�i���R�F�CTXۗ-$FЪNϴ+�O���F+�5}g ne�W]���AL�N6���L%�"|�D]���Y��kZ*�4�V�B���R����+� �@,�q���B>�Uy�����V���W�R$X�Yg����d�D#;�)�F��Qu:Պ�­�-��L�W��N�l��U��{���ʒ���Qnh�}~zIBvOL9!�5�͢�Xj6�9j�������o��v�P	�|���7Z%�X/�|Fֶ#L���k�O�`W�%��Q5����Heq�Қ��nO,[`�W&o��Լ�
� �0���u�+�.�*-Ԣ9�� +j�Q�U��[LX��v�o��Uw Cft���z�<z9��3��q8uY�v.�64�~���9$Z�x����F�M[q�����qL�(��t�	�tU��ڏڼ���O��
�?qO\pE�29�݆RdJN��;ք��P�sN��Í�
J�|C0����0�J��NM~(PC Z�����@f@��5���Y�ݰw=�$^L�B���zW���QWڡ���A�`���7���5���A1��كzw=r�v!ݒ�΅���u2R�A��B���
$``�2��yj��˦�j�z�#7��oP,�2���{l@l-�|�-��b��֭(��`	
�T$��R���g�(�Ԉ��{�?�@p{�OVj��7n����Qm��j��P�*��NR�����=X�� � so>�����c�6@��u�5���?�uK�-X�6���109g��ޕ�aج!� ځ��Ce^��%�{@V�a�a�/<��+s��8��0Y/2Zh�u�i/(W�1o&��rڻH�S�$���z���tY���%�i�Lb��
:��b'�KN��]��l�_2�U���ʷ����*�&�ޟ&uș3@����^�b�(�M���� �e�	sx���>��i��oBM�N���2���W���߾}�G�a�Q�]�dT�8`�-{����ޗnF�E"� ~�������z����n�,��*.zh3[��64Wg�#M�	W)s����4�X�mh���z�i�K����em0�9�TǏ��ځ��}�Xxi!�|��oxaWł�ڥT�!ߪ���D�d�/�2�m��Ф���6Ր���	z�2�-%N� +	�6�j��jCUgs�ő*�8	W�*K2���E��õj�E���9+CQO�W�:��S��U<N)���}�5��_�h�~X�� cC0��y:��9��Ȗ���{�U�,�3
p�~�A.,�h����1�84դ΃�jq	h��&p�5#�����\k���V��)e�ڎn���1��G3Fn�gյ��������&\ڃ�+��F$���s*�6.�~W)�<W�9���a�����6�����-˙p�����(o�:L1&�?�ݞ�P|��M �7�6�pp�X=5OJ��Y}f�Vy�RS֗�l	8���.���'�rz�g�>����.�X�:H�@��*���^����}�8�UK�4בR<2���~>�U�0�Y�UE2S�D/<���^�/Ы��. ���
�U�z�B몜��)�H�� ի�L���+Y��{����Nf�d������%�i����A!D��g :������`�K����T�ƨY5�,��CsZ�=�(R\qOV'o��}΋����~��eXTy�7��L?�<jl-+(��*"8n�\;'n�?����m��L�:������'����1C��}0� ����d�F���|�gOظM��zX�?��ȐQ̅N�Ukx<����t9�wn��
1y7ڧl�gٖF��.����u:䪖$��=�L��~�x�0���[.���Z03_t�S��8�r�]��Y*F��,`.�ч�-|8�=� �o�M�q�]r����
c����]=�b*�>:0��5�=o�`)x�/�:hÙ�Ž;>���v�O��Y �y�����C�m�}+�+����&dtoo8C�a�{D�D�ȟ�C�ebV�I�OP�/һgpe$x�Vv���47�� %Ԗ6*���C<*�#:y��.I���]c��׽;�C�[N�V���i(�Wx|A�?[_�D���HTHAH :L��y*7�.x`g_J÷�(�q"�{ � ٗ=_aG�/N���V�&�5�����ke;���:o����T{���6�"�6J��_���g�����V�j�"��x}v^�`�|���;L��/�o��`�2q��1me��P��Q|q����Ã����ƞ@g��T�(��:n=?��� �ZJx���W$�Ah��)A��gl��bz��hq2~��Ti������w½r�`��Y�o��ɇǩ�C�������qRU�B?�lW��T�X��7�`��m�����G
�`�,*�N��
W~��\��nO��jl��]�������t�㢞��b���>���H��+�D)s�aZݥM�"�l�w7v*�cA.Њ��3ǦWj�>(B1%��1J�N�,ѡr���MMy���}}<�����L������*�1m���ك7�^[̅Y�nud����^3��APs���:q����!��}xz?���/� ��L�1|
��Z��j��p� � �V�h�&�Ѳ�G�Ҿ�����q�&n_�/C2E���@G�٭=��*��Y�큆���D�\Mh�(�p��g7����$Lx豆$Q�IV��<�[�ޤj��ۯZ��q��t�uŲ�	it;ż �([A��f/�N'84���Yޡ�c<��tw��Y4����jG��:ʅ����0�!>p���f�F@�xK����QW2�ͷ�Ɔ�J��`��d���#O�z��
�9��rn��7���s[@h�穞���i^g�6�h��
��qM߃�v�큲�G)�[� 2
���4fTU��4,��U��zhQg�=�Ļ��_�p���}6c-R�6��?����G�`ڶ���32��3GG�^�2!��O�	LEI��&e�Y�]��Bs�n�
�o_�b��t#2�;���%��g��3�%K��&�g����>��ٲp���Hd?8�l�T` 7���촮C���D(��p@d�գ��w����<��Ż�F�g5�O�<T�����C���ٽscivd �Ѭ�c�T�]�2�&͢N���r�lF�m̈́�l̫6%EvP�^�+��������#�ֈ;|w���5��`�ш�l���Ǯ��V���"��������K�8{��h��Tyg���C�lUzPpT�����"�� n$�q�,��{]�	�i�E�e��Lq���F¾A5:�4l��2<C%\�b�V��"|u��픅���������9�_��_�K��~���|N���/��DA�28B�3C�5)1F0]�h����Y|�v:��/ �bn����-�K~�D�1-Fk��Wy^β�W��k����b� ��z�U�^��s}GS��gָtЋ�X�~@U��(�~�����?�����V��e\��
�2HJQ��h>�-,7ԛ�E�\$��z�9�| �@�'�F�aKg��oiS] �;.�3�p�o�o���v�/�����_��X�~�{�/���U�g{��t�0��'U(+�3�����>W9M����-�99i�l�Q� ��VX�#a~��m��#�Z�{VSF4oPU�(:��$��n���+�J�/-�����̸K�o�5����]4Rl3��/��>�2�v<W!�dz�l��G�K��r�﫜����E2o�X^L��� �W�O֘]|~�ܚ��&�[��,�Mo�����AQ#6�R�m:m��%n��~�D�?~z[9��H*��`_�1ѐ'�������M�N��nF�a�W��;�	Y� x7/7�����")��x�[���~d�өU�8��P����	��3�,%�����^�m\hM��S��q���c@�.`a�
P��-�{�����f�_���<W�fܾCo�\��8�(%�(��}I8&�K�����,{zo4�'���߻�{�['t5�?�C0�M|�0���������T�[?e�u'dp[O��m����%Jr����f"��	#� �������ۺ�� 5��P�ʵfީٳ����^iuW��k�c���VH�Ϊ�^�� fA,����2zb73�|�r%�=�J3ѻ>�B��;,�$G4����ɟ����zږ[���0�v�t�e�� �kFQ��k��
_����4|H1q��h�J%ώ ��#M�����	<K��'�i�1к������/���mK����<��7a�Nӗ�w��1Èu�i�Zb&6�d���()�u�VC�EE�Ɖ�-"�J$}�$����8����/�±��Hڤfc*�8XNS�lg{�0�������f	/�Sl��>��аJY�zQ�c�A�с?�y��qJ��P�-�r|�߷G��sr��ۏ���ߙ���MU4^-�����D�}��K�Đ����)���p��a���+���ڕ?���fP��pJ�l�'b8�k�V��ĺ�#�=��1&onɳ�n}W���a�G=�e�K�1+�K5���5���KH�M�r������O>y�����i˶v���������+Z�j�Kɴ/�A������n>m�����n�桏5�&ン�Dj�%���>�O�J����&�|��ap��H�+�`�9���?vb-h�b*ֱ��XK"j6�g%��e>w�咉�7f�$�ݨ�O����N�����2+U�d�/�Q��F zd*�گ����A�@.�?ћ$+3u������T�D&Q�� ���>��Q�]bgjtk�DT���P���L�C�ZKڣuM�4O ^����?pW�MT�i�E���04�1R[�>xB'P��1/6go�4�q�ӥ��,�������
tM���ǽ�L������n������td<���v��:�����2uc�)k<�I:��h!�:�]��	z�}4�l��[��f.;I#7�u�����1є��C8c;~g�QH��&�����΃���S��ٸ�y����Gk({�fo�f�gʌ3hI�*x(L"�/�b�ڦj �ok�e�5�=5�8&��Q��9�n��R���#mq��J-ɣj����?�KJar���d`�QK?��"��e�,���5�f}L�����¥�b�2���*����TTW/vYJ�1����,>%�4���=�%:(��O��T��À�3T�D:�H}֣�z�_ڋ�O�����V�tB���\o�E�X�D��T	E����w^C`��c�4��(P>"p !`�̍�A�<��b�$h���R9سW��ޏ�S1O���P6w�B�
y�>ͰP�Ӥ�؞.�$�6<�Է��!9����wpF�!Õp�R�űTT���6��@�-i�([�P{��P�:���8��r��ja�+z���?Ԁ��M%v��ʵ	�@2&�I�_��#��Sb���=�w��,�p+�ڏ3�'(\�^�yN�'c��`7O����Y���aZ��%�������|"�_�[y)�B���c�0���`َ��껔� �3[�5*��XD�[��b��_�����pF�%ϱV����*|�����l�ڷN���NF���mT5����N��]6gC���SB�ɠ��m-�~�D�ոZL�ɾ?٬�;����@�+7DPAyLy�<��C���(�|6��k��)|���8�ef{$=&#�0V�I���-���["F�`I�q���V���$�gZ�̕J��!���95�|ݎ>�Q�L?�<R �Ȑ�6�8�U�4��s3�t��6�9�8=�0�q��iS��1��3�>Eu�[����-�ީ��j^fYj��c_����j�>�H ��:�L�w�w��'^zҧ�]����;ad���Ë�;��'E�b�c��2��d w:�z�'FJ�:����	~3	��J���z�_��Pw�	*=�M�q��ʀ�]�����ļ�m��G^^�����dL�	�O`�E�`�YgA�x �������젱�rˊ�9���e���m����9��O�z�`�&1=(`���Ղ��cU��p$Z��H���uH&�5{�A��ְN4�3&�S+d��g�Z#�µ�
9��1n��[e�h;1*C��	v+HD.àX���l����ʕ�/IJ�g������4D�j�vo�x���I��/���� 0��G�fe
�0�J-eMh����iG��O�j0��%e����%O��2�+�$
iB�y�X$@\�Z��J�EԼGXH�)b��Qج��O��&�M�u�l�"g!DN��D�̂�у�Å�?��^B�Ъ&��-'�~|��H��;{����+S�D~+���d���b����#|һ�@3ط��EPS=���\Lb�]�2K
��N��WU�����]�M�:ôOo����:1��%��>�]fN��/6�N��M�F�gZa�Y'�R��2�Uy�Q��c���*���_�V�w�n��j8��Y{�=����my�
%��j�y�Is8$5ѳ���|J�I�ӸL�`�}ζR�|���ۄ}�:5��_�L@3�nm�;Pײ��tӲI��M��>�n������\*�,|��P�K�
uaQ �;Ly�ف�8�2����#R�w��Z �JlMM6叞���A�=� `P6��+Ɇ�Z������e�l�#}w���$z�콚x+����|Q�)Pf����cEͶ^H�xdЬ\���y��?��op^�-�:�q|��@�3����1КUw�\J\�n
���2�����.P۬�����⠯D�u��+[���	�|3��c��znHR��� ��#*W~5��cf7!7�ϡ����aь! ���[�f
sZ7Q'��r��Pϒ���_�߾Bo��Ȥ������t�ā��tω*��@�<'��3Q{�vY^#���
���s���n�6���m� ���h`W؁/�4���i'��S[�7;�K#�R����oM5��0iW
�4��0���"C��;H:I�Wg^�T�Qx}���
Lg���>��R3�m%�Tߧ��8��vPy>V�8;�]��(܊~���(e#{�g�(���^��	{�y� R-�ެ0�P�O�X��ם�Q
(!�GC�v��8���:Sc�8��D��|��h�X��l��G�0�� ì��!
o2����Dv��n�U1�#�H��܄���zY0��zwz�lek��g⤲xg�����Zn���ʀ1~?2�֎�1A��}S*4��{������o�v���5.�����t�,qރ�6�����Ըk�¸�y 0W�ɀ����-�*�6���"Rh
�^-��m��R�,��	��^�<(�U�;;9����eb���PY�ϐ����a`X��K<<7Oƞ�r�G�^�9B���b��ð���-Kc�N�&,l�v4 U�)��v�4������Ϛ�Xڈ���W(?ٕ�!�'�f�����On���T�O�^��!�&��#��Ӻv���O<e��	c"��}	F�_ aJ�F1���"��m�Q�O��b�§S%�vB\oө���WJ'<s;���l��4�� ��Ę��ed~�0�5��|�Q�M!�)���>`E�G>�䯦C�(�P�*ggh8�� ����_Kn{�%-����'�����̀�~�޼���~��f�R uQ'��%l2	�ͅ�
B�0]S;L�^��ݳ@_e#�(ܰ#��_b�9�n�&�χ\�H,�5��J�#�<���:�6L���������\zx��.b�5�	&��9'���%\�BR	\=�9z�2M�%����ެ>�n�];��F��.���(��[�����%�AWq����M�oA�6�RWE|�2R�հ��.4͌7BHY�>���k�����{i%�8��O,�&Y�u�az"�#���m�r�L�v<Y���5����aa/���)��ҽڴ*JY3(:<�fh�(�"���m��F>�M���.����9˘8�m��49>�l�� ٥���-�I��Q��	�#6�GG�L�:�>��fx(G���j܉���z�lL�|E�viN%\(b�h@o���kp�7��f�܊?��>�x�$�M����3��juXY3��4��d�HYMpN�l�K���b����H�`�x�w��b�E��Jh���3��1^�i+'G56�����9��-<���|�"�˼�g��/�,�a���6y-i�-��Bb-�0����teB��}�>o���6��ː)ђS>H��-�dӥ��'@C�����ϋF���L�+K��\�e�0����%]���h� ��?9�q��MF#T��L��eW](���(.`N�PVX跑��O����5�b:祥�3D1i��o�v�P � �cף���x���*������_�ɑ�E�[��+!���7h𫯪t���[�p!�+Kh��p!R���K���Z����|��'��_���Rn������`��|���E�Q����X\D3�����Ǻ� ��>�l� b�_�SR��(�a�`�i��/�,ԥn�!gz;_���G=� ���JBQe�Q�+w2��5WՄ�I�n&N�s��r��2+|Q�u~ͧw����a���
7K_�
+��>�U����I�	<lre*i��=g�cY��s`����w��6RH6$�d��Q�Y�Ah���]"�e��c�"��'s���&�q���gE�cݯ���^���"L5v�ҹ����ct�]t%S�%.Aί��a���OՌЇ�T+�bl���`�/��]�|���s�/g���V؅E�\�G��w�7`]Į\?�����_ ���uw�9�9˓��O�O��]<�%U��\�3(.�[��Dq&۩��^d���U�<o��P�t{Xw�����&r�M��S��ۀ�ݺ�����-^*s�3���H�>d�W�'���.g�xf����b��C���z���CLd�^��G��$��$F>��#y#�o$Z������2�X�[]�d
��kl�n�NէC��\�r����%���-p	�G�Gӷ�n���)ql����띐S�5y2������:{�dn@�W|�O�� w�Ȏ<�?fn������n�YR)�CILED"E �b)��)dU"MݺB��{wX8L�A=���H-�͡�����0 _z*����^�X2�E��y�����<��5��Jf�`Wphk�)�=G�4a�Hq�1ǡxŌ p�Nh'}��]�V��!�ry�A�ZA-C����΃Y+����kf��s��5���-u��xF�kH���B ����A՝��
�.��mB�*�K��؈q9�`�<F�0AA
�ݣ��t���J-� ������\�V�$��G���~X��y|� �.��$�e�eR~��Ĵ(��c/��LV���§Z:=a/����$�@�Յ�2-|��: �S�P�c�!
Oz�<�γ�,��@�ȯ�H������J��!ku]��������XK�X��O�
4)lM�,CD��T �菄��%���*��T6ی�B����=��)��1�b���f��u���҇ڈ�A��k���<ٲB`��G�W��(p���V�L!�z|��"kp|��W��o���<kN�����%�C��K4�1�W���)n��NJ[g}��(��}$���kA��:h����Q�N�J�Z�;H�>��N�a{��`}�>�W��z��a���f��Ƥ��l�e�_�̀�&�w�׿UΓV��V���T��tn���RI!���.{�rt/���}���-�z`�ޛF�}O��\	�Z �#V.�T���N�����Gv�b����s��^ZQ[�1��3��ovn�^ZqL<���}���Q#��Uix�������C�7��3���a�?�_P������4�"��o(@�P�>���$���K�����v�V��V�-�m&!�>l�hD3�V��*Wyˉ�X��m��J%W���n�+z������cu�}-s�����:j�hCuY&�t8�E%�u�#:J��l�V>H��9W�:6�p"����PZO
�z��x�>� �"Bʎ6^|�U!� ������NE�?� 6x�w=�n6��Zh���bŢ	c�7�7��տ#��J$ɧ�E�a;�W����<��,��O.`�	0U�#�x&1F���������לZ�?�s��
CP5s��^3t�Ԯ��q<�q��k�	� �"�l�QbݥgH��W��3OR})�@b^�H$�J�#LI�'�l)��1��@V�����,�_�o\�V}�=;c{OZS��Ǿ��1�1�6PM #Ā�	Z�2�P��0���T�G�OV�#��M�oȡ/��%��j���r������L���;�
̸fް��2F�;��gײ�-�4��<inA�к-���h �S �:o�EY�Z�>=���סw�6$�~�=
��{�7�
��H$��K�
0�x:��!�j�&��Ҹ0��G\�.a;;Z���d@�]8����n7Ȥ���5�g���hܲX#4�ֿ�r�jA"-#fgm�ـ:��Z	�����}s;E�jj��\ W�_�ң���JS߲���W��� :ۋZ8���=8a��C2�4+]�\�{ē��Z�x��O��j^km�e�ʯ�O�jF������i��"��zN\��U>�pZ��j ����\�Y�6�dI@���@��f)�z��[E��K��>A�.�`���hM�^QY���%�Q]�Ѿrg<m%2�_��9
�2����P��r$�aw4p��
�-Y�Enպ^O�
N�=�v����,�F��ptn����"�+Z=ŉ%pi�o�s��d�|�MxK�tæ�z�T���N7�&���ҽ�vs�_C�	������^?���-����pgd���� �����H��,_�V�sq0Ι�-H�$��p�]/o����F�p����x�e",v��'2�2�I&�p0�)�h&}�[������9�q ^ĉ�z$���̘���k���>,
>h��:�2>s��ď��xm�}��H7��)kl1\Q�KpSE}j0�>?��r߈n$�_�f�d�w����y��ы��ս�Z���k��@+A%# ������QS+T; �8��䢨�Z	#t.r�:�*:�k�_�ρ8=�� Q	�}����'Kg�5�Ň�Qv%��Y�,�c����:c}ǂ>�w����В��׷򇌕�q=�r$��x��b�
o�	�	h>�&{Uxv�8�1P���� ��?#��qg�4	n�=S-��6l�3 &�RMr���5��⸽����}�3�Zmm�4�'p�; ��1~�a����D�Y�$�-�q��C����Zy�=ĸ�W���f�Ţ.��,HDa��[V���?��c�r_��A�dg0��0���g�n�E������:�$�*��4p�"ƛ$�do�� 2�\b!��$�w�ˇl�ڭ5_��'�B�����r����PAYtyd�N���1,�.�Ѡ������-=���^������lC�<Q'�����vVWo�e�י�eĖ'�Z�]�y��&o#ԴN^pI}�W}N2f6.��j��<�ͥq'��P��)��G����+j�XG��Et�J!	����#97����q����A#
�	������7�=4��|���W�4�e�o�ΰ\~A�f�z���x�DXf��焾"\l� BC�3M�ڨ'���)������Y��>>V?aA���!�CbY$��I��"����0��Y����op�S}�(��2%dN����Q�g���s��XW��kg���*�t�/�8��/�4��,"w���!���9�^��Ƴ��X~�-�eM���j�PF�����w<.E�]���J�k��5n���ų��ҽ�dj�������*��o#`!�*��VG�KN�ڤb �� ��ՑdbMc��u2��]hA�w֭��8���QQ�w�όM��n����l�;ih9s�8�*�lÔ\6)��ӯ`�i`���c�>u�\w	>����<��P/ !�>�q��C^���I@�%R����qg���\Փ�mشۅ��HG��e}xj$�N����p�f��^I�N�~|�,q��tHMlF�+d���V�	W(i���֮�*R.�y.��]��Jģ~�5��t���ԑ��Y2 ��]!�/��e��c�тZ2��f��h;θ�Uj�-�O�ÃKwL�%1a
z��X4K-{���6̪A�iGdԟz�:�V��l�#6�㰬BA�o�܏.#���a���\8���N��<�&��4*�y�k�We߸�e���C2RfZ뎡h��6��3A�f�����H�p�o+a�mte>ջ�8��' �VY���:(��������*�He��%���\�X��@w%�|��;��l�� �En���j�Α�
,[�f���Fg����O���� �ʀ���; n��o� ��S���zv91��tb�|h1�e2��U�&�K;�%j���['�v	�W>�f��\���YƼ'��v�*To9�Q)C���zۑm� �%���!3��y˻'���s�-H�௻F���\����xp`����*O!AH2�b����0
�vK�.µ�c�]hƲho�4x9�Cg�I���`�)һc�p,H�_��;&ˡ@xJ[G8���<�A�'�`C��M��h~���@C�Ya#�R�UI>Ã˗r�Կ�P���q�W\�$�Bʝ���b7��k���Г�Mw>���W���?>�?&q%�s*b����[����[�d��L�
~��{�⹘��cǺT���z6��+F���]�յ��e}P�n�V�-'B��cA�3~�W�[��XVS�taO�$��K�8T�8��<��	��t�����b��}�0mCL���(�$���&gl1C�OV|\�z������;����Y[���C]^O7�t^62��t�-9HӸ�:�C��Z��9H	�����rѢ"��XLN��Ȍ��;�������^��W��$z!i"���55E�������B��S?��=ܕ���ń8��⟜�u�7��=g��4}\��;��9ڏǋbv��:ė6��X�� �~�ħZ��1�����i�9�LP����Y��4�/{ j#�%\��O�-��әzR��@��̟4dE:[�ئҕ$$C)6��Un� ��tP�4]��U�;	���x�%U�BȂ�p
�+����>Kw<L�h������s�c��OD�[��mw&�ǋ�(\c�7�u���~�J�)���ƃf�{m@g�������'I�[��:iR\.rӠ����X�U@�GL���T�`6����I���4C�����)��^�dO89�0�����t�[�/��0�琉(l9���4JR'Q��w���͎�����&������w��4Sah���>LD}�Ϟ)<[������)�)<ͱ$e�E�Áqc�2���ӠM�~5j���[��� ��_�k�^��)�_V�t��v�Ɋjr��s�~V�Jء�x���q�o�?���2w��,�>6�w"�Y�7$�J��י)�l�W#�e�a���AȤ��L8:le��)d��v��K2���]:�j�~�RQ�'�����aGW��[����jǪz�F���g�ͯ�����7����09
�ZC�>T���_r�>�5"������d��z��#�t�@��0�K�����yIF���N�p�70�$d�J0��1�)�q�h9���Q��?jRC!+h'|��c +Ut�E/����ڼ����\��j�aT��
N���n��Ƴ��A�>�xw��L���W�"R��͢2^����V��0�ПU��'XT�x�=���4>�e��x\�?w��}�}'a̢�`��O�Z��1�Џ�=��P�sa�c�?�	O�؀ϙX	�)�.���v,Q`�K���d�R
�5�aTLu���f��q�:��;�ҧܗ�(��1a�.�����P��^GXf��5ps?���>3�t�N�\�z��[T*���X)^�ж?O�i��	�Hi��3i���{E��z]ݿ �+ڱ)�3�޺�{Z'%�y)_�w
5 Z]�����Ƽ�J#ױ�E�u��jb�Ι*�I0��W�kx�3��q ��w�	`�I�t��Ÿ�#5�n��+�X�j�����};���m32��S#��v9�Rdd�C��R��1°bј4zsŋ�j
�L���P��ER�a��d�p �|d�i�B��u������(�!�Fq����ظt(�����2��F47W"��;a��E��}ҝ���b�,煢S偰�Ǡu��V��&��{d?-�N���[�M6%<� FAN��wL���e�����&�o�H�e�����F���S��!Ǻ�~vmKM2٫��DBx�2�ٛm	g,G��R�G(�TeZIt�`e�Ď��^�'5��%x$,�� "�(l�n�˾�}������b	���T�ۧ� {�][�g���I���G�_��!�'O<&�ҺE�_=n&^Fv6�:kpQ#�l�`����g�Zsk�B��p::Ҷ�@���������z���tC��W�3��D�m�r��ēRO+v��?��������@��|��{�_�{�Ҷ,�VS-H��ol5���_N ��ݚ@� w���S�u\�q�2�PA�1������@�����4��c-v���ƹ�^�m��*��lj�y�'(����J+1Y^���j���ۯy:Q�(�����l�U��L
u�R��Ts5�d@ >
���W��Cn�7���aг����-�%�%&������l��&��G�a�%g}?ɩ�����η7J`�
��쒥�ݬ�
0�"�I�In��s���	{�=i����7)�+���Io46�M���w3��c�^Ay��\�݀9��	Q\H�����+u�S~N���,�v�l�7ꥆ8�[9�1����"c3�����VxIY�,� ����a�Aj�|��[A�A� �Q�i�5��tv�D�!sE[�����u���"���Q�2�KO�=,��y�wb�m��u�tq>v��7r�O�$��xδ)�x:!��KF)kR�_G����ϑ6�ѧ�X��+���,�N+�;��(�h�E���d��I�� �fpF(΁Ȼ_��Hmc{b<�~��{US�#:� h�E���Q�s��]���Oh�$}L�y��ɍ�_B�y(���e�������&S�5!Ԇe\C	��ˢ$�5K�U��>��sX)ễ���#��3��Ɛ�κ��m����uo�ݪ�y�+0Y��G�
�)����}!���L��'I�&O��3?�m�	�b2A�r����JMQ�k\���g���O���0��^\z&O0���Ə~�����t
��nTƶ�Z*�w"��'�;&	j�̰��i��|����Q�}��\}�:��G��z9�-�T�|D)�7Hx�7�A��9��a�,�=����tiM�}
���;�
�� �օI꫙��q���꧉
&ͧmw����$���7��*Xe��ZU���N?�ng�j?��j��Vy�nҋ�%�\V��z����p6S×��E�%��X��5�Z��7��b�������SYh�e��:\x-p�eo���s���`1��}��ʘ�0f��T����r��<Z3�7f�g�u�ٱ_�������/X�m�}�i~��KK7�R��o����9x�����HF~׶�c����c�7��a�̄5��Gz>�n�q�P}���qp�^~+�F����S�x꧛����k��g�GN�`Ӭ������	.���-��6r�����v*Ǯ�/�¥ſ7^r1o��j���8=��E�l��a�X
gǸ�ż�CmA$��u�g[B�RÂ��>S�(���3l�ԛ(xF6��3���e~U��G�{�AH�p��\��"�#&����ę{֭yG�F��6b�0)g�������2/�Q��>�X�]
��������:?$����>�Y6�4�2>�^�\���y�m���|���6��3`y���?o�.�+�,�_�|�}�p�"qu�����4�%akG��N>R��0gs�ʌ��6�m����%Y��=��*:�Fk�W�	��Z�F�O�{{��
)�����pK��s�h>�ض��ҩ�̹����'��w"-"&�L*��������t+$��4*�S��*���eP'.c���N�*�:��Y�=�T��I����M_)��h�r��bz;3�C�8�_٢��p��R�<���z����.��<]�,Hߏ��'���UW�&&�����⑩�>l�]zr�+��:[�5����+��ބ�aJ����9'n�d��E�	 m�$�m�p"��A_��	�[���h��T3���z*O�.ԟ�fr�׺U}�Vg(]�:3s��!��ܫ\��.�|^o4�On��Q�y?(��
��Qx����n�
4�&_>���TୁO���$*ն~�mʱ��w�)�:8�3f���s&����?a���`N�4�hC �\�
���Uڕ>�������F(�L�����^�jr
�n �.]z�@��WY~Yؤ-��W0���&�$G`@���+���fu��)ӊ+{�}�z:���M��f��"%�c(Gf����iD �4���U�lȈn64�?��.6����䯟�����eΑ78U�Z첯����qlv9)�Z�io>�f��/o9���`f�4�-�O5R#�(�$�����m��:�l�\�F�-���& c����ÚsО  =ԻT(R�Bk��EA8T�C�D
Ԁ���ߴ���Mͭ��)�y� �`�'u��U(A���+�:D�*���B7��s�e��N�KwA��z5B�{�,��$�����|�О~�������βp��̠�y�>N��?T���̛^���y���WYB�h�L�S�Np���4�biL�^ ���8/R�t���m��.��>�GN���,��2��[��sE�����p����H��	)���ӡ�Zh�`A-�a����g��3����'���&C_�C����b�օ~u����ڥ�]��jX�D����OVpZ
)����Zs�aOu�A��`�\����aM�x�ھ�8=S�fE4�{&����"�mgh��k��zc-#e�/�x7��S�e�)��{v��gAs�ey� �����o�u�s����CC�]�K�t 
l�2�D�ľ#+m7>�\�؇(\ ���n�<^��D?�L��+أ}jH0Ȇb*�Kǣ\Q���釅���ZA��<g:C*�۳���л�V�I5�)x���`�/��嫛�傖�
��؈��T���������Ѽ"%r�)f����FE^�(Q��蠨�����a
�s��i��7ϙ��՛%�9�ں�z��ن�C_Y�B�_�e&Ϛ1j��Qܘ5u9ru7�uȑ
3��"��@_�1+�~���IC�l���MDJPa����u������L$�_����Y)�����e՚�ot�#B �&`B��D�W���>�c���+�e����zN ?��ts;j�0R�T�R���o���_�����iM�Bքא��:	�`�bz��A֓� 	��1g-�%�����V���'ZAH�PߺU��ް:������WwY��Ȧ�NY\�k��O�y�V6��OR�~b"ŐV��y�O":G��}Zܯ�<�0������}���/���� ��{zK/U�O���b4��?n�W(Z㤆 R*�͈�c�:"c ~FV�t��w�8��<@�c-��!N�v}���@=A����0�V�7e����}�a���!d���h�؝���������;w���b�m�G�8�k�:-j܍i���b�ѫ��=ЈH/�.��������!7���mT����
�|y��˳�Pe�'����'�m!�(�VhG�py#�k��{�������U5DL>�K=��Xr=�D�L",V�"�O-K@q������W�Ջfo]�����6��2Dw�Qв�����@������-G��/������X%&�u�mԛ{���͋\	�/�WP�_�����q�I���Nơ A1*�g���o�9��G��Ҏ�z�j�U�T_�\�Y��Uc��V�.+�""��m�XE
f\CGp@��ܓ��-^b����E�&gf0.�����[-�ȓLPx�U@\b�\��@?{��$E��L�1�y�g���`��d��7lB5� �&N8���Ҩ���J7��]*ۺjv��#����F�䉀��h����9H��İ�����24��sH�k��

�b��w����ց�>ḧ�<Iz�iZ|�ܿ+��ʦ�r@�pu�~*hV���;)�:��������}`�������rA����>H3��X!"�FCb�!��J����1�=�6T5�:�����Ag��I��SPauP�ԥ��ƼR�;	#�;��+.�-�֎ȩ������p�ʤLv�OYL3��K�(��$mW�3��
�@�r|�)�>&�xF�	Г?�?(�hVا�R޹s�67n�?s��w;}��Ά��L5��.yfi���RN!�g�v:­�m�I�d�O�$����V�Ԕ�c>lAڧ˸���*- V�+�q���A�*��	즦f�Ta���|��e�`��V��>�n��r( x�΄�k�_��dr됪t{	��϶��*LU�����VE���f�4�:j��!�0FAWrS�ϡ'�qɩ.��b����H��;A��IC%���dY�L����v�%N�������䔸>�&����L�`�ʰ
d)qJ�b���deyJd���6�|��9�f޺J����zIh+�ERjGR�m�ߺ���Bu:�6�����W��b�kY��(k��B���a�w����B'Y�N�$h�{O=X�(\A"�>�3-�=�uE��o��<�����)�~d����f�H��"_�� %x�Rw�xԛu���(�J\�����|�K�I�v�=+=�|R M|\!�r:+|E�﹁
�
��d1�ؾ�b��r;�մ�.('ގA=��{�D���B�KlZ\j��Т�.��O!(H ��]�,�2\Y���B��yA*Y+�G)���s~�tȑ.���?7_j�l:Qo՚;
�����G@��]w�6\>���>#�����尦yR�o�ÖaQvK�P�?i�j�j�V%��.��	���8�d+8���!��,F�� ��pS@r�α�F�d�!�M�T�h��穙�]Ų�B5Ӳ��0T�����%Ѷ ˛H+���±�����+�X� X��e�l��9�x}n����+���@���������̆6�l��
�b��^����|��"n"S%v���JD��~�)qD�\��}���w�YrN��uco`���GF�	�Qor_\Đ�BB��I��>ja��B�y�)�jo�<��U7���F��n��@�J����ԁƭ+��[Y2jj������!9�f��33?`!��)����S����(V�Z�-�G�n�H�C���_ж��?hE�̾B�M�	!�|�+���)|� o�	�|�p{ħ;��Oi�8��Ofy0/NQ�i�R'Cl�'��J����Rx�Z	r��=�g��g�N�G�3�0�q_in>���u��D�j���X:#jFē=��e�TWou���2�q��i��w� U�xp���Ǯ��x���W&'��.�h�r!���f��I�V<)�S�T姠
^'n���������y���FŐ��`����6�C�wl�a|$!���ғ�-'~V�M�sޏ�_3���ٺ̶� �����X]������i�rƆŎ����q�T�ɣ��,��s2[,��7˸r"C��������ʱ�ԁ	���Iv�1�����l	�u; l�������ЩGh��!�I�磔�ܵ��!j�yR�ml"����;�D]U�/��#�Q��#���fNS.n
A(~/���+j��7Zͧ���O��m"2�7���M�Ru�Ԏn�X6���W�Q�Ӛ3S0U�Z5�R��[M��ջ�y�2&֔)Q>2��P�T]7A�3q�f�j�yw?���b�<X����U��V2z�m��o���/;��H��zE&��p�	O5�z�0�\��ߕq�B��H'����[<׉�7t:i��P�;`�_r��Б bU���F��w�*Q��K�.P��qR .�ֺyRa �����6h�u�ͳW�a<Y�ѵLJhUG��= v�ːĊ��n���v̑K�e��E���_.�Io)���}*�f�R����/Q������@L���G����
��8�߰�~���í<�kP]" 1ݬ���X�29�N	�x*ܽ쀿�U6��<m��t���n��ɍ�!�"7S��Y��k�V����@�
�D���POd�0��'F!��_Ŧà���:��u�M;�*a����e4��'ط3�2�/��$M���Σi�g X^6l��k��؞�T{yqz�A��:@��	d��1��Y��* _.���]�b*m��K�ۚ����{�� R�p��	�]v��X��/������U�� ��Z(�٧A-�ܧ������C��&0ڠ�͏�o��	�pGg>�����X1��!�W�Ц`�y0I)�{rG�l5�wʵcW>/��F�Xu�����x�e���}<�K�&K�<oQ��ʜR/�h�Ɵ�'��I�����S'�.���u�2�UwC���B���ߎæp��OSw䚵[d��4�=Dyå�.�s��?Lb2/�u
q�Ɂ&�|Y��uD����:#ǉ�=`k��V�.�;r�@�-�Ԙ����S4C�^�pT�������dh)��Ul��<8��:`�ĸG�}�0�Q��TO]bZ���#Q�ɌdB���Ēx���i��4�ji��5��E�&����m"���"�B5�o�Pz%�^|7��-��˰S��NЍ\���$x��Y1p����P�z�_�-o�jt�<=��V�QT�T��w�m�Y�e�+��7`DyX��	*��4@Z��	���R�+�h�l"���*,���#��J�>!"_�FQp��+/�B[T��nq9�5(�t����,Ƭt�ft�#��#}\:����+��� �;��r����Z�S䉍[ͱ}����n/M����_.�/������@�9�S�>���-���P��:�zU��h�O{5'�&Ӏ��F�\��K*��&�w�C-2�{	v��H7m���� #�������H��Vk��o����@R�+h�(3�Q'[�ʳ2���[�L��H�F9��C��p��:��K\r���>Id�����a?h�=NB?&�e�4�l[):C�*�, �Ց���ӎ_s i�Z�%�G/%	$˄M݇�,���:���!���,�?��-*JL�I�ص�1_;NO� �A��3t[����1ؼqv��1K=�2m�#�_�N�j�@��=O'�ump�>)K�H�3z7o�J��>�員�/	̻�E'�9�|���.�E6&TbA$�(���n���ǿ3�:��B������ֶ�̍4,Es@�Sʉ��B�i��6�< ��0�Z8е���:����'�82���۞��ْ=8%wd<{���Q�ܹ�
1-q`1UA2�-��8�W�����w\��;ͬ�T�u��ɹVg����iP�iZ?V��,�Ľ��L����KJ�L�V��#�����wR,�MX�`�2
����$��ĥ����(��PN�}༼"V9mrQ��9�iM��p�V�8�Cnx�~����ީ@�`rJ�o/�H�ھ��dˮ���뷩FF║�F�U�ST\�R)�����w�V�اe�"�A4=Y�<Wn@���*��{���r��6���9 �1ۣ��A{Y�]GF����-�!�I�,"�;��E�p:-띶��(Q��8�������F�:���sy�~Fhb2O&�$3��;X�^����G6ս_�# ;4�0x��de�I-�YN[���)&Z_�Ɨ�r�%�����_q��9f��Jǚ&���*U;i�&Lq����u}M ����i3(W��!�ee��=��K �f�ya�/	���	�;�G���-e\�&��hb݀d^ӵ�ş^ز�[C
��%����Wy�M;-��6�NM���#�',��.s��a���1Y\�]o�/y�w�q�1�o�ruS�U:/ql�5mz�}6��7B-�C0|�Wvp\��'�|�#�A&j��S�b��̓˹�����I_������r}_p��G��{�p��E�O�F-�^3��~�J�X^��lZe�n0����;��rTwt�7.���?�Z��y�k�����M�5��E�C�-{c;x1G%��]>��������.�'2[b ���$,���~!Ap�bY�:�h����a�Pcr�"p%O۵�9��HY�鰽:6%(��:Q�tg�/ x�`�Ǌ�^p���Cd��-x�܊������]��h���Lc��j�F����x��o�T3"[`���Kw��H��ޮ�ܞm��M�~	ꄬ1����Ν�� �Y��zϲ�Po���V[�3�&�!�;�����������<��>���륷c��C�X� vON���*C�0�a��*�T�L-����f�/�׿�ƺ�O�q���o�c�-��l�<��`eO��;�*��2�S�Zu��UDQw�Y)�Px�����?7���C�>�U2�k��W��8���
N���E��5*t�^ ��������n%gbXU�c�"�Uݬ�RP&�l[>���z�H_W���eC�jʼ�tD�6"��?����j�X�о�P��k�w}����>b�Mg��.a�NA=�i*�Un�1Љz*q�LC����]�Ct�/,g@׵��v%(��&��6�~~�\K�bF�fO�k�w�����o�C�xzcB�q�9o�xD���ep�]��|n�F�	�����k(���i�j|5��%L�5\-�\�u<����O= �`t/�R}���Q1�i	��l����e43���^EtlpC�@�^T6�tD3�&<�"��t��V�	o������&������9�[�7=�~��uht@�y�']�B~����-wt���c�ޚ[����c;�0+�����Le�&�&b���5�4J�gٚ|�,#b؃��!iuUr�s��y�\#)JL��
$3�K�I9�=k\
��^�|�I�Rv|B��E�Ӑ�m4�L��hg^�Zt6�Й'��-�� �ᑰ�/+�+�a�{��3����;��Z}�@# �_����M��T7��/Q�["jp�N:�>Φ8�f|�%b�N�1����V�э;)�뮥��4�m�e�[(�K�������A�b����0��q��=��v�ӝ¸��4�T��)�Ŕ@��? �uCw� ��eiTi���!�&���W�`6o[z�쏍M3ay<��JL`2K_I^r�Ѧ��y��F2�}�ɾ�JqFCˋl;�gL�G��7�op����oJ�<�ҡ�,��<������+N�"R��6�������#����TT�����l����)����>��ܼ�������Eû	�����l�����`c�vƥ+W�7��X����/Rg?�R/����C!J�_]�Z��X8[-27��<�9�﹂L?TPj�[c�]�Gw���OB�p<�U������d1��$�Z�}���I�����N�_��,$���:ƺր� �Q��Kځh��)$�!zogG/���'B���l� ��O���\������>�b
Op���3�Ý�Q��(�{<�b��:�y��؞jh�����d���U�?'�=`s�l��D�7��=��QE�壴�2ʙr^-��!BS�@'��Dl�C�YG@|�)R:�x_._��1z��^��H���?��(���(@�'����H�
p�����v���;����<��v��3���fCת �>�4߻δ��rI���xnv �����q���ve_d:�h�7����gw�n� ��W0?a��\u���#���|����SZ�~O�Á�}�<5x���iq��G�������U��9���������LǼ]�T��D�W":�"�U��@8���cU<T��" ohj�d���P�g�Y؄$} �[#�#���Gޥ��n�!�𞥱r_[BiCU��ģ��9�4�x�x�*B���jX���w�/B:Ք��<�"%�T�C�b?��\t�=)�Ǟ˩�ϥ���^:|l�X�a!�R�ܰ#^1�v���Of�x��߭�i	��79�#����g��R�=���Tj�T:����H�v���4�J��[
E����O�m�)�
B��CU��:TzG�?��/W�Qm.$]�Y�gr��҅���`;绿;��(�뙽7(��A�5��*�=���<�D��Y�|��`��ԁ�j6_.j�<���8������V	�l,�&i������RC�y�'��7S͠�gM��`�� ���=P	���yP� V���"t��
4ć��K���L����?a+��?�R�Z/�}�3 pj{�*`"��p�R#E�$��Z�B�0�0�0���2��8�lgg�6q	��t�m�Z~��:j�e0�6:�,���`1�q�dET��3���l#�Z�ߧ����>�8T,�{ܤ�1#ṷ�T�|�򮴺JNղ��Ĕ�\l↿e�O>��%h���<(������@����C���%����'P`�o�]<?6 �:�o��$�7�1����>-��%dUm��E�1��Q��~=vJ�c�[Z9R��r�U�$'^���O#��NH��UH�0����Ztr`�����#�~�Z�~����2�W0}�]�3�R�3���|7:{^R�6�����������~6����ִ 5�4�"ħ��P��a\�G��]���J�x�e����Ki~i��Ʀ���`�7^Qm�>���Ƥ�&������XW[c-rXtWJ�2�X�i��%�DHWj����5�|XK.@������$�E�u:+�vw#!���}�(��D��H��[fv�����in���k���rj4�
�n5�W�m�������3�@d����,��ޣ}�(��;����?g���"fV��iK����ݾ`8[P� �\��nH�5���֐�oa���g����`�Y����|�\���0xF\lO�����K2���Ե��Vp�&3�RI�x�D]��X�:s������\ܽgz��]Y�g�8��P]�~a1b�P�\��y���eQ?���:�2wu ��"�ϓ��Wb����]����Ё��"C�d��5�T��� �c�����*Q��1*˂h�����^����%�����&
ŗ�M�����[�A�ʕ�C����ڸ������By�M��O�7��V�S�M}���N)��tz!����Q��Ys�h�s��~���X,JX��av�{Ld0~�0���'Q�V� 2��tzB���8-�̇�����o$���q��ص��áMj��+�d/017Æ�w޲s���8�	yb����:\����!M���*�$c�'Yt��&����������:������;��&��nЇ~�܎fg�ۊӂ���M�ʇ��P��~�ɧ�G,�+�y@evG.!�ҙ�5>���Ҋ"�byEJF�D�Z�X��|�Y���q�1�TM�>Z���}^Vn���TO�PJ���.�X� ܌Kpx&����]�$S�l� �bf�&�҅��_y�@I�Y��Y�Wc�s��Y
���tc��]�Gr���Ԕ�9����]Y6�Ck����ӗ(hbgG�>����q��u<�~�u�������l�o��E�+7�j#Ƙ��/e��?���$�h.��v��DjǇ��Ы��#�-�aXl׫s��>YM� �d��V�k�3G���_��2���_�.r㮠�O����6W��.�T�b߻��������2pT#z�0*�3�0aٙ�C��-������K_	�Fك��!v���ŏ��~=�i��^��@f����9?ʃ�(f(7+�}��n����X��9@Ok@lGx�ebI9ؚ�S��[���s9و����y�N�Z��ۓD����N�#Ll�;�6}x�$�8����2��
��*���6�z���;F��M��RU9luM���l`��5��/b�7H��X9xs�x�ƶuUD`�/��
�~�E-�I6l��:�u�F����Go�� 9�'U�[�-qZ�\�-�s�C��~��	��z����s��)K���)\!v�׵C_�~�`�"�"r�
�Qk]�[�v���D�NK�%7j�`���ȡ�%�̮�����]cS� ������52xAw]�"�o)�f�XH�l@����T�vN�'��A��f���!DjX�8�k�񍧟XK��k�C).�������PM2�<t���=*ߟu
��+k�^��;�� ?Æ�<6a������D�.4�W5ěvS�PL�y���[�4�g'��Ϯ񪽙�4�]�~ڂV|
c�
A�\��e��y�
�~$��`C�[@6�S9oc���eQHs� ���֐������s{�s%��������dM�BU�i���Ƿ�nr�6ޮ�^}K@�5H ���2�<����	���.K0k�}tpG`����:�����w,�n�0jJԥ��ˈ<g'B#��;)t`����*�|�:�ޥA'GeӋ�h�|ߌ�Wّj�c0UPgno�z�-X	�G�k7R�=��Ղ�m�(�@M8�H�m�g�%LU�֍ĉ���N�]�z��J���j��'�<�t�T���#G����[+�X�cɯ7$��ʇX�(�-9�������Q-��	#�6�o����1��M90g���Һ�&���!�J�uD�ʶ�?��m#�i�I�p��wK7�8a�][�!_�����d��H۩�0m��&��9fRz'i�r�t2q)�c���l��t�扂Taү1բÙ8I4���ɡ|����]�������	;D�^���	WB�^�Ż�23����Z0������U�����j��C6�ў�)1[�rN�^3oy5H��ŝ�I��WCDKT�Hj4�b�p�����Ze ���3�M�=�о�R(��1x��m��R���a$��ת�j�l��@�|.���� H��4�e�	5�;Ƒ��J�O��u���l��X��ڀ`Fq���<~�O�F�]6|�O�%c���B��}�Q��p�D'�x��Y�g��x������G$�Y��)UdWh��V��O��5��� G�h�ș���@��Y)�����˃{�T{�)��HQ�A
������a K�R,��I�.(�Jp�@����6��5�Io���ɴme�)�t�ւ�>�)Gfm���r�h�Htyz@��7�����4�P�� �>�Ѩ�B�`l]�?�$�����0�|R9]Ie�Z��f;�CX���=��,�M�?t��N�p����-�[����:�~�{�WG�K��j
���s��l��a�a;>u���9�[FBĎ��{�}���?J`W҄��U|��EC���Ġ!,o���}y?�4\�♔�!#{a�엟�כtq����n�վK\�bLyua��?�1}�͘DS��p�~ܒz��[�*�����/i�EU�~r�����z7�����:Uv�SȻ��pe�(X~^K9��Q�����)+�+!b����7�(F���g8��V�����N�:�u.t�(�y�����{�I!8H�U,���H�+��<����Y X�ǃ�~������P�|s��p�tw�@�Ws!4e��H3q���l�7�G�jE"z���-����)�m�d	߃���+t!6a�-��)��n�x�-7/`6x�ev�H
��C������2����}C��I,ZY�"�[,:�Z�QBK�Z�٩�a�#��&�\a����~.436��A�>9����w�1���%��b�8�7aL��5�)b��*���9a���m���N�q�;7Rp�l���P؛ŴEL�e��S҅���c>�ji]��k�'��T���.���p��A��昋�G���l�q��aK�U�<*�SM-ź�U�C�q���am'U�u]&9�٣l�������w������|��"ϡ�2s۞�s?/�N���p'�i�"Ɯ%�}�����T�~� �*ÙLm���1L��La&�h��ʡ	�M%�o<��M�fe��x�i�L��&�����;���C})����r�U�?��e�����E�&��.�Ay���(��Of�=ۇ����,=\����{��c������],j@�9��g��Q��%Ӫ�D6��K_���̀��s�)>��kQ>��2O7PsY��1���m�hm])͔P	�` `���3'�-1�]���뵳M�}�����h�bf���:����O2�yC[N<���Q��9�����4��ͧ�䪲�
E�[�����*���)���Ա/���k
?�*k��S��Xc�@��N�G���*�����	i�JgH�s헟S0�\�1`L�(krN^��'	���i�,\����+�ޘJ�i�P�4�x@�ka��w!kbc������Ɵ3�&���m�]w�i�/��^�u���t.��\yj���N�)鋔�}������e*��5z�`4�%
{�Ndj��'thOP�*,׊P�$��E�ᖶG�"S�eQUJ5�U��tn�/C��	�m��B'���;6�o_:}�9牘~���p�X1�i�8���\�5�v��3���;QЋ�.��(uPJN��8}��=!^K��!aq H�;���d��qz3,�c3���z�"��:Z��)�l��a.�iɅ�Lo���(9���s��.����Rl��j	xi
k?����|7"�xdT��(J��PID�B��zA���R��; �Y�<��צպ';��W,�#A���t�M�.�(�=$�QT�b��X��>�N{و �4� �u3�K��|��^�kwԵ=/��O���i���q�lvo�'�}X��_�J���E46K��?d@F�y���TV�7=��h���8~<L�$U_����(��bӝ�W �����y�����,UU��(TE�~��� k��bm��?^��"��ӭ'p�	i6-9 �qF�WZ��~���.ۑ�>.z��^1�X>-��e5'�o�j����U���Z�q{Y� ��]�{�X���c!�El�*��(�&��%p����ZH��iˬ���£p;�% ����#F�&<���q���f�����P�dV�ߛt3uhoe��E���=�����h�����m�"�s����B�}�S"�v4AR�ʘ
[/� v���������:�h��� 6<S̢Uz�kz>g\�w��Kd驫�rcDD�Gu|�D��e?DT�T�JOt59�|�J�@�=�p.�ɜ���D��3�ܴm�z�X;��m��U�'{�m�2\��#�調�d���!R����c�|A��T��ap�DGP󜚻p��d�ӷs����]��a>$':&� RH>�fz�㋧�-?�$"s1KjAE�����Z�:���b��d�2vkM �X����1�m�6�<�~���	R53Q-�V#\���s%��^(����W4�%^%X�"a��kux4�V������'�0~��>��W�Z�7{ax ��@�����H�16b'����2�'�N��.`M-�M�r�w�k�]\7q1��훩FQ������|p�&<�>K���e��L�����ՅݫT�����f;�*?+�:���_�f�Q��5\�l�e��`��h�Jʯ���۶���jw�{+4�,�*��'�҅|�0\��j��n��fG-�3�`��F���N]e3-L�g�"�x��[��[/���|Y�Rۏ�2�Q5샽w ��&_QB`�z�՝��]�Y����mwi?������OAY] �&��Β,�ڔ�����,d�#~_�� �� Ξ��Ԏ���e	��m��S�`E���Ԙn�Ǩr��I'�9"�>���ё�%��w����g��~����n�b:�G%��U~{"���l����+G���0�lAO��N�wJi�[T�u�U�(��l˜rfЖj���=�v���f�T��$��5�nF��,�z�A��dG�j0쐍~p��a4N���ڲ��ob�׬�_q!�)�� ��,y�FdKhLǺ}V�诐�Ԁ�VN�{�"pۅ�J5Dڵ���H|����Q)�R��o�q�$nn�FS�}�B�J��M���u&�o�����!�I(�ab�b��h㗐z� b�
�":�Vg��0����Xg��޴;�	!D���N�KZ�Z�n� Q����U��u큛�{ۑ(�ߜ ���n�ڷ�2c��x�DQ��20�0d���Kt�`�mf
�}reZ�C�|B#�#�������)�vl��=�ی�=��u�p:򦐖kVU�D"o��k�o|Y2���q�1��� q�^�.hC���i��-�[ejm����D#�������������|Y�s9p�f]V��Gi L@���R��{���7��l����S�Ө�K4m1[���%��S�7A�e���ϔʏ1�t?�?f�������`�$l �f��J�ah�{�`P�S�9͡�-�b�-�Պ���:1�1p��M#�i�����a����Ú�����&'���'�ZY�;E�$�;�Zxh�V[�-6{�UO��o�{�X�Z����������\��<�j�R���F�v0�ٖ�wR��n]6�2��d��$�.0�n5Ib�Q엊�[�\aX]�74��_��d�
;���1����f�9���gW �|ѝ��2�����'Qtd�{ �kO�]=�4���|̄am,�"Ұ�P 	�q0��쒆ߛ�ڍ>���Z~�<�/30&�mM3�u�`��I���BYa:C����wUɗ3��|]sY�>�	��K(�e�p����_©���ơ�&���|opP�F�{�kgk��Vߜm1d�|awɹ+��w�Hq���,�Ѥ[A���hV��-xӉ �Rl}���VW��7��5��xeK��}6S'�������Y��6mn:o�?�z�,��]���}q�H���ew�O1\��x�O1���D?��xg��`n�2�F.fZ���R���9�����y��\�9���ҽ����ɛd�\��B!x�A�id�������|R<�gHP@W,����BD�_�5���6Iq�,_��l\��m�N��}��$!�Q�ڻ�a(�[�U9���z��j�>}4�V$����.ܭ�6����J���][kl�D�ldc������V%ɠ���d
��\�K��j�7c�p�I�����b�,n���pT�zϸs^J||���D2o�?���M(����9�.�k�Ss
�$�MB��{�=���Wq=e��y"��о�73�!~�EEG�tOn9��-ܻ��rk�}��ES���dٶ(��[#�Ѡu�������֮�f2}�_N�ܰy������c�`����B���]��!n;Ew�Т�V���e�Ϯ1�.�� u���RH���'�K���AE,�P��	�~�Y��h�Q�9M�����h*�D~� ��d�RزI|kڨ_�O�ۛ����"��rׅ�@Uݭ�`�'�2���4ྏI �iXn+��~f�+�-@l�sd$O��.�� B�R�J!EjRՀ���IΦ����{��1݀((�<���剱�sn�L%P��C!M�z��Ɗ*�O�&���P-&����F�%n��$I	�аyI�>	^e�p}�u�����#�b��a�S�ɍ~��G�&�ϱ2��� i��]�	��h�}O�:�8ܬ�_�+���F�h�Z�RI�LW,���������ʭ����	z"������k�����s 6B"J�� �z�����j�����IMDü����8��Zn��9�� \S	��(����l<�pe�ƥ	�Zz�J=�u��xP���9�!7�h��@�������� 	H
�s�D!�5�v���S����a.ti������x���Ի���nD}����<Q���PI9�vlȔǥ���1%�qAu�w(fW�`l�����N�1>A.����B9k!�8~oA��U�_?=円�@��F���=�|�ڧ�����M��Y�4�7F*ڒ$c.�-�q	B����� 9�ߙ������y�s¿���L���]�Y#���^�/���L��'ۺ�8�D���'�~� ?�NY�P)E��?��eS����]�88�TjVc���D2�ߣ"xE2�rI�\�ۏ��� ��UTkM�wc%�&h�c��1��m�<d���(�Ő��s����R\۝�-7�1�%~"�����Ŧ�����ݢB��u�>�x1�gk�o�+G;v�:�G�?�Q5Y�Tό�{3	v�o9�Q�m��٘6����kC�v��L����S�9��ge$3� $�?��u3j;&J�� ��1�މ�/F��m�)�{���L20��o91�A�F�]�o(���l��v�y(r���˛�s�C\0�M�z���F�����Q����H�,5=l2ɘ��:��̒ wPVh��ڶcn���!��w��0��;�/��50�U\��n6��.�齖����rپ��>o ���˩�"���!��^� O!!��Rk�����a�WZ����~��d|!��R��'<N�m�Ď���Ǻ=H�8���P�c����,4e��$9{�j��Tc߮�cl�w#�!���?���7��>	�'y3�~�=P:$,�����[�\v>�|7 �[8hP��j�o��X�����008LN�}w�pP6>��ȣ�BwGr6�_`H=脴f��¢@L.�mG,/'�zښ�ނ���)-��6�;��#j�X@�?W�D#N�=�GT�VYr�����{.0]K�1��(حڗ\�y=1�L�\���W�JnmU���M�S�ZL?tu�h>/���մ�Ḝ��c�b:6�@�s^�*n�W�w�l� 2Y�3wQ��f��,�7U���8�^G����i�B$I�ƃ8q9���J�����Tm���G�mܳNt$(E����T���M�gE��1�n��9�T�ԃ\tI�,g�20��Le�5�5���Cw��HK�j�2�����h:��ì|��L��7��&d5a �$�R]2T��������%-�0��i}����gζ�� �<G�n��f_�2�,�cc���<���E����+3*��B�oeZ�	��7V�("˗_q\������y�����s�cQ�E��Ң��K�_�fO77�<B��}���s$ �R��g;�7vP<����2/�� �󻽓�w�Rի�o��UY ��Xͤ:��EM6Y�����Uj�c� �)���Ի�
�no?�xIu����\+e��6�zMEYx�����}�+ a�k�V(�N�̐���|O�8�|P>?�㤊��h���AP�A���͇i���3Q���:��	y���Uu�:-p�w�V ��D9��G�E�L��y�Eꕨ�L�{��K�Ԗ5[�K�+afX��~5�y𚸟�!���7���$�Y�9
Yo����5'.��}C&ա�Itk���t���PM+X	Dn�3i8�5�:������0���7wu]|a���ϱ�{�x��8�D��K�Y�J��RBjI#���$REՎ���m/_���+O����}�;�Z%#U�=�7��������*-��xS��pߘf�W���	2!� �S�^��66R���W�0�'��~%��OpR��3�sG�z��m��,{���V�O���v�nfU�:�ˎ�n�f��b]`��?z�[���YV����B�j��n�Ů���1Pe[����W'͸�����Y7C�+�n�Zd
���\�����ӗ����Yr�Ie��a�m����p���_�w���M6/��F�O�������_$��bO�󀿭q�n���d�r@lrlB9�	a�_�ye��8�+��$O�N�5�8x�k�%��K�36���W�:�i�����3�Z\�R$�S]���'�ۀ���=?�
�FD�f�n$U�� 7�ݥßF��������Aj����B�p���f?��Aw�;:��J}�qQ��Y�J~$,E��k[#"m���E-ݐ���l3�;��[�Za��'��z�I�>Ҁ1�I�N�E1��]�W�F㹔ʻ�oǈ�<�ѧ͟�H�.=��X�Ccͬj��wK�C�� �G����|XqY������0:��]�`��W�-O{�i\^�n;[�����K��2���A;C��|~^�~���T���N2�^�R��)E'4�7��whn�A�[�?:p}&xb�o�F"�r|�p��Y{�	�3M�*c�{#M'�vY�8��g'��5Z����?��oq�q���?�@��ntOq���>~Us0e�:���i��b��	[Y
 ��z&��e,$Lx�F\�y�y�����C�Q+R}��|�4$�w끫f_nTK�s��o��E.���j��c�d#ݭ�bQ\�ōV��u4<:VG�.K� ,ay����h����Q��� �fN�Q�֦t���e+�%6�	��g�g�J�%��SZ�83rʠ�m�A?�z�)�aԥ�A5�BL��c���0Uw
A��e��׬�h��l?��>�"��ѧ�6��x4;�����o�� ���'vX�#���r%�	�� =���(��:��R��l�O�!`q�jk4��3�[-I5��~n�����2!A����Uua�&����e���6����t;rO�����D h"`�݆��|Մ����|9F�G��R��sjs2��u8 ��'l6�(v>����_�>��SZ��i�01��ƣ�s���@��p�l2�@�T �vLN`K���������w*��Ǧ�IX�@9�6�Ś^�G�:p�iXh���i{;�zRm �1H������/��"u*��n �:f��A7AR{����j���8X�a��A�������y�&[$y��wǔ�?�.��K+Ǒڬ뽨�>äBs/��(j�y���1�
��!x� ,MIiLr&<i�榞�q�,�W�"'�6�}79T�D3r��~R�r�W*d�S�������R�i5�g5�j��i�/���ۀf��k�cЧ�� �v?w,��r_�yÏX��C��=�L;{��%�^��|��دr�b}T�U��`^Q_��d��A��x*:��\����d����"��#(��8���n�UQ��@��G�}�T�%AY{�ͮf���x_|X��>FN��HpKb6٠���m�.�1��xD�i7̢g�Eo�	�� ����_�d^l�O���ƶNez��v�}�
���.1��[�lԸ�MwpOe�e��	iI�V�{�i�O���5�L�-�X���+{GP7�&c�$��7�C;0c��a�<��7��!�[�u�����|�`���K�@Bq��L�\n����1���zȦ=A�'�)!��,�W}�9;5�W��D��h	Φ]�?(
2�'�,�{E���[�E]
i�u߳�ogX6��H��%T�X��z�7�C3��Lo������z�/���rU�'��Ԕ�ia�~
��DW�ֈ�r�L�2(��{\K;�,����q<\���Ǝ9֎ǅ���ﰿ0.&������d����HYW�}ǥ��oBax�O��k�ÊIH�W�c�^H���n���a�����Đz��,���;+��p_�pR���Q1tH�Ѵ������l��#o��C:��������BW�"��B'�p���?_��)��H�\$R��JPL�,���)H�����!V1��x�%��PM�(i��I�) �4�"�8"�;�m�vF~�;~�T�ڶ%��0�K�j��^��.�%觴4^=����F�t�g�v�c�fm[{J�1K'y�<�C�uI%h3�kkƭSkT�ZZhd1a~U��֚C���Ό6	;Ģ�*��v 8N�W���g�I\Evw��5���=�		�[�\frq�WuOqN�uGA��Yh�]��3���*�]�J"�/�N��P�SkE�1�M �����Gp=+�G���dx�����J)P�@寵��x���	:��g7�P�T�Zdg�U����KunoD�f��H��Q��S��Ț�~�k��3��E��r��v��:'�<c�`�f�����g�A#�X�0ʨ~J�-Ԯ�
3�K�DCb�7!�}YB�a�9Gc[P���9�u��)KXK���t:��4eC�q�Ϟ~o�
G��&�ʚ�
{
��k�f�>O<R��7�^2���[oM�����6:?�yi�)�����K����DR�ю|���=k�~�<��ۀ������21��ݐ��,�ٲc3я�m���Һ���l=��,�g�6c��7/o@����<ܜ��wea��awH�CIZC���W�G�5��.���t�L��>K��ic��;�!��h��w��H�	�)D��|��Umn��a0۾�?cJo��7��K�>%���wJ	x��iR�.0�(ظ� y��K�A��D�x0��'��h�)K�0��s�e7(����]�q��[�%�XJC�;��� ����P�ʡ�I���7�[�B�i� �yn�#����j����s)� ����SK�v7]��i~ȅ��|�f�5ĐZ����w��nlVR��]�����w��mW}�9B�9�(��%u������I�+K�i��Ա��
���+~Ys�#Gj��� 0�<dB	�\��0އx�&�S�ְ9=I(��}��W��t;T1�d�m��ۘ�I/�hF�<��{�ٱd�.Xf)��7d�y�zf
��`�����2@^�����5�r/Tv�C�}���t��Zލ�Nl�-�6wm�J��q���8���!����EĻ5 �%�-;�yV��Rf�V	�����C�%��YKPF�( uV����;3���Z��F>�9NE��-2V7;���|I.L��s��"�49}�ofM$� �e�:��ʲ��.�f_�*�lk2g��2��4��3p�^�����?X.Y�ht�t]����-��y�_G�^A�?��O7<����8� �?Q���pA����#��`$��[M6��:/�y�����Aۑ�`P���<�ʦu�G*���&��*���2�{n�>l�D���<�ҍb����`��<.\�������d�Ѯ_�.	CF�쫫�,I��>����h��l����#.ҟ�l[+x0�q���_�:��e5�L�p��F�.�u��Q^�R�vb�Co�Kd�ir)q��ؖ8T��^���d�q���t7�¼CQ�͍�6�8F�NJ;c'SV��\��v��0�4=�B}8���q�h�J�l�b`�ZQu��t�od�&)ά��|��
 �n"�R�h�a���#��Y<ۥR�ua�r������ak�5b-��R�Wn��3u�S0�v�%"�:�Q��!�E=1C��{��Q�q'^���q�w4ϊsc��� ��0q"�J:�Ćت�hj�2�(/��Xy+�K������o��Hd00���+S�m�^��63��n;�Ϳk'��S}�e�bL���"}�@�R>]���M���ꤙ|wB�,�]�6�Zl����T��/@���V=�TE/�^	Xg�m�W�c��S:i�aFQ�R�Ӡ]%�,.	>�\K3��=�ҫ8�.:~����˥fp^'��G�齩�����7���IYQ;H`j藌Ǣ���ע#V��j۳-��l�s�������	��/�;e#%�;��Ơ�7 ��rB3�ݎ�OO�0�J�i�^u> ��2�:K�T����y�9��o�ڋ�u)���,�@J�7��G�{������~4��v;�j��
�M��X�.v�>��a*�wJ��i	�����l�X�k��j�E|��R��EM�w)�_/]������5�e���N�=���\���R�^�W����%�ٰ���ٻ�{S���5w@�쮎�W8��Q�<����;�\��y��E�m�ē<�����eo�猍z�ߦ��~#E�ǁ4�/����kVV�V��bw7��q[_B��r��ML���RӰ;�OG8m�mspi�U�l�.�w�g�[�H8 os9?����U�i\s�K��}��f^B�b֠��Ҷ$r��GU����T�U�+�@�gD��=��$O�(	���~�	�'��$���s�Q1�cy_"���
W�̾�6Hed�+���݄H8��^r��y��x��Z4���}�x�e �BK����\S$}�L�a�y>Ү
VQ�M��4Qޘ�V}��N���j�?.)^ ]E�'pI��X�k���g,z����_�p�\P��W�bBk��p���D'��,�+T�N�k=�Zc��+���P)l�ɅJ� �#�1]Ӣ*#3ۙ���]���(����?��s<������&�HP�q�˚��6?����#�%�i�3t"�|}�nby�������cU��ɼz_���Fs]ឲ������ztRHc2BE*T����PP0
EE'O(9{�;;Ŀ���)>l�9Okg.�H*瘷�Qܸ������ڙe������,b|e{I����9#UyX�wp�aph�;��7�|��Y�yw1	U���Y�a⎮[Ol��]� ���{��g��t��6�_�T���I����w�t8�/dm�����X�Soje�%6�P�� �C 0pMÒ.0lE+�%n,�<��H��v�"��V=�'�2�I�*� �>O���7lc��~�V�����;*~}�,�mZ�`bX$��c6��m�n/t��U'1U��f�����������0<'K�$bS�:�=�0��Z�|ۆLΆK�t��'�=�ҿ$�]ў�R��$�"a��uߎMgS6��Y���e���/#éV����vis���4�<�X��Q־��Re94$��2���R�	�8�K�3��ic{���HO��M�o�t��Q�D��n0h��V�c\���"��J��5(Z�پu������G�eLỡ�n���eXY�񯿌R�('����b�� ��sTf}�$"���k ��A��Wv���4�nk�`>�_�m��u��^��>Z�l�#�o�5�(k�뒺�Ë���C�hg�% �|���9�|n��f��'~LNx��D"5��4-RS1�Z����#�i�&��	�e��J�<�o�b�RO���t2d	��o�����t���k���`6�޸KS��1O�����������DĢܼ0�ޢj<�\R�~�Ɨ��z5��h�0�6�3�ר���+�_���~paus"}��}�9��i���!>�*r̗�@��J�0ç�5C�f�D���b'cY����q�XbW�o���ax��]#p�]!y�e�}�=7ّ�F@���U0岑Y��b���(C����߷��-�{η��y�bG�v�P�
�� �}����L��P�LWN�O@�r��]s��W�-�?�.���뭏=6�zhP9�}Ѭ�k��$S�����X�ʾ�Fw��UA�h7�C0p�V�U� �{����<C-h4�5���?��wE��C#<����hy��ͩ[a���bUao,0\穴>�\���ĸ���0е���tf��ꚽ+����t_�J���y1��5�?�wh1/}D�v�z�`�����_�H��������|oЅ�A튄����t�	�'T����	��.�v�G^]t�uY_�;6ϻ:��#̾��N!�|�k HA�6$k�5vP̆�鐥d~�^���67_�9�g?:�%=�����Ɛs+�g��yk+ͩ�p���,Zf��3��~�/�=��ֹ>�w���7�	�:�8��b�'�����D>ղ�Qo�e*HV����!���__Т,�H\D�n<zJ��]��q��,�z��P@�6��Z:� �6���/�V��mOP�n��$�`�]w\�4�
�G̉�<NТ=?��| ������#���YI>�ڭ�,�,'�|<�{��7r
�F����]Bģ��iM�������R)� �+M��
���<C!�M�r�/���)u��T�gU�I����iI���R�e�D9�
���g���VЫL���@���˴�j�l��״ִ��_pO6�a(����>oh�]�=�X�і�T!���gH�����&�Tr��`K�.�n6.���{�A��1?�d�qp��9������N�W��rC��H�z�����)�Y�;����-�qj��{+���5,/�����C���5o�,vg�< ����+�#x��+�\��EMXl7����uS����g곋<�l�J4$���0�9��B{H�#�gT�	����B��ψ2��XM���	��{�>h��z������yQX"���J�T�/F����o�0tR��D�5M��#x�3Pm?b��5 �]�~�%�=M��b{v�ah�H)����o ,��R� <�e����K g4x~:�0�ʥ�"t�����KS���-��H2�?�WR�f�tq�;m�݆�d�ך�)x�yUU9��-�xA4�+���*��[&U�0P���8�@7�E������2o!0�������;�d��8ؿ��T3���A �V���>��B�����ޒŞ�%`Qv*6��Za�Jzh�;1������n��:O���E�.�W������˝��PН�##�� �?d�SGI�b��A��  HFbS��~" ���Y���vLlI�ը�k�,>
F�Ӧ!�H�Y!$�Y�@�}}9����j���2(!��|P�`y��DQ�䞻:����Υ'v��v�e�/�ˤzya&q��T*�ᬑ�l
�~��$x[+D~��{C��]I0MA���G��_R�-)��:��B��0-�H�Ԟ�	@�����Q�z�NxZ��է���T��c�I�btd>�j&W�,S��|����TdtL����Y�B�����̺ؖ�2&Z�I����9���(h�����������wd�I�*�Ǫ�Zt�쮾m�u X�N��k�z�S#�=�.p-�$���Xv2߰��H��/<���-�	�Uw�5�)h�嗼�C�0���t�������%Vvp��,*:��=��z�t��LZ��bO����y��J�X��nB-���(L|DF�A:�<{��"I�ݬ�q/A�}\i�&�¼N ��ݛ�ED��ʔ=�� �$VK24�ޢ��$�-���/�( ���ȝ ��c�֤V�����1��~V����Me�7q�m�C�*��mvqWf	�)zeb��2.� o[[�?v��j�&]�4����Q�XxS[��Zʗ���*D�h8��g�
��3�[r����Y�Y6�G��0p�"����������8��ۋ�V����bY���Z���4w7
;fVJ�̑3p���7�/�P:�Wd���@��ǭ��(����)���s���W:��A��tb2Yy��ke�׸ WɛT@[��c�����Y�� ��E
�T�Dꆁ�������W�}F^o9��Ox�/-az;a�5��P�d��ѥ�)��r�7���zI�<*�
������&���90 X�!�˶����$x?%U��H�#=�5--�}��9�o��������d+��fbL�*�-�'6�\�`�o� ��M%�:x;� ⧼&O��Y?�tĤ�yU���D���s��c6��q�S���,}�a3f�!.�f[j
����SR�W�I�Q�k���ނ
�\�Û��{�Ԝ[^�Yq8��-��,�/�ztd8II���0�L�����́r�J����)�����/X�`�>��Gt?_�z�I�[[cr��c)~���5'���e�Y��(��-�2׆B)�9��)T�.�	�t��Y_h�L$=���	��AI�%v]����rS�F���kŶ��Q���3��}��U��t�S�}�=k?�ã1��e��>��ӛURtQ�D�c7qW+ ,6|5����[�.'�u�ߺ��m/� Or !��=R~rH�A�K��#���x���/���+���P�g
�e�}�#���4d�I�r��e�G[h\�����^�={21�X����պpBꁎ�<5���I�nr�.|)kz+�w��h���i
3$��(�!�ktbrN7{�e�N3���ii�l�w�/d��͆�5�d;��ԈX�?�I���L)g�Y�&A�O���I~L��E�� #E��:"�8Yy��;*���E6D����^h���	����`֫x�i��O:��5�Z2i��VzL����a8n@$���=L�#�g@�n��H4�]���F_�f�������g�!�i��� @X`""��Y��W�Ϫ��0N]�b@�����"lh@xcEr��*�U:F�d-�s�X��O���/���:ߙ;3c)u��/@��3�Kj�ͩ
\��n�_	�J��^X>(��i@O�꺐U�K��>:��nY)�<��{��w9�ɀ)�Ӑ-�RI�9xT�eDO�`.R-\peu4�򝊯��IU����koxk���*�i��+΂�F�(V��(<l"\&!�P�}<p����!=��6��>h��WK�~�����<D��	��I3X=�F���=��6=�0�R�4�N!�YL�[�F,7�/V	AZ��.��"!7�u���W�����"Ee��,�?(�,��	08(���_��]{�U��=��$���l*6u���z Z6Z��BU��ʣ*��QB������،��7�p
䷣f��'	��1� �oi�?��r���zT�"�޺秎h�WSY��Tm���>�P���d�㞐֯�2��V������x;�Úu&&�+핖��/�O~�����&c�R���7vUc�HЈ��K(�'��B�ڽ	,�OvMjm�RT������K���%���0�դ~�R0:R�A:�̈�Y�rlIT�[�e;�4�4ʴ�/bɤ��󑙰�G=���߂�e��/����r��c��{.'Nd��dP>��+5r��n���ɲ����Z�����+�����JSs	�b����nyϼ�]��0<a�2٬ÌC�034��E����I���v;�y��f3�%u?��L��a:�n��n���9d���G	���>��M�H�����ԁŐY���Pgt'%z]���bQ����wJ������ǜ���9
��}�	�52'�k�e�ɴY��0�������&>��P�@	`���)hytI�G����=N�B��t���Y�},��'R�����
�89��ɀ�PA��5يP{�"�kE\*Rଙ?6�T�~+��,͠E$�t�q���5q����#b7bƏ��A��1
!����Xlb��u靵�Y��tP8u���'��3��[��Jǀ��Vy�DZ�v�������!���t�M�#\�8�J�#P��� �mb ����*~6��~�U��#Ѵ��'�����F���Y_��"�"������S�Wf��f�ДP��gӿ�X������J<H�ᵏ{"�`K!몬�����uX��2_Ҏ
�,(.Gi�x��=�`�F��&��N�kQ�C*�[p�BR"G���;��Q4�C%)�ƃ�/�\Hl<��1Q���ӿJV�,xb��W�&Ֆ��%����?O�f�	�!ci(��&�+T�8|R�.�8bȧ*��|�~�Ӓ��@��ޱ���\ >х*��5� �= w����~��U�d���٣G\��n�\�j�~���܏z=wy	�
��O@�P�L��~eM�{�ee���x�����w���z$Q��:%�N��֊pH�䊲�8�ւ��:���u��e�.I���P߾�@	�A�	U�k����֛��nu���]�M�QG�u���~��.K�j3��
�Z���<5�8ꎶ�d��A�~�g�eUs7T��q�c�~���.@P(�c,�7N�VW���Mp/Z]�M*?Z�8g+��	�+Z���k�k���X��<�L�9r��gê��i^��{��eC^�M��b�	���A���B�&{+#�<M��'�
׈�(��@�Ail_�F
�vmDb�����_0ՠ55��`S7�&OV�𾼚�G�x�.�\�4i�"�j�5V[!�B�l�����;���x}�Q����:XV�BJX��ل[�>����r����#yd�w�tO�<�n0u� ��_�+[aŚ����mY6r��E�QKMEF%ؙ5�j���O��5w���z�����Q��cVSEńVT��Ӫ��+�{�Ԉ��6^�m��5��E7�A:�5Ԁ�	�s�ڕ Y*�3d���U��o��:Ha�
!T��n��_�0��X�߶���{X�I�?�����ի'2a;w��Ъ�y#/��艪��)GI�J�5Pݚ��sӀ����~�A��#`z%���E���E ��+RZIc����S�v����^�$dE��Ŀ��ΣB@�X� d�xWi�4$'i���'���	<J��Ji�i�y�7��Px5�"�rZ�0LB�Z@.�i>.5��c����P�a�<�œeky/�}�zc:1��g��J�ݏ����}-$��e����[Q�ʤ"u �Gl|�c�Fɲ|�<�=����<H]9X/swH<K�F>���<kG�<��'�F����U�����[�؊��
'FW{����AT�2��/�F/���0�M��B�#R�����󲸾B��A��&�*fcjh]�	vj20D����3:e<�Nl�ߪy�F��X�lq?���o�Wo*z�
��H��v�c�m���$z��(|	 >�#:�/g�������꼽~*.��A����1��Fa�]��R�|2�QG�UI������F(9�B�3�������E=��ҽ�i��{	���Ct�˗MtN�w/l�7���lϣ~�[�?���`	��b��8����]LG$������4�i��v��H��AI���z������j�7W���}per�
G�U]��(�4�O������g��O;��0�~�̥���_�:Q�[xs�(�Y��Hk�@LPl�卲rHR0u'?�j�ݝ�|%@02 ��nN�h��~�"��2��=� �4Wtw���]@��H��rf����n�nZe\�w���FE��8C���Q�qӼ����i�F#���Ǎ���Hv���������(P� /�Hf3|�C�w����:n��Ǒ�� �q�~KS�Z� ��.������)<���xƆ0x�#�Ϡ�؂�X��9�'#��l��n4zkܛ���J>я;j��W}g	>�o�)P����bW�+<���?���A�1TC�����l`�+N�>���ƣ�;��3p&��~����>�� G�_S�AlH������TĞI\>��_dǛ�U*�f����|�:�cM&cOQ�j��mԨ�>�"v����tx���
�����	߭dE�J�8B����b�l�3͙�l���֋@W{��+3�gZ��НH
!I��n��c]j$��c��Ů-�"��`f���W�U��pOb�ې�}'#��Z��x��0# ��Sm*�U��b|�k�����:��!+yt�Â�B�>�͍��o�^f�.�2ʙ�p&����+��ُbqpd+�}�U�S��{��II�F�`.�x��Sd�󳸙�`b`�1���˓A�^����:���p�)&Q�,݉��є� ]����z5Z�k�s;ͼ��[#��Q�eP$E!D�z������p���Ӟ���!����g���9��ME�|�c$����~ �w ��P���ڎs��ID<��Ήf�����FF�A�N2*G��]�8�\"��0_���H�8i��,=T�-�k�s�좜"��6Dz�v�ܴBD9B��Y�N������=k�z�)����
[e��@��氟�t����c����3�`҅�dqu)r��`9i�|�Đ�x�<Nڑ�S��2n2.@"UvυT���5^�&l�{�U�e��Aj��'�h�O��h���/�I g�
'@(�趰&�MG�O��2n ��+|tA�R��t�RJ��DLu�#�8Kp����U x�J�'�*����ͯ���m,��m
Va�	�-{/�݈@��d�'�Ua�v]�J	H BQ��܈H�/� M�v��S% �iFг�ef����!l/���C�>���II���3��E.�~����uf�F�F�����Z�E��s����AO�q��\���Á40I��h��t�4�{�j�=�OsV�s��4�Oi�.Ȉ1D���?�|�ts/���RS�Va��K�k�Q�[8����E���8����cL٭�ٿ��֌RH�d��������.��+��U�{x�b��_�	���H�vٕ�Ǳę>��������Ap��S�X����]����1�l�P��+:��4;�����_����G�[E�����}�]	�Va:���Y��u����lE�B:F��|Dʫ��A0�e��J�'@I��U�$JB�t��"|�����b<4�Ѵ_+��������A`zA�>���hc=ѽmO
���*��ys �D̬���9ۋ�!�6ˑ���Fe�J�85�ɸ%5J��{(����/u0'8և� �L��^��o����C�A��3�"
��fĵ`\T�ťkf+"�,�f�'�f����l����:�!���T�=�Y�|�(qȭ1�/Б�y�>Q�.i�R#���[q6����g�2c�ʵ�>S7��񐪶ͨ�������4e fv^<cW�#�n��6��紒Jgִ���34_�^H+�k�9#�+e1e�ܳās�P��,Јu͓N� {��a�c�|��3���-5��������PPq.w�'4P(p	;T�b���1j����5�?4>rz0�DHh�='�ƀ�O�練28���G²I����AeH�t`�t���B[�0�9$.���+�/Fd8�!�1�y5LUͽ~p�݃I�|��
ےRP���h��ܧY-����{�/	��'��gB����
S�O6c}���}��W���/ܱÇH�JR6���G�-7l�x�N���>�L�pE���ށ��zD/�Z��P'����1T�A��^�I��dgXf�����b����f���9|�h�m.
�9���P���w�{��O�Ƨ�mD�[�
�X��z�=r��&���2}����ɉl�̈Mf`5k�`Z2#4���M-���Sֈ��\�&x��-W����I�?"�T��u߄Lڙ����i�x׾�����^��l3���=�DIE�R�=@�u@a.�Vz׮.�}�)���}6浹�hX!5D������*���(������bf�>*�+�r�`xCA?D���k1�Os'����tӢ��������T�θ�:���q�,�}�g��-|Ex�_�W+d��< 
�uĵg�Z<j�\r�f�Yn�p0�q��Gs6#�RxYN�����צ�wE	/)��3���)7��8&�3��|"�ܘ3%(�RM�����<h�s��z�S�3G�!���)�� k���a�~Z�AJ��7�3cq�k�@��/I�6�qH*�=Oy��N�Q���SQG�����ln7g��{���qw�!�~{��ENvE����SCR:1<��
݌������щ�4D=�ˁ���'Ed��9���RC��������Y_���H��<���6]XK�m|-�jfxnm����JMw\�͇�j��l\Bs��`���6w5�� �"%��9*"��1_
*�g�y��`��D�a4��nN�ĳP���P����Y�E��tzx��-V�1F�I�7>*���0��ۗH0��6&٬�H�N�#sn\���)�~���M����g�_p)Dّ�!|]l�g�#R�TtO�$�/��?"5�?v*���J����F����P��ジ��%�����f�ڒ
�~Q��4l^�y�Q�Qkv�ю@(�����oi�\�`�u(�-��/q������ch��� <��VB?�Kڅ����Pƙ%;S>���ZS��&R���/Z`�I]$p�e�_NU��q}���{vp�������р�� ���.�,����롌��`-�EO!S�֑����w�E����[ҵE�^�6����'E`b�
�c��w��SoL�Q%kV.�|>�噳��\��9xڔV���"%���ߙ!���9' H������#ŵf��k)b�f]B�'M��h��-�AjP��&]��}�)"����X�J�WQ������;��
$�{g�"~�*;Ro��D]���ҥ`���}��j��A����8^Bk-_d�o�ފ7Ƿ>'L�;ȅ�z���ĕ2�/�,75@��DD [%Ƒl<��`.���@jY�B�s��qIZ���G�ae�^�������zM8�VwO����k��K�!x&D<scR�Gl���-�(�f����9,s-���eFlj�5�E��c����K�J�ۮ��)�����6��bP�X�8]��q9qy�����М$?*ɻUv�霎�u��ȧ�(�%v�=�r�A�Q������|%�
��/��WX�_]2�
3������%����]���$;/Pۘ9������3���Ð"���w��Ey�B�]���9��
^r���*jȦ�Ip��=R��rW��^C ?V٘ؔ�bX�X)�������_���8Kg1�zRAJϣ��/r��ľ|�6��X����1ݸ���E��(�S�t2�<uy�jclڮM��(A0�����7z�'}Nu�tt(�9x�Z\�ܱX8��.�UF/���:�Ղ՜L� ([Jm<�*�A��?9����w�\����2��gGVx f�|�-�R��y��O_��-��ȕn�ůg=Y��Z�.�ZL61oſ����H� ���\`����ئU�i#���X^-A�BS]�cw*���8u�.�@���Q�U<^�F��h�>�/@!�i@�� ��e`���1?��˷.\!��[xC�#o��������&���w�R�I��zzq6H
��N���T�ܗy�|��~@Z�u��|>�z5&�1���.��-}�r�-�Fz&8�#u!\8f�I��<�1.^ϳz���(�++cMה�qǡ�40q>����
���X���#4i{� ����_~���?�D��:m~����{���*q�Zb�	U胗j,϶��D���������}��)���LF�;s��9�o �M:�_��]��'���>���@��D�(Š!G�^��F�i�+������F
��(�	�w�d	��'��@2B&�O��#\�?A0l���f��2	�H��t��֦�������M���I<:u)�vSʏw��z&!���:6�+�{�9�>7�%�m��y�����X��0��W��4�<W�0Yp�ҸK`�����ih��_o3��;^р�5�ԭ)�|���IL~ ^�"�ݦמg�o�a͌��]6/~�:�;�dd���}�Ԧ��3��jp����w��<e_�(z4���=�c���u{��}0��JË��յ{�;[Kn����]"��bq��zn�=_S	M^c��<���G�
�ȤT�����.��(�߰��#��M��+��st�E[VЄ����˪c�'*𾝠b������5_����!A���������O���$u��5�e�x�n|���1}�0_���ں�A�P~�@P%��Cdu
�M�n�.�r�|����ZLm|;��z2�2�"o69@�$V�`�T1����P���+�{��M-�s�)0uΪ��:ͤ=�;�&��/�F��u#��V�A{���Wk�v�����Tz@�U*�E"B�Y��y�~�%L�E����{A�
�����k��~�
�� Ƈ���=-y����<�p�u�X����8�pM�x�p�tpw����:[� m�AI�̚�����i`a��}L�\F�g�D[�7l���|�-wR~��N:P�n����ˉ5ue]H�%F$@!p_��>h���cbC�3�K��~u1n���>���n&���݌��\�j�Ŷ���������χ��Q���PMZ�3\�3[*��J���U}��W�Ң�����&�׵6�;�X��T�W#{��-��4}�����pj���*�r-�H�!+ͼ����Ȑf���KZ*�}FS����zo0���W#-2%�w�3�P��g^
0�w�i�� ��d��ƶt�,`��o�$�ؽYzв{�4��R�,��"K��e��&tV�Ɇ�BZA>��Ud�>,H���MDߛ�uC����҇��&^�J*�s5�� 虚�`�A��=༒-6�l�uG��l�&�M�)�"E�Rz"��q�ln1`��H�[�.�md!oVp��B^�R��M?�i���~NB�a���6s�ˣ��4C9��P����t󰎰a���2=��Ի��<��v+~�F0����H�@N� �JF�	]�r���ͫ&�5I�U�UkE��x���Y��Aɑ�����e��q�O��A�6�9)�P\L����>��N���I��"Jj�18�b�?�U�2J�[�N��i��(a6��4�$�Eze�V���ޗ�"�^xWI�J�Ƀ�S��y���*�!Ӌ=����i�LG8$���32�Z���L�9����hBǞ�M����n�-����~N�"T��[�b��_�0�ذ� cn�&�$/M�7��<��Z>�������wN/m=L�,g*}̇YJw���g�JQ��{��cG2ky� ��ݭ3�R��a<��,a!?]l������ϰ:5<�To�����}n1����5�I^�(�LK�cz� �ᵲZ��Gn;w�P�&X	���o��q �)�}@G�}�لA��^E�ZB���!��t��ԑ�(��T"j�,H�	�z�j��~��������O�jy��G-"M��E��G�%|����=/�S���]^�I*(��
�)+���A�t�4�׹�k���z��tn�=7��r�X߯M�"jd����6x�BX�K�(�~*߾#��Nd5�M%�}!���|1r�n!I@�$�h'A�a��K�v�ܕB�9of��?C��"eSq\�r7aTp��勞=��;^S����r�!O�7�æI�j���T�L* Ԟ�+��ε��c��.�%<4�3���V!�M�v�Q�Qp�
��O�^Z�5�W����<DJ�p�,i�	1�X�J����'#��mX@��^d����0oQ��
�#�{�-(���Ml�Pm!j	2P�]^L�CVj�%��no�hŐT��p��:r՚A�eC�vG�����~iZ�!�w� ,t��yן�w��I���U��M\����H&���Z�
)ˎ�=啔������/h���n�W��hA���,Op[,C�������k2*$���aR�S� �Y�/�Y`b��\,�T��̐�bJٟ��B�z#LŢ�S�{U��<<�ì8����'��`�zP@���FV�Y��/ԯ��K���tl�r�
+y>&�����N��Vf�ϿJF�y���+0
皌�}�N�v��I����B�@�m�	,2�{�뱛��YC{��4��q������%����-oҼ�LL~�?�ùE%�@�V3�@|��/�D���:ְE���H����'�2��]�ygA���VZ?����]��U��g
V�߅"H��i���qP*��o�Y6��ݸ�rb�RCh0<�|Mcz ��`�ᙔ"�CS7`5�"��D��Q��߰UdO�IC�2(���4o<�h�n+"
%y�m�Eyk.~��Z��S���}}E�D�o���Gm�+��8�,04�I%�u\�P�h=;/T�l�������­<�˕T�+9��L,Ӭw �[��xR��X�i=rgse�IO_�a`�0���kd�s*�o�(� p[� l�)A��ڕ��@�p�_�IA���7��:�7�v-ѡ��g�#��H��9`gi%Rf"7���B3*��DW��Ż�O�;	��s�:y�`y�lTVB�P��$�y֝W�Tvc'�Ù\*!r�_G׳X�kGm�s���o5�$�K D�;_��J+_�U����eo(�b6��VcC��x#�VW��H�ex�𑠱E����E��@U���8��A��f/���]�k�;��b�e��JY�t��f�i��v�t�����i��ɾ!?�zjZ
Q�q������P?�)\�&I8�wv���-���nX���֨F	�5smA8O��W�5�{�2n8���r$�^)w^�ЋR��uș>|��E�A� *�>mX��ĘSůDq"��q� ��8|��Y��^���ԤGnT��.,o�CxÓ{��"�#~쯋��"qȦ%�%��;\�BT�G�L�ݭw�4@2My'�R46�7\a��8VRL=q�f�e�.bp��#�X�=��ը<�}h���A�������k���Ł2�@˩��%��=��^ �d9kL!����9��x�v�İ��[�!�}����,��U%�ޣ���l����߳�&�����*�V�$�Þl��7�H����7��ڭ ���Zi�ovpKc���G ��������N�#��ԩ�?h�� ������ �0�D����j�>�H�aA��1<DX�)(0'Q����i=��:f]T�(=���/F[����KbD.��]��\�O�7M�s�NJ.k���`�����ŮN����:R�q����G���T���k�C�ڵFHR-�����|"��7=ڡ!�D:'�c��r��z��΃;FF�3iu�N
�D=n3`��2Ү$���3�=�H�m��`O��������x��%BY�䏨�����͉��ݳ��:7��}q�����:��z�)��u�>O��#�m��T�Qr���Ԓ��GQ�*��-��rt3{�eY�o{6'H�s��{�dڔ������;���9f�1��uԞ�t$t�k����5,�4��'b�J�oF��U��>��	��"zڟ�@�}J9l�	�|�,�Z�A���X�AX�6�[�-x^�Z�d���;��[�4v����t�u\�D뇽��ԃ��82�y�IuH.��y칯�ϖ*ܨ����6�9��n�X���V3y�?Ek����hl�t��rx���4���2���Ƈm�_eH0ʺyZ���<k6iR��t���(x�Qd-7�
 ��@U,p`e�����YS"�cD#q�F�*�<��R�紵�*-h�mb�[@!}[��чZ��w���ut�2p,�+d�aKL���w��!]���T`I��3�,��� L���}�l�]d�6/m��22~�����NMxiV�^��K(�V�Y!��Vڑ����ښ"���Y��b9���ܮ�����-H��3��s��bk���_��Q�����h@�����	��x.�͈nk���Z��ڥ��AD&!���+n"�g:���mr��,A.��d��������6ǶW��@>Z�2������*6��r�8tg�SR�ؙj�x�ee�@�
�W�_�Cc�n3�\^��
�{V* j��4��.�aiB�J����6.�ڥ����p�	�r���>�3�,��g��,8�U�)oY� �5��zĝ7�)��T�w���N�Q�o�S��{�yoH���p2ͭ���(X�U�!��r���;s7�l�w��l`qI\O�*��GZ�'�x�5��쮏�����:uc��x��.�dt-dr����z����z겾��]��e{F�S!�`5�	�*A��\lm�ue,���=b�9�6�E3��Ɛ	DkFt�������K�\�sCn�&��HM��rs�� &��_�q�)ޑ��]k�x����Ho�z��c
��q]����@�WEU��k���jF�.�q4~�,G�č��.X�r������PV���ۯ��M��F� ��|�MB=\'�x��8����wXV���yY�GΧC�ۙ�
��$m��S����w`��
=��4�W˳���3�rL����5|����7�4�`��(8�
wg�o_��%d4��T���.���&�������{�R�������ZR��m���a��}�qW��#B�残q�~�{����
��/�9;�o�+�$V4>����í�r2H,�u�x�qeH��N�x@���0H-�I�F���+/\֨1����7��:�����D�(��>�X +��#v��x� �1Q�Y�[ ��QU5�#�b�SY�@�?~E�%`8�[Ɉo�|H��E�΀'�U�"v3;�qA�!�To>S=�I�% ����L�9��UL^�n���Ăl�2�L����pgiI��`��H?��[Y�I@I�i/�q�Kz�ʝ�H�9@��r+�-�d�9�d���H�z��~�?�5�W�ҋ�%�[�ճm���kK�`�a4�j�NL�5���t��镕αz���������C*ܨ��0A�-�o�'�˩�}L�1FoYӀHho+�z�pR�M�g;]A��FfP�&��Z-�Nu�9l�kP�$rceI1�/7ڳ�5�2���ǩ:[��kܟ�sYs\Y8n<�����\y����P⎭H"��Z0c���e�&�;�l�z��P�GB2�ĵ�_skGzi�i���BZ%�lE���֩
��
�X'�ˆA5���:�i~$5�
oXy�`I8F?�E��I~�{*�q�626;2\_�X+��<�ι�$���Փ�M�+�X:�X���vF�����`���A:�}�5��a�F���̦���ů�5�1�
I�RR��6�'	W�w����cz�ݹ���F�穉����7c�G����O�ϗ{n����kܲA5��q�T-�'�R� ������%t��*��$���>�5�v)��a�����>���5c��l�ⱘV�]�/�|Ti�I��ށ6�ߍ]�M�<��� �F���V�e�%RĚ�3M��U�r�OL�*Q��<l��j7�0��=��_�y����m ��Q}cHLTPp9�Ľ��i���
)��������0E����"S*Rr�
2}�i��YL�q�*�oNS���b7�0�L�V,��N��2I�X�L�h����G�4����V�pH�ң��d� �y�߇���{�$�h�=L8�5ȎaOp�~��;��X� =!u��&�8���2C��Y@|r�ր���C�.���>z�9�˫�aDH���釾)K����q2,��|l���Q�ĝwd5���Ari�+�yh�IvHl�ȓ?3[�4��EíU��E����[�!*�#��TO�i�.A2���7�ӭ�9��2�H�O��J��V�@���)��uw13pr��L-l9�/g�������Y����΋��M
��I��K�����HÍ�	�_�w~X��G�hm�����u`Lgn��	I��l�>'B����GR|�1s���K�	�y�#n���|$�,��C�RK�I)��i��S��!ӫ�@�v�І��5ӿ֋�Y0*ٌ��^t��Uxi���N�x���v"���_PN�*�o<�s�M5k8B���a|/XVn�߻��YKdk����<��ۿ�3�[�roi�[��&�r�r��]+5�t����7_�ћą6���{9-�K�X�����A�����i�6\FXX�	��ig.Q�����3��M��ce����F����W��
���XgUz��n��O��>3|���0�Y����C�ݮ2Q�"I��	�q����!,L��_��D#<U�}��� ��^i�!nS�C���_E3����?����"@h<�6��C�J�e�h��k�a���e��o�<�*ƫ�z�;w��� "�ܻ�?�Tq ����~:�>4��d�k頒�5"��}�b0����q����©�꓏m�K�k�ML�C�Oe�}���������k����O�^�_ ��ʫ��i�ꖤ�����@����1���fk���,�t��$.����I�1)*��YP^܎Z)��'�,��q�V��Gk��R���ۃ-,�O#5��ڭys�dîn��: cO�%��1�8v�x���YG��cX�W*���* EY(��>�8P{�~F��TAӺ��\�}�)�����"���\� �	���O0�G�?�d�#��$�ϚG��F�q����PRK"T�]6n h"�'a�����a��| �puحSIu�A]b�� ����j�K�[.�4��X���?���#�/ 8y���+�_����I�R���cv
W�w���7w;Ƥ��A��ӑ�fǄY�=�Z�*���!�f�t7�nb[��m�N:n�ꦏ�F#sW���̞$ddYסI�˘D?ۈ2�2��!un��Y
&=Ʌ���O�n����
&�T��h�(��TF!��T�6��6x���Q&��y�g�U2���27/�i�_����q%��&�[�4�c�&�Ew�\�h(���U����o������3
�� D����q)-����w�tuuΡ��cͲ<�-�f�Dw��x��	G̭B:^���1=�s�H��7��PV�`�b��\[Q�+S��G �PzGSo�F}R�+:Y�.ؤ�E��!�W� B�	�RT@��{�Eq�"��)�!�h�a�`
�ٍ��AM$�׳��B�ꇲjG
=���G�R?�1}|YYb������X�!�"�:�0+L?��Ք����C�����q�w�C�r�iF�Xo�N[5F�D�$?b��oD���@d���JZ5hS�ڵQ��r��H��(6,M����򨖯�[���w�Bj�8�7ћ`Ke�@��S�3}{�6��O���x�HO09�,��ۻ���$�X�������EyH̻k��v�W�����v�h��.�q�6��y���/�Ra�������i~�t�نC]����$,���@�=z�ݢ�ߙ�nB��K���⯯�e{��	ײ́��)�_�N����h�Bi�6�۰2�=h]�fQC�iSu.���L�v_�`�(Sl�40Ura�Rٕz������:ޝ	��4���A��}fZ��)B�NϨ�'�[)��T�e�/��o���*��~ʗi0wh��?�?1��~���N s����l�q�W8cNj�Q� �iP4&�h�9{��L�6(e���<��#��qv�2��^��N"-Z鷫M@���P�:�8�nm�*t�*D(��aa�]'�ql^r��փ��ґ.Ro8��a\�@�U�K�����{Ð�Ey �"�F��W3q�Ud:RT��v-��N�^�I��-=�m��f�N��U{{K�����Z� XT���ma_�g{��B���_�\� Wo'�~���'7�R}���d���b�����O\��K�SPw�qqܞ�)]�F��y��6AF�C�2Vmφl�-+W��1a�z�%W(�~dn��۫Ur�{�2�8U��w�����`_�Z;k��;�-��z@��o��a+x!x7XǙF��ԐN�����^w���N�	��D�:���DWzL�Ҽv �b�	�~�1��T���-��0Z�`��(��J2N� RF^A�$B����'�e�Iw�=2�k bPM�T!�څɲ�����`��^�����1�uq�������Uo���6l'F�Ů�e�f&�..EIư�Sc�Q߃-c�(���4i�d\�P[/�U.�u�{����ndE��o�`�¥k���j@����g^�:���A%���\�#�e�t�����_�bPn-�D	�=�CAnr��
k1�W��k� ���P�9����#N��?El �p{�{}������/Py�7��0�쬖�ٔJ�P����H�e��V{J����RJ�=R��y^d&���e��}�6;�+f�O�4W.EŹ0G�s���j�����_������@!�����ff��z3{x�)��?Z��]cVE}ˈ��]��b~cP�L��#�u���6�;�W�{��>d��ȫ�����Í��=��8�gb�����i�A[NI�E�Xa@�%���0.��f�ucaN����ٻ����U�4'C��ž+���o�T��z�1f'�ӆ�[Q
���+~�c�VQ֝��?��U��K�!�b�$�&Cr�͓u�&��ޟ(�J�cI^V���ښ��'_+�P34촥�zfR~�1�om��0�+Xz��ѥ����xl(P4��~��NtL�>61����$��)׮q*z(�$5$�5��V��I�Xz� D��Y:�U�G$֩X��ysV��&�xi3�v��6;��r3ຎ�Z.���	�_O��GY���������S�$ v�H'��zU�$���bc��nnϸ+ui'#�+�Gu�PI�[��L�(e�ʞ΍�Y�s��Z���6���C	Шesr#�Tl��^��4��]�u:����!?���+��_ͣ��ˀ��V_q�\�H1��฀�`�Xt�\��M,��L�X�}ڡ���Y\h�%}��-B8pd��[����9B�~���5���G��OѤ>*�:�
��4�w�%^�g��`Y�], ʙ������k���I����,�k��[� A.��o��뻧OmD�[�W�Oy���Ì���O��= �:�~����'�W��ok%i��>�N/^����Y���w�f����L��0�����k����5�W�8��G��6��M�B�c���!���بv��0�ੜ��ٜ8�q�6�l0�JD7�Y��B����`1�o[����R�_Ab������3j�X���2�ÿ��ޭ��V�Caʵ����n�oL��~���/��&�~"�{��E;Z0~C��]݅��r�Sbw�����F��Z15�E"?�.$bwt�1f���&q��u��Ƙ��}�䑀c��<��BL>yˡ?4�nI����ibH�y�uVt��E,mr\1��2��������O�Yא��٬
[��ݺ])R j_�!���I��{�2��H�ן�A�ԛ�}���4E(�T�n6H���(�G���eȑ�&n,n\B\d�R�.d�H�qf���2dH��:~;x���-�wCIAV�=
M�?^��.P4WO�JLX%ږJ�m?T� ç~�G��,w�W�0a���Z���/�e\H���v�~6� �`6VKSA������.hh���Y*L���<%�Z�����`��v�Q�v�
�EZEx�%�slxbX%.f>�״^Vg�h���uCtW���Lh*�C��!�e�0يx3��u ����<��f�HF���ү����b.ܡwX���4���̰������0|!g�P�5%$�\�PMY��񭾦	<�b��5�G}��L<:�u�t�\���� }f��V���>�f]cT�|E�T�>Q��4N)R��;V���o�	'辋�a˾�3�Y�P�$�v`���7Y���P��3�0�59��&N��ji7����T����)Nf\[��[k���a�� j�	XF�J�g��	S�K"�m��6inH ��'�8�v=+D�ub;��s�C�����ˁ���	r_YW�Ҧ���տ�޻�M3����s]�w��;WΒs���u�Pk1^�m-��5@ހ�K%A[�w_>�~Nh'.�n�IP�0���ӂ\��r��S_6�3�Лa��'�
��oͼ�-�g�W�}��~�{l3�DP*@0�
"����?�y$l�O����Ap~t�'��$�_�ŋ2H�,[˯Q&F�Bs���Փ���Ӗ��4s�,I�H�#�0��z����Hn/��=�]\up":�[�y���{R�y
ƫ;��?�zg��4 �����y>]s�p�n과�ST��l%������cT͝Ii�<
���g�\��\�
���}65��0)%�l˯�F�w½w�)J��x���-T��]nJ`�o�p\��ڢm���[�kz� *�~F�Fc��z!1�/y,`ԯa.- x���μ�	� �_��w����?(�yՉS��gF�m\7[���\�u�4^b�b)3eDZn0�I�!x��]�)A�`�uΨ��,'ym���^B�&.��!�@H�4�/;/����U�ՙi���ſ7��1JSE%U�Ha��hy�z��;��:�Atp�4�?��h���$���,bYq��俋`� �uϭ��=^a	8�N~�tIX"xx}^z����Ԥ�xh3��ܠ�zK�]E�:�ћkU!�������X7!1�LԶ++�a�s-��� �G_J���.s={���F�eF*h�^�߹Y�b�V�6�P���)��)CKS��^�����*�RoX�i���KpfϏ7^���p�^�4�&p�����P�:˳����z�D�ޓjV�\2=j�򎔆v����b7!���	}�Q4�"Nߑ"��G��{������Y-q�U2t�W&q4��Z�hz3=�\�e��E�[�Z�����ϓ���fRS^��DA�������3��h�#eFPLs���w�q8�'�tin�ce'���?)9��+s���\~~�4!�ztТd&-T���+���t���F��+��|��Unc��/�M��Cv��6T	i�[�n=��w)q%"u�K쿝ГA��[T�9�UV��������+y����m��d����;�D��>�?&�sR�V�>����ﰇ��Q����\<Q�����x�6��m�uD8��v�Ąw^)C!
�$_P�o���Pl���uƽ�3��X�d��< ����X��=�@����dnR�}�d��r$[==�cY�XS͟���a1��q���S�s$p��������(�>к�����&o�/
e�)�Z��cڹ��NĨ��!�ݛ"h\�1.c�����+�aAD.���6����3Y�B�_(����!bx��y0+�h��W7ks�2X���"
dA�+e�4�2G��B69e�"�{R.<z2�>��#\I�A,�h=!\h�۴_#�b�z(PBڏ'�_�M1tU���lm�I#�K]b��q�W�X)��EɒWS�U�DҬ�μ��`������U�d���U�!4ҷ�1*�o��?��;�4��t=�� �H��q>Yӄۃt�07�y.`3��pt,����Q
���	��ʚ���̮%�ޤ��}5d��%C������Ӓ5G͇>�"~b7�[l�J�����$���$o���?�Q:b/���Y�.~HB]��2a�4��Z��0�p������ZA��!OJ�:u�ȃi�}�顢�pɺrS���r�&B2�`��mtx�0>�Ð2o�xmt�f���ɮ�����g���5�]C
'�\J/B���K[�GV�){)�&:
"<������n��F�����*��f��|����CL�q❮c&��iF���Ӟ&���Ώ��*F���8��3�: -���&��D_Q��t9\3�B"��yb(c�:%�h���q��.
NS���w�C��ӎ�l�����O)[���#�]���x��4�GB"#9ѝr�='����>����EK�:5��[�n
��9�rc��2ݔ,��޷�e��8�U���C$u-�O���X�TN��G���XS�uPn���5��:GZ�p��+�Y=�@=e=��	���Nw("H����`b���q>�|�/�!1�σ�_ �b�a&��~��d�w���i3�#�ߘ8��^1�2�E�*E�]�!kQx�^��|��v���1��K�Z�X&,E����K+Kx:v�K_�a�1K#ZG��}�j0C	�HfDъ�Ч�֨)>zp�1�g}+�?�x��'[�PԫPfY���R!�0矰e<O8�G�AuETzu��U���K�Yق4�h ^��h( x�j%�3G���&R��}N��� ��,^e����N�`�jӛ)E�2�0"L�a�s��{ug���$�#R`7�G]/�uy��P!�o�S�b��j��$����J�G_��d��º��Ď2<#��'v��U$ou3볐C��Yt<f�:��U��<y���o�Y�t�՗��VT1�_�m!��>�'�x^��V9"o���5��Ҽ�&�߁�%�"ph�ET��g�����&PYc.��M����NP�3�xeA� S�'�%�s7؈�ф���rx� K�ɱ�����`���il���mH
a��>���S�fа��Z�ޱAc˵�N�ah|���Ɋo8�$1��|���V�I��[�������8E��Ӽ��ic">~�`�}�U] �&N��r�9��-j2������7�ۻQ�[*ﾜi=,��b�С5Y�b%����[7a.��AH� �ڢ�H<+�X�j���ft/��ɮ�*�ʓ0���~�L���`��l��`G��}�1�^W��+�2��E��$���)w�§�gI6��ZS��@�p��\�dS���3�����,�E�E��g磇�F��3��V�z{/'�Nh���X����r�a�bg{`0���b1�G��D��Tݶ9ђ�~�PX�h���yF���(Wa6M��M���^�
H�2�W��#���[����(�ЛH����!��<	��1���N�P(�����Kf*�%D���� �E��#�BC&���7�Kf�n[q�M���)B������0:��h4�ܵPZw���FHX�oc#�2��GV2�ӟ���ϸ¥sn%��i��tsH�3l���P��AųE6�J��m��6�8%���(��^�X}Pp�) ��oy�.<��uz�c쪷C_i�5�kB>/�3�dW�Y�`?.��Q�(&�{���3q�į�3BY��Ͳi�?pTb�"�k�� ���Ra��T�T#$��]��p4�;ɘ�*�N�L_�^�����-V�2�]�t۬��t�I��g���t4�$:fǋnݙ7��8K~}���R/��N������Ϋ�����s��v�O)%&�0��\�uAŀj��N��7���#�^K�׏�� �5���Ͱ���%��$ؗQnH=ȑ�3U���ԧ	؄.#nqvhM������rmt�,�g��ݿ�"Z$�/4�7-�5$Z�Fπ����"���!�����̯g5���1�5Ѫu��X���:Y^���?o��ǳ_X�C�}����fuӋG�i��:k��v�|��t��g4q�J��a(�=G�1�Ě���1�;AH5����3�[��Q'~ �ל�������y�q�d*Ʌ*�/�����]E��Z� Vg�������SQ6C}�m����s+��"m�䘛��l:���Lq���j��"���" �9Ɗ8@g�-�u��Փ�g�V�"�}1�ku��[� ��izv.��bC�D�_\b5l̜X��&&oq]P6��4�{!p�y����~$ (�����M�<hT4�r(�9qe�';���A�ZP|�yJ.P��Ũ�*�������#�1���]dRk
/\,�b9ƭ��&Q���R��-k�\����?s&T,E�S&�0�C\�Bt��S��Ш�S,Sx���ol�JO�H��4g<@�Zv�anT֓�<����l�e�U��U^1h���[t���f�;b��|���|D���FC��vq��_r@�8�O7}	�I�j��&��x��.R[��N.+O�6�q��E:N@o+�ܛBĄ?�֯�s^��q������4L��,�_؏_��3��.�C3�����2���z�ҕj��ڬ�C���)�bs�u���j��f3e��8��#�H_�6���eϰw�}T�cAQe+��i�16����~�W���Vv���J���J��Ė��y��*��ԃ7#v�R���(�a�H�5�wY#��@1��Z¸n�7�`�$;{�^�S-���ga۝�=�0��(Đ+D�:�i���&.K�U��;ֻc�8*�8�o�X�X�^ʖhY��ݣ�A���ia�مwʖ�{���ݿ��jX��*�
�HJ]� S����րD��
����A���{�%�Sl�X�˖'�S��t�n�b�ͱ��߄��^�JDH7R.��~
U�cg�q�c7>N������Ìw%�I����O�$n��_𥳐�2"�$�-���̻���ݥHc�dџ���j�:7p�+6AM[;�I���X�xV&��`mϚ89����i ���R��NO[y�U>����J�XҤ��@������e�~!�wWRc%�����$�6���ݓ���ܩ�)�u���+w����|_�K�$	v�A�K�,���&�Z�$�a)� a`e8`~�۵藚X	�������{h��jm!Ӛ%=�E��ֺ�%s����`��Q�:�����h#��)[g���� ��"�n$wr��|Tby�����(���Ve|5����Ǧ<�Q�5(&�>�1&��
�M[�'��!�H����m�B?�:U!��(����ŊȔB���Ґt;�#	�4����$ǆ��O�?�I{b��ܟ��,u�ą���+f@��M^��7�?9�5�%S��ׇ�s���
�H���^�>���m��A	諺C��
�b�p���/�����)�7��E�e�$l�g���N�Wۚ�J�^�[�.���R^��e,@�[;1�=BӇ�eS�����4K���#����r�p}�_�+��S����Ðf{�D��x+����R&�d� ������|�4MW�WW�,��KM�j�����CZ؈�~��Cr�P��Һ��_�w�K�C���<�n�7�_iT���9�	����Y0�߿���`�^�������/�A�w@3F4��+�*�c_�u�w/� ��S	b��l? F�;L��Y�).{x?(�v�o��I�PU�d�Q ���f����F ����Y�E�n�n)b�2�����	wG\zrf�Z43�ם ��1͒��t��� `��\ �[�o��lu�
 �fv�%���C#��:u)"��+��8��9�ဨ㼵VG��g�~�mX+Mssb�1����`���r(��x�᪣)Y)}���qC$�U�O�d1!+B ��B�c��l��e��;o���;�O)�)���v�\V��Y"gF,+P�x;9Rq� ~��l���3��Mն����@��W3����Z��w�fpU:��'c�l�\�v�D��Ț}�y�s�/�t��o�E59�&-��7S�4�Z�o��e�aF������B��"\	+aF�����Na��+�BOq��N$T��S����CE#�a|A����t��l�M��]�L���D�0W6��Z�����2����goϪH�F�~�n�L� p����F_����3i�QG��҈�ω��Vɞs�]7?����Y�\}��MЎ�<M���P��ʺI�*�ńr��Ջfԑ�����"�sˣդA x� u�U��&T��@(p�V��	fhk����e��U����rFe��NK�8/�\�-0<N��+�n�96O��hU��w�@f�ǣ�