��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<JÕ���<g7( �^P�}<r&��+�����9�n�c�0����a����!�6\���c\�������cn�m>6ۂ���|�u��lWk�t���(��'*w�"�2n�E]�K��^�h���F���\-I�u*UW4�w:q�m�.����U*2�p�Q�^`���$��'��4i$�0�"��S�D�h&˲�m,�IPy�ј��4�����ڻ����Mfj��Jro6��Tq��es1���z����t������ȺR��4���Z�*z�H���Q��j�P	+z�����K�X �d�؜_ݹD��f�.`p�>ڕQ)�fT����^Z�WqG?��V�.^���ؾ~��<aK�
�T6���"�P�6�ߵ���ټ��Z�=Q�rT}A���>�e0C�������#�/�ܿ��O1��$�� +-D�~��>3?M]~�,�⨋��4�\��Y�2�`H�u}���w{P�)g��&e�����7�P�%m#F뮉�FV�~��uy��r?1�}�FO�c*��J�Z=/$ls�įB\b��r~�
�k�?ۃr��&��=ͮ�e���y���D�S�Y��?$���wR�z��m�wG��
bi����{��ͺ(e�~����s�q{@W������7��&�|�~!���-��^l �5�:����KXL�HO�J%X�r��R�N0#��������WLP��>F;���ʋR�M��ڟ�7ǅ�9���u[��=$�fA�P
u;����=-�����|~�I�x��I:��|�sEK�
ke�Κ6s���Cm�����y�s#ve.�w��?�c�"�(!������k����Hp�&�<U��(I�6X���h}T(�����/ޫr� �cO)��dh��P ��#w���$���Ǩ��@��J���'b���Н"[6�_z2�,�T�Ȉ)Z��1UE(��z���0�Z���w���U��,x�	�v��$��~��r����ڋ���M�:���ۓDK6r�C̣���c�N+\`|[�7=_��A��/CA��x�<�$z�����~��VBkc��k˘���w�%?&�7��y����j�~��7P��B���0O��H�n�"K�/g���ٙ�Wԍc��ة�-��hN���)�j��>sZ��T���9"�nv-J�<@�:�I-�޵;#Ӹ�L�]���ݾF��p����dqJ'r L����<�}�x .d)�t��V�~��:bE�� ��&۴����0L`�c�_�%协_|E�G �g�6�W�Z��zM��NaJo*\z�rۖM	)8F�8�_$�d�X��M�ƀ�ͱ�i�@C�-�~QȈ��̵??Vfʓm��~�T�Q�qrw�����ap,��\����;;�K2��Ֆ�sF�
��akG�J	�=yt&Q���8L9��5�s�Es�PO��u$[N
���K�K��L�T\����k��7���I����������!�UG�f��� �ſ���7��@0,���$�CQͼn>�A"F�m��ׯ+���<:{� ���N,����A>����XF�=�΁,�n���cq�w}b���h��[>m������g�*���P8�1�$���=v.�_�Uآ�ӭ0]3p�!���
^,�Fj2?jqo�J�Hej%\�k6
�J��d�15��ʹ�6�7�\��b0��üT*�(�hj� ��6Ⱥ�O���<��H���y��g;���p�.%�Y���?HT_Ѯ#�;��ؚ�.b�=��yd��������,����M+����I;G��{���(F�u@�'�D�HZ2.r�I�N�9\��DJ������)m��4��ķ#<��� �	W�)8Ų���-��/Y�T*@y�|�$=E0ٱ��<n�pXJ�Qb�|�{��>M�XU��g�څ8|Ge�>�ڱ%==�Zx�u�q����/~]R<�7fYg������AgO��u�|��|hc��1���e��q������F���h*�y��bRd�s.�7�wAw��8�[�������i�d˫B���c��%Խ$:�� W�C~�Zo�x;����b�&��{�-h�
:F����f�������:�m�1xXʮ��<�b<5��;iO�m�&1�����HQ_�� ��EQT�ΎdK��fTk���e[Ƭ�C9�cM�K��5���) ��T���qj%��-S�?�P�/��U�8���úP[WB#3��~��7�~���mM���lq�kj�c|��[&�{�G[]�~l��sD+�W�~RL�l�T�����k�(񟃬K^ڪ]��\���{�DRB'<aXq�8��)��1������E�)b1��)�%=��q�������f8��bŶl�? i��!������7A���O�ݗ��m�@FY����2�����l�n�xjGt�`&�0��~ż�[r� QT���ej찲�SP�>�=l�Xg�b�:�����a��eҟ�Qd$��P�T�W����(�BZ���͛t��8�o�Ƭ:�(�]�^���Ĵ��,a�X�(,)�7�`���q�$��Im�]�VP�e�yY�/z�L��	��FJX�A��Rg�/\0B��)�(��!����F֏��_9|�=��@$K��`���G屇���ȳ�yM�>��m�)c�Hc&>��R6�(B���U#����{]�����U]���t�yGx|M5�S�<a��ߜ)	\�G�>5S$j�Q��8�2P�c"���W��c�r-�u ̝����;C�+Mʞ GDԧbiSsR0����<i�\��vO�K��I��Cܼ����d�j��޹�ԋ���H0�-�Js�9�8�g�d&���Ŷ�����G�\���md&�������i"�쳑�k-�E��r�.u�i
y~Ť�����_��C�-�E1�(h�kƍe��C4�v�|?>D�q͢};�3�����
��c}�R����D4�׻�u�sŇ_8�$�FMcDt��L�}_:�D�.b�|�2um�ۯ����������tU��
.?1�"�Q����L�H-�3z7�ouP�ޖ���z�����qqv�!�=։�|�x��L��msH�6��:�CE۲�m�Z*����!aXe��v:��Y�<������)6���Q��H�Cř;X����A�Ǉ@[>+�`U�����ͬN@F9�$d���a�ݱ�W� z������������i�%-]{�i�?�+�v]����5{z�s:M���;	탦�QTl)l�X��Fh��</���q(칙������Q��	����-�}��,�>� ƅ��EU+�ߔ�j��`ʟ_�-1uv������}<X{m2;�1B/�q��ZG��z���:�oY,*�te����M��U����a5wOw*:�0ͱ�ި� ���Y��9��g�Vč<�$�lmq�Oi
|)6��Gm�'![4�6�}U��v�1���IuiF�
��iGc����>.�P�=�2�r��*� ��.��n�n�`_�k����(?�>�eqoYxx�4�����WQ���zD����˦O˛i����$�
�i.pD�C��Oh4���y��M�������� �5�n�F@%�fv�\F.I�d%Eۄ�*��pyh�Z�"}�cV� P7H��gd�~{g}�drq��Y"��0�3T��M��p]�$V�^���yM~Λ1ep��\c.j�@� ,\�a����;�m1m6G�؞P=��U��,[�6���j�1�DE�P���To��i3�.v&��3�WTI�I�br��j�'T���A�TNR�C�v�^}؁���U繝��hQ�r�w0?��SK�!R�ڭ�)�+jL �X��;&��A;��}ܛ��)8����
����(v���>r���;|�g,A0:#�v�B^�䮨6N�yz��T~���A�V^�jʚ��k]z5~L�������#.!|��o��ͻxM2٣%�Mt%'p:�s�@>����x�X��U�<�Ƙ���(�s��+�Q�rDв�W��q�G�b3u��YJ�yn�	Hf"��ۆ*�{bnb	CQ_��P����<��l�tJB���A�`i�
oG�]��.�6��S����4��x	����V�B�UL'��~��R��{6b8x�RbU�0�/rQC��#�[ 2���<�^��f�۪ۀ6
���n��am~��!�ZH����0�^������b�.�w_e�~*��O�õI�VL��A�Z���O��K?�t�e�l~[
��;��܍ ��ZXo�ӦCXg� Z)~=�W`v�b�����C�*�Ī]��wud�N
ŠeV�mv�¨�#�0�F���p�OtO�:S�*���g���8A��bP��a�(i-0��0���' �=z�kge��-r����?%^i���v]��6��y�HI�kb/��(>�=����G¦��ˇ0�2y�n�|L��?�}g!�N��)/8@צ��㷆���^�����yz��.˟�@�\W.�2x#3%&�PYz����ƥb�+����c��*c&�����;�HP�^�J�I���wSbM)>x���� �1:�)��'L�U�EC��/�Gp.1����� N�����3�W�{�R��=�6i3�B>8 D�R�gG4YR��h�=�[)s�0�@|�沝��7$1��bpc0Y_���aU�|��!��gr�<Bw�a��z��c���&j����qd`v�����VeA_��r�r�D���$�Rn��5Vs|�m�a�yHl��/^[�6���nh�ٳ��O�ͻ���7�92oI�y���ԟlyt0�����ͩ����3;��mT�q� g��b������lI?g N�?�9���$���t��OP�V*ʥxtNE���go<"v��|W�R�v�U�4���*�և��-���W��9hhv�]�~/`"<ĕ2�\��ڭ�kz7;�W$�Ծm�:!�@GxW�P�I��}����~>#��>{�H��6�}��u����Q`�[���(�-�e�UYJ��/r�#Vs�>k�
�mO'B�V��xu�V�^�U})�^J��X��u���g�q��������[Z�r�Q`B��^�z#�X�nF������t�
Z���H�c��z��ǖ��XaMgJ�`EE�mX��h5K���E�u�ڪ3�a����=߭�rC>��"5|i�I��*�ր�=q�Һī�"�4�x.�8nC� �{��zq�ً��*#��9����M�v>ƟN_�8p��W�u�)fc�̠ �lֽ5S�;&��W7Eǖ�ۆ�5�*�\Ye&�ZH��F��Iv3���� ��g��/�z[��WN_̀T�u�rB.���N��d|c�@��wgJ$O?�>53�%�9R�},JX�	)cJ��8��{���sAn��O
����ós#�e8����VQ�@�}O���9:��jI��ˋ��������
,P y5__X��[��T�s����
��9�I�,��D�i����1g��C ��f�4���x<�{d���=�o���,~�ȾB�E�K|S@���,�MB��奵c|���y��X�U�
t���#�US��I���PQ�b���=����`���@�^6\o�r4X�X���_��ޕP�gs�v�#��T;P/>�X]�1h��'?(R�'�����"���Hdz6f1n&��U&b�3�S�J=𶜏py`���<7�mL��C�Fh���d���>��֊���M�oH0�C$�P�>�_��=?)��Z���m�߆��O��B�>��<��v9�K��L��;u��9�%Xx|����2CԼ���'J�뿅�^ukᔢĈ���VD�����ZW���-_���>���qWuۙ�H���Q)}��G;c�`�����ڴ�#JZ�Pzwc �R�;�:� ~MUP�	�-S��+"�	�e�����|2=���˘������a�	�ޭ�ØkaY�e��
.Q�!�1�Z��g�����;	6��y!��{ U�y]'.5�(�պ�g:�t��l�4u"�K����RI����5s���{�YPca�|렭��I
�������qDhɄvw�_n �����P�zi�h;���'2�K�{	(�v�G�����+M@�NK���𔋺[�{%�n$V]=��U&9֐���+W�&�pP��D>JӜ�'r��' �.l.��~Z5���� j��;���R�G�%M]��
Trf4<�A8:���_���BY��]�F�ƪ�on�)�
�d̀�	�aB�Ц��v��w�^�'������Z�l���$��I@r�E�$�>������Af�
ԗ,���;j� ��?�vP����7�7:B�PLJ�{�@d�-)�џW���T]�Y����~�����:������������<
����6��0�xv��Wc�\ȷ����k���i��>UΪVL���������IQz�K|��$P?-����	�\I��:�&^��U(����C.�\�50`���]⺄YS!�;"[��������N���Mq�j�*�|��慍�D��>�g�	���7�m2A�~\�d�ڙ������Ȋ�FcL:IG��/���~vz5&�K?�4����`�9�j`x��T�
č�'����"86��c~5/4����� �{c$P �TJM���i{�d��$�6Τ��q3����:V>���0��u��RX���:����h5�f��f=�����i�d�-�z��~6�ݒ�Jv̂r$?g�&Q��%����s� ���˹ȕ�
տ[�A�е0}�C�W�RnЀP|��_��H.�;MX��0�'C�v'1�^l��T�j>5h6��7o���!@Y'}�����nyG��$ʴ�PA�%�.��B��c��tN�H�{_�R*��)~�?�q��mƟ�����H���y�XF��Fzz����,���P�N���Q�{��������5<p���Yf�ar]����Ƒ�s61'׷�gVA��~�Y�8A����Eu>��Ã?�q 7L����O,�_��wr��� �{	|:��W��%�#��e�kd��v�N���]��0���|ј��)LnN�����_�ܭv�'ć{���?����@�N���� ��Rf��!�eXva��j�����+�pM��[;DO�|�c�ҕF���t�������)?�`<ʙm*��������2���S�Y<,�A>VӍL�)4-��qɥ�t��mm��1:aF��+�u5\'�8e�9�jً/CUl�X$�5�w)��m�7ZL?�H2����=WEx�:�������M��9 ��y��uy��Λ�G�#�G�a�̇GA|S<֔�8Ѻ��y��4��ġϓ���I颒���J��Y�65�T�@�Vġ�@��5�:��-�w#���+�=Y�5$(��ZP�p�=8�e��y՞��h�S�^�w2��|!�47)���Qh��X#Z�}�n�O��fx�,1\��&�@���MV�Ɇ?��l�pӍ9�%(�+3Q3NTu��+�a��l��F!�<U�F9(ܥabܜ�=ڸ��������.��*u�\�����~�cm73�)x�.���*��dzs{����@�� Wфuz�/7�"1�(LN)�\�$�X�'RrJ�fJ�c�z�������R��Ik����ڒv?�*|�-�p��>P�5�����x> C���NA�-�V�ڤ�����{�?�j*�KJ)�o�dY�C+��rM���}�L�����v1h����!�5#v�����ێ�H��xu�D,8w )&�~P9Z���N~o�Nl��:q�&��%��&<����备}qf��g# Wl���M摮��Ž���M�կd��D�!�´�/-�[=�"����Kv�=��Ы.�/�˰�n�@*@8B<���S�d�z%R$����/�B ��޹=?3�gQ��t�%��H��327�b������g����Os�Ю ����4���4����6�YWTN��q��-\Y�ԏ��W��ӗ�^G���^c� l��ET}�s����֪l��	#����
M�!`l��s�u���;��M$ׂ�m5���t���f	
fmq��-}3��r6�Z�M�*D?تJH����'��5�B��A�p!|�������Yn|��Lt��aF3��p���*��3E�E��!VQm-�����g׾�m
.�F:������BiD�2�FC����8]h�H��Sc���O�l���
��3��NpVeGG����N#ǳ�\u���m��%���(}�h|���Zb��A��S�E��,�2��Sr�c>`̚QW�7j|!<R�DЀ���'Bt�&5�B�\�
���~nؓ�Q�,s{�Z��䦏BH_phFy.a6��M���D��~w\�7S�)��q�6�z�˓#
!-���Hd[R;�@&WQuI}����WO��F: