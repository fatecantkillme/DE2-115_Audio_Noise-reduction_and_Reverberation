��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<>X�8���#1���bO�'����F��dM�z6N��$$�A Ӭ��)�q��u��ZH�i�D&Y�YŒ���+��K=r1�������w�1=s��3Y6�*����Kto����5][�����هc̶8�N�RB����W���H�c#91;�HS��B����V��Ӯ襀~��"k��,��*�R�,}Lr��˒�O�������:��$��כ��A{7޶�Wg��䶝��#���>B���{Jt�o�ʦ(h*���7��x(cK![It%]���=ys̽ъ� ��f�ۙi�G�hT��4ݞ�X�������-i�i��t?�)c�#�	Iq��E��c#]�L7Z=�E6K��ELqZ�?��:�<j]����]=�D�O| ��y����y&z|H}\XTh�j`2=��ύ�������i�����:��7�ʾ;��Z����`7���'B'#��;��d)�Z��ݠ��$A���XJ+Ւ;��÷ @ڔ��=�\ �T�U\���@���ɅI!�
E�4�b�^��<f O���7��:��2d�H�����Մm���'#��+����D���?������8��� ��֚Q y�*(R����-E�H�&�iAn��%d�!眫�w��F�-v�������K�����->7��� 3�t��n�#��ȏ'����I$��x�����N4T�Sݡ��Da�O5Fޒ�w�#����,�H��NiV
��q�} rp�
XjD=��x%u�v��_U"�զ������[&��q}�<��@Ρ^���-*�x�f�lE<8����f���x���gE�O:a�f?ۇ>󯰗,͓�	��Id���_�<9`�eJ;Gc��{c+6���GrH�m��n��<�茅��Q�u2�d��q���F�Eh���x�����,ǰ1q8e��Z UTl^�/���H��؆�x0a�\ ��c
 *��y�H�i���j�G7��?�
R�ˊr��m8�Na���`،��e<����L�R_9
�C(�i�"��d�6D���x�*չ��^)�JP��Ck�wgr���[���nѱ����cٺ�4?�"��Ck��%M�f*]�yգ�nC5�\��s����?��udn��Mr�5�0/�.����`�tnm��O
rs�X��!Q����a�^.o�{�-��~V1~�5o�5y��9$^"�Ө%RQ`���:�R#їF����N�w�fK��";��������!�M�V��㎨�2:�N31�laB@��B�承� ��x�m@��x���[^����j��R�:��z7�>%�_Ļ�����d0�q��O*���'�l���0.x�J�W�>
p���[Qn$������܁Z��rTQ�(���?����>_��Ud�+-�fc�ׇ?C���:l���fY�h�t�0�V�*u�ʤ�(J�i��ͳz���M�Ne߶$ ƥ�屓�6��Bv��a�(�k��V'�̓����R�bY�9w�pξ�0�ūU8��t�Xt�p���
��Q����}�׊]�����@c}�=l�U-�{g9�29�KO���ڣK&���S���2�5��c��ڠ��I��3��R�����?!df�I��ź���ijI1����t2��frz`\�K�@��S0��XûiN��/@��-�Ϊ�%��8C��S(�4[A1l)\]�Ԝi�a��t�3������Cf�������̣��������v�k{�y��䛿���Y�MP��3I��9Ҧ����~���C�c���:���6��`aփ�Z9�SvA6"�̆�&� y{��͂+���A�Z,>�N��������C����f���Ev��$`��+9��� �v��hQ�Lȱ�t���9�Ӥ�+��1ʯ��.x�{��X������d����'�s�UwU�}���5�
�2B�q�L�Q�`5@�]��_��=���C��`r�u����ϷP��^�y�>�_�q��ó6 sCy�=�c��������W��6�п�	r��d�H��|o�0f�>�����3��� ��TylP�Μah��X����f�Gue�K��B㗢)P %E�������G/�r/ԩ�=�%&���UK�9�'�\��B�Ӷ�!��U��Qt��\2Ɲ�)񁂡N�����S��6'����9U�e�H^��Y��":�n�ߨ^��O�=�49�w�����$�p ��$X���Z~ ����+��V���?g�:�r�=�
Lz]NU�-W�jÄ��oO��\���`/�TU��Z�R>������B�S��o�
��u����5@�4Ԗ�֕��*�Ů6�.��Y�t$�R����aԶ8*��x���n-�x��H��G����AP�{�VI#�ɢ@< ��cSC:C��gT���ic�SЩZ��4�٤ҕ������d��B��B��T��4;�G�L��?�{��?{#�<C$w�T�H���ȯ���'͒��&~��&r�QF�PM��kt�$�^���3c�AS��W5��ޔa���×�y����������y�O��:u�i�A'�-��}����?
���x WL:������ɱ�u���������\�ӎ����Ll�I��d�|��fWC�q|q�H���B2�Y��!�9��2Čد�2P!�x=i�5�DJ�:J��.1S���g�Hݗ�W�Y��� ��i���3�{�\��^հ{��P����9��-�y�I³)�25*���*#U~0X�h�����V �Z��~�(��&Gd��f�ү�1��7��㔢/�6s��ܐ��:K ���������R�aW�q�a��6�d�-Hl����ą��!~<��$A8���WS�>i[��~�.8_�h2�}YLkB_8{,k���-����.��`E@���2o��G�2��`����a�Kh3���%�F�o����h�C�HD%�=�k����ƅ0�x��G���a%܄�Wy��c����Q�S�U��C���J�/S��k3O���{������)ɸ�$���/k�ٕ��Q��p�0���d���3� �'��wH���j�w�oN�ZkT#��	u�OH��D)��tSh�"šj�+��󟤝B�f�l#f%ɘ+��&e���j�V��@�ˮ��[�\)���If*�]6�!sXqɥ�FA:\6�na�'I5O<�H�ɫ���Q��J�����t�.���Y���^���8���X�έ_hȁ/a'��F������E��T�1+9q�r�	|��|Lx���g�	R�4�6�3��iƇ����,���G���ڹU���-�O���r��aC�nq�'3~�����W:��	���F.A$�R�͕:�{�J�(����!��H��j�.up�em�n��a��H#*���?}�G�I91e83>D0f�2��YLw��O-]M)�8�F���$�|�D�!_�Bko �q�KV*���}s�F{��΅7�c�{�������To:�!�2\���.�]�$gpYTOF�G�fC���֜hl*�W�sȐ�3��H0��FZW<�=&����y�Dw�	�X��2��I�cTy�^�I�MM0�2ź�=8���ܺ��s�Պv����*m��!�3+*l��!��N8s^zс��B�C߶�9G�����xV�F�џ����-�ßCD�;e���و�٠�}���b��=D�)���{zL�����99rQ��um����5�.�nO~�V8���_�6?1U ~EJ�`NuRCG}]����&�Z!�
W��{鼃�:�∅��w*�J"�b�`|�\B��}P(�Yz���
O�	9J�Q)g
�EQ�~�rB���5��U��W_��)���[�0%�(atx�~�-5~(Y�s4��b&��i�ɪ�Fw��[��2q�� 2�$=����ϟk���Q���Yi��Ѓ3M*�!��F��)i���O�ݥ�5�ps�>Q�*ͧ�-us�􁋉�%1ʔ�Xۺ�}Y�e����I�jg���؍��9��Cykz@�Ҳ�D��'E��
'/�v.�z'kq�����y)Up�1����c�%�Jl	8��+�i����b#�rXEJ}�!��\��9\�r�^0���J*�b�u)�5��,� /����YN�bPg]�*�g���v^G�`"��h'�"�tN>K)�;c���K����Z����]�5�x��v�Y�� ͧI�|��b�T���t�+�g�Ah���$���VR��C8���^g�!��.�-2v�s�"I�$)rX4���,�E�"]�j�6�8ڔ�S�$�5b��˯���.��Xp`�iwo,m�\�;av� cx�/Q�0���3?�&�/
��b0��ޏ?j~�O�H+��+1��V�� ��{��mq�ޘ�B��U}�����`��s�oX��p�����t#.�߳�q�]���?���1�s��/���H��9(j�u����\�k"���F���]�������gH���H+$�8�z	!_��=��K-r�~��L ������씥2!���X��p���߯r�f����B��˰u�Z��s�%���L�$�	~����:y0C7}��'���Vx(o-.�MU��w�2wc}Țz�?m��5���?�хX�@�F�,&1fY:�b�vg�����M�zB'*�,�A`j��Ȍ�O��l݉�������YtG}��T���� [�F�|O�KU�`����VA�!B���9�U�n0+����1�蔗I�:�t���!C�	���e��r��f�����6i�:ݳ���yj�b�!>�T���1���v�i2��J(^�'p����Gw�5f��p$S.z��'����$��f�o�����ԗ��100�s��h��6��`���uB�3��5�B���wrM��O���Z\�`�L�솶��X�qf0�CWPR
c����Q�9���]�H��O� ��[{TJ,N��k��O�^�1ڇ ��N�,��T>�`��{��Ȁ�\�B�CC6�n�/���	�k�A�cV����q-P���	���q���r+�#�c���M�l��|��:Vkh�vG�H�Ē���f���<��f&-����Wih19U~e��1X��Xv����d�"�VuOhv�΀���<O;���9�W���8��������|B���eg72u�_�\$���c�_�y�Ն����yѠv.�������PS{,�+,�6߼^;��\���0X�����h����ۀy調i�I��CyU|�����c6iǕD�	����W���,/�fR�ʺ�颱�~G�l��ƑWT�8���(�`D�N��i3���}~G��u����ɞOǱ}��T�g�ɻ����l�3���|k�w<��	����5�V�YrIߏ�Pa35C�-���]Oj��tȮ����p���H	@L�u�u 룎�����^^�|�+�|���뇙����y_�(%���u��˻��b)�X9����~�U(^̈́k��g����ծ��hU˄�Cǽ���
��]�@ҵ��&v}���3�$���wP�8%��1:r���1ǁY}F(�I�+ܫt$�1�ñ��lfh����ؗ�e�ә�$�RBυ���U^����u�P�� ��Z��-_қZ�	��r��
�A\� JrY2���-He��q���`��C3�Qu䴝6%cXla4L�P�e�"*���&�<�T�X6g%!���0L�)�hؕc@Vw�xT�:%(��`]GF�5Q#��9��i׈ms��鐭K���ο�/0��X:]�I�J��J�5�����O�f��UJ@�o]�n�t�b#I���"dӑ	��B���N\��L{}E9��m�۽
������$WtA{������I4���o@��CI��@���\6���@��*Y���1Pl�&����61W�~oM#�T�T��B�f5�9l�_�; l�6�������w��f�U�<V�OW]���=pp�Xy��� ��XZ�m�IZ�AcL����3ٴ���U�4(hg\w �d�9��D�Q��i�� c��o���_&���_$֟P��l5��Б� ����-�?�o�-
�P٧�)fe�@���:s����ϖ�^?ndG b��g��`qm�ߙ&%PF�����f�I)�r�����=7�cT�ϲ��`� 0/�8f���=,�3ӽ��e�ڽ>�]c����P-���Ƀ���$�����w548�X�+�7-�+J��j��|y) �M�� #CzDQ���A��9��� ��D�IP�}��c���Tz7���:2N�	=1��769�������	e&����@��m�v��VP����l�����bg.�<�R$�\�~eL���w�~f���*�2}^.&Դ�a������ΘΑ�!�+��YӒ���c! ���=��.�Lv�훹M� �;�Ab�B��M{a��h��ӜG��?6�;K��!Y	`@��L��g�BA�3z
ٕqa�/)d�!P�$!D*?޶v5�p$��o� &4eOφ	���������bK �E�2��.H\��.�CB^.3!���Hă�]h���m���6���9��9���IqI#�7�o�o�}/��H~��B�US%r;��vr�jY���pς�GZ��n`��*�9!�5J����z7
�.aJ�|�l��1&�AK�rx��\���eHD$���J?T%4�AS��!�,��J���S������\r�8܀꬐�X}4�f��5C�KHg���B�@�Y�%��Л���'��nc��ܒe&��Y���e�w�y�lsg�`j���Zo[�\��J��\��Oo���?�`wz"�I��iٮ-�Z�ɀ���a,�ֱl���	��~8TKޤ�IW����4d�����t�iL�Ei� I.�F:��B�S�����g�T����A:�	ٴm��Hj�(O�t���hM�l}�����f�"=,Sȫ��xh�CMO��������.��^U$���e�B	�")Jx_2/�|���ڨ�I�H$��z�>'� N��C>.�*��qt$B[�ssE��y���Z�Gѝ���F(�������MIe��7����\�҃"���CO�|�N�5�B�w?��A�ɚFo)�ujk�Ǖ��j ���>�57.�*b�ދ��O-^�Z�:g�/��,�(3��6�\ɢ�G�+�-��a�e�j�{[Wݔԯ�yp�@帿����o��^C����M�Z[P�a�V�4�������F(7?�6��%ߎ���TK��JX��5� ���~�x]{��\c@<	ͬF^(�a�C\�B�.@|��0yJC�^# )�#�Ʈ�/��:� 6+k$�>]/B�ԩ�������Vn��|�dn�����_��"[$��R�����4Z��O�"Ck3�8w����';i� 4M=��%ȰGRyʥ[��	u��^&�������pY(=�0� ���j��$d���~C��8�.��7+�Ur�:\�O�?~��r��D�έ�:'w;��n-Nx�T1C�b�P�d�+�R�J����L3M~���?��2�g�f;VK�㆓��_y~�	�`��g"=Le׺���|H��h*�� c�ԇ� ^6n��j�a%>���ԒY�A㚵#gH)^uJ%�A�����C�%[I�<��&�<�@��J� T���ﵼ(�\����o���K��/	���(���P������W"��&����2ʛ#MF�oT���V?��~og�d�S�L�j����}S���9�b���/���u�d,}fӢH�;���(�7��/�t��Nu��ncN�جp][ꕇ�7!֭���u�*���b��՘
E��N�_�7Z1��z�����Rp�XH���nK�l��k�©�s������)��d�ߛ(]��(|��'��r^�Kd��bg��A��dAj�!	{�ֻ�x�L*��r��"��i)8�"L��^>��+���jN�r2!~�_��a"Yk����- L�1�v`/�Ԑkh�?��O��J9�Ө�꟞�3� 7��޼�v3�����P��}�0&�$��X�Te1�\ȱJ�3R�EE��E00�F�MVl���C>�l�U\`�327b�i��)��y��3�5���}F_��ŀ咽��`Ԭ��U'4��Lᜬ�p�Z�7+O�=xRo����"�"�qz&-Qsڐ69��l�5�I�J��1��!b6  {C���JBp����&��a�e�~5��L);�q9�:����<��ĳP�Wܿ0�W ɜ/�9��'`�G�� �#[j$�c��[j�L>ɏ���Nቼ�76��D_~�w���W�|���3y��k�/762ڌ�u3�`�&O��	p�I��3PE,��u°Ǐ�K���:�h�e"/�R��b������(��v�W��O'��Y�0����m������@�~,zyg�p���S�_1:ŃD%r~:���){^��dk��l@jf-�n��8~��Ow��s��� ( )[�/�2�7R�A�7�����mx�qV�$e�����ūӔ?�+��O1������_q-�3�
�GΨh:�5?Vo�&���i2H>�`�M6&�����ki,�y�3Y縷W�����n�x���|8�d�n&&�)"����7���{��Afq�+g�\�Ç��EUDׇ5���M�O�l�{%�Dt��]�p����h��C���iE�; ���M��j���(ʯ��7|/�kȶ)@?��5n)����Nǹ��/֬��'��3T3�+F�r�m/���*���� �G%�����6p�.2z��a���ƶ�wc��X�v̫�=��(ͽ�\H�#�t�h�13�s��ε�����X�����oD�3痓��H����8�u�l�Ն�*㽻�"���s�8�>1�盁K��@�g���<d��2��&�7���8�5X����[����5|4I�����h�WD��`�y T�1��dU��x����E�n�\mGp�ÍJI�.ܒ�o��6��'���d����'��UA��RL�����og�@@Y�� ?=u\�H��g��Ԥӹ�Er�}���^�z���� {O��o���7�+��(ga���^��0�7�z�4YR�_j�,�%�����j��:��ॽ�MJu��$/C��O~*�F-�T`�Vq�p]>��E�����Q`����J�<D�Tm�I�b�e����r�%6W�e'R$��ʮ| ��u0��V�&�s�+e���$��	�`�R��E�V;^�������J�tލ��`�������D�Yh"n����U��׆�ޜ���l�Gb��)`ʍ��ב�`��g���=
�8Qo<�y� Nέd}���>@�Q�����o-���WI,M�-+�����3o����] d:xD�x����iM�fOΤf
H����P�B��(a����o��H�J;�8�ܗ�@{U�6\��k~����+���FϠR1�H8�r�[@��[���_'��x��/w�L��� o�#\&���r+����H�M�}��ꐲM�����2L�@��Nx�j /"B�+L�2FR�l�p���`����M�K\�l=%�X��S�s�P/�4��9��3�np��z��4򕭏�?�-�]�j��]c� ės|KY�ui6啃c�.�H9U�Bŵ�^�<v&[���H�Q�ߑ�&��;�Η�ѸL�ۑ�= u�^/T�uw�m���`I*�j�P����b���a#ƹ�X%k����O��ܲ	�i{s^�k5Fs��௿�	7�dZo��%���o'˶����jo��D}��W>~�/�k�N������bu#�4uRºZ�R1f�c���'A�������Ń�J�^�k����B[Ur(��=�ЯJwB����$��	c��0J~l����$w�+�(R����H
3���T�JzT���s���:�r3�Q�2����9���F�~7U�gn�P�G^m}�oZ>
�^fl0����P-3��n��c�"[�pj����$��ü���~�g*}yxH!�V�tQ��fAٶ]J�(%8�� ��@�a�諶a3Ž���&��������<	)d��,��*V��d����Bk���wW���k���GX��1 q�$�$�%�y��_�����7�j��󚅇-�0X-���X0D�d���8�F����Ok���+�S�_h��k�_EOd<�b��H-��[$Y�7�����m50�n<�U�Q�.�'�A����ɼz�/�U�Pώ�Q,�J:�ͺ�I�����q׳s�&�&{���	O�w|�\�|��綂K��q�1h�S�������e�����?]9B���o+��Lw<�Y���{�.x:�}Se:|�b�܌>�A�0��M1o+�Rn�i��N1 �[l���|���4��i����h�QPE�����v_5�YfU��˅
�$�S������[R�G�+�yȓ*?#�l�~$�7t>�_VS,ߘ��z��)���x�� 0gk�g�g�x8�C�#59I0��RO����~V�I����O��5�Tӱ@�_& �с�'Z�Q���D%�o-t>nf��i{Z:�ԡ ����9�j��j����M�2X{�N�\�{w�f�o�t�H�y9�J2���A�#0Gv��S�� �l��Q�a�B�3{�N ��t�1�R�k*��bM���?�,��rj��J5��-gTܒ,��>�F>0f�\I����c= �uj�$�q{��� ���Fo��U�wMD*�y��T�4p��mPq��D�.R��a.ֶ�n�L��῝�K ��*�|��rh�>@�G!�N�X��,䩪5U�y�e=N�'���|��������)dƦ�><1JT��Z"�jIw�k�3�*aW�D��le�Ȟ2P�,Kx�k*U'ةP��Dy������ۻ�k1�#�	��F�T2NƠ�[������z�{�N&��������](�3�yZ��SE.f��v��Iљo ��ǀ���:tf��>�M��������f��Ykގ7^�u�a��������2g���o�kmj�j�����E�C�\�fiU���	���w�
32H���B?�N�L~��DV�Z4CL����ol��:���C�t�m�� <��p#1�ӵJ%�[
� ��oΚM.�����}ϊyUsAhsӢ����/f�vN�S*ki��.��%\�Yv�֔�C�����fF��$����T]�YR���	K_K���.�f\�J�lw(MQ�(Y��'b-�=�m�0H�݅�w�\�mMO����mAE�u��|,���G�X�M���mWޚ�����O��Z>Kwb��޳�q�A�BFB��!GL��+}�����o'��{O��Vc��$@�L���yޛ{?���0�������S���X�1I�^�o��2�z:+ ����v�A����[mPm�S4�K{3�h|sK��e�e�Q�Z�b4�9��t�,g��^n�b59��'ċwu��aY�u��ؼY��nn������2Ow�P]��6Z��e��= �4?��j���vp�i�i�|���J^���_��ڦ��e�-��)ss�
Er�[T�ĩ��jy(Ӂ�)��=���cHv}�Ȇft�s=�w�2�	LYR�k�r~��wͿ��4 �߷h }&:�0ȱ�(Y�|>T�-&!v[�/������T1�u�'��l�i?x=�T���2#*�$���� �����a��zM�|�Π�x#��s��hD��Y���!.���Fr��&�]�+��c������T]�D�s*�W���6c����)F�ڱ���Vjao:�߸��:r��Z˗D��ژޠ�0�70*XJS]�g�ë�B��՟�L��Q�Z}�l�|H^XDݩ�����h�x��c�R8 I}����]���5�֤hmx�n.+r `�s��F���u��5�ӃO�)��*��
l)�訬`��:�m<��2�1�������kcY靺���S��y�9�ш0We�!���!��'��m`'6דU9ӒCłhro�wj�+~�2����cP�����3��zfɳAWn&��rm{a\��c�i�[��� ���(����Pb5�o4�n��2�B��be��$���T�VfR�^��&#߿¹5S��y|*�d������PLB�+��֑�A,�)á~P��9���͚X�O��P��t$�WGr���p��oʛ�!@�U�02n����v��s�a1j�/r1�o�,?{C.��;�+_�#L�v��Lp?��)�q���mi�P��_%�FvJ_�{f�e%u�X��j-Nh��{��Q�6��T�b[BJ� <�f�Ht��?���"�c��8[o�+��a����.^�E���b0������d���TT�K��Yq,Š���苜��������;K�o�w�1u;j��JĲ.W��&�	���!8���[��z3��K;�i��QL�(�F�)�El懦��I�v���FW��@���y��*�\�~�m��Twm����O�dK�����9c=,J�].��ðp��4�q�t���A|d�c���>�;����X��^�-|_gH"��"O�tX��)�^�ˬ,��ߏL�h����O�p�*�m�@����8��$�v���IЕ���V���2ĩ�	υ��Db99W-�
��B`@�b?;��@f��Yl�R+Z�9��K����8y�[Ь�J=kW@��_���i�?��Q~�D�9c�����c^]6OV��O�T7�k�N��*.�VZ��K���q7^��m8'
���� Ұ�$H���r%����a�2+�F��rmg��ɾ5ց�g6z�򂡞���_��Pr�U;]��L�L87����*_�������+y����U�K#R`��J����ͺ	菌E`MʵoCS�-�~Ⱥ%%m|i<�ϳ�Q�1
'�G;��=ޞדn$�[��ʋ�R H�M��>[�^���ѩu�����k7�-?��_෾�BqՄ�&���%��6XrVgz�g��I�D�cp�N�L����Wvd�~?!%G�)�%�'z���-�
�0��*N��T7��zж����_��3rI��:����\׹p�ئI��B�b�>�eA��Ӣ}�!�N=N���<~یo����q��Hc-�鐿�ŞqxY�7]T����D4fD��r��Z�b� ��"�59qy��bh��G<�������Q)��^6�D��z���Y`=��GOi�bTI�½���|���I@_R�ia���I��Z�X{�Jw�N�
��8�7g�a'r׮�K��WP� �?�V��v�t��e���(�EQ�������<�����A�3�5��� z��uf��>*&����H����sQ��C��]'+Ҵb�2f��F��Z`Я=�),!s��O�Q0����+�z�W������gy��PG>�O �o_f0P:���_��w-�ZB�C{Y2?�,��攘�l��=E{@ah�FeB���h*���yJ���/q���֭%`n����SY.c���-��L��-q�VyhP��_u��:�F�l��ц/���m����O��:���гＯ���ЃUd��*1w8ɸ���;&��bH ��R�'�6�P_h-h��ꀔ��ݢnfE�w}蔨�7�s��$�mu���E��T��\P� V�L��	��u�z�S��jOy��0�x��F[YS�������UFھ��B[���u�D�?
�IE�<t7��U���Z��x_.���Fਬ9�_iq�`��kZ��{��e�o��> �4ݑ@�����p�l"iwV?����G
��-%��z+���~f��� -D��!&p��6��HX�nH:���=�z�.�Cs�g_���V�8��1�ro|����zs8/A�%\�'S8S�.�c�\��=��0���8��0����<�`�N��kkI̙��ᇧM;��5�-n˸g��]����v�Ӈ[�~}�Am�)a3%�hF"�X�m<'�@bEN�a�`FȰ�n(V�oO,��> 1׼! ݁>������?���Q�#���&G[�5�v`' p����w���	;�v,�ѿ����!�J0������bK��E�H��n��Iu����������S�T'��!�:ҳ QOP�8 "`�3���^B���s��-A���prI�]�t�!�٩-�uZ��UXH��YuZ K�}6�B)�QU��}��Z/��18�"��(�\c���zhzv%0��ô�C=����W�	�9���1=��  Hf�H�G��r`i��o���v�p�I����/6]uʒo����?��
�$�ŇtDܨ��ϳcs�,�^���y�[QM�r'�=��۱����B�z����O[]�Ji�����U(P���,~�/���'_�*|��:�r�4J���A+�AvM	(����m.z�I����X�чI��^���$$]��`���	�1st�6>[�v�$7�-�&�&�p��4҃�L�K5
\��6R�L�]�5%��KZ�7Y���-�Z���ӳ��v��þ�i����ꌱ��r�e���	��9�L6���!Y��Zc�Hq{!�r!P�[ޜ��Hv�����H(�yV����s�z��Fm�<g��')s�������4�O����F㳈�J��Q�\�?!��cMl����~��o��B���$������@u�8�$"���D����P�O�e�P-���y�,���^g��}��;{����)��ٯ݇5�"����:^��}��?��oS�?�!���b�6�+r�j���b
l��bo��r��k��a��K���9��Gf����i�BI|'��c-������eəB�_H����I�,#�l��PU�4���*��] ��fy�L^s�N�e�+q�.% �>\�0�'�gh��-���N.c76����fJ:����Ů�"z*�/�8^�2ۉ�p����+͖,Q����Fh�Rl���˨U�0#��@�y�_^�)54Y]��w��P��7�'�#2_��1Z�A�
6��_7�^S�m8N�\/˽�@� ���B�����գ7�m?dJ΄��a]��6��@���,i$���R��}�.��#�	~k�n�5uz�M�O@��)7������:�f����_�����+.S�Q���R&������>��BV&NO����j��QË�2����u���YR��'��� �Z�D\�Mn�$�hyc�!���Bd!LG�t&��?���y��>�n[o]���3p,[��0y�f�C�Z0�_2i��N��H�Ȯ���cV����ڄp8vKЃ�ھ�S�t���IsD7�ɷ/�cj�����(}ND�1I@�Ǻșl^b����SWOh��9k����d=⢀fK�*a�k@?���4�F�m}�����c1{�1@�QA�9�blY��Ņ�����G=������y܋9���H�ӝ���.��1<����
܀�<!*�05�vV�&Ժ�aЉ����\�> ����:Y<}27QE�q.r�G��RU$� '�-qWt�^H�]�t-k��,����f5���ʦ+�f�굈��ɶ��mH���DIr�o������"�EΑ��3�=�p��:���	6=ʐ��c��ia&7���95���9�9|@C&;h$��+��E����~��`˦R�d�Pթ`@��S�mog�� ���)s|Ipu�ＭF t2`V��\��K����=`����pu��R�$ٜ�k��Z; :�]�3�C3%L/I�C�����g����&���O,U�"�M���`K���z6�U��X��o�:M�i3*���ڪy�ٓLH`<B�����خ�{-�C�:��-����eL؝'�!x���Z/�=u�l�.�c�4�E}��.m�z@B8��}���K�kl�g��|�q����(�l��`�Z��<��<��^r}p`V�$�gء��9aT�xM'PX��y�6��Ճ6Y;D	1�w;�ҵ�h',U
r���(����n8�N�
��{��'"ygt�I�q�ù��q0��Ue��F���~����j�Ep�L���Ҏ�1l�?DL�z���1"gpy��:�ftX���߹��VC;�_����8Q���t[�����sS�Pw�^��-��FT�7�hn��{e���=4�%��_�ng=���3���@�˳>�6��,�������橣����(̢�T�BM�H��]���`���a��5hޅd�uv5TeW���s}{�#����c]��a�^��n9�B�K�	�j��~Ώ�=Ym.��$�,��[��Il�IZ�@�)�N"��H�Ϡ��'�2��8�ś���b��n���l���Y���U��z�N)��{�m;��*�����ʠ�z	!�j�J^%�|�4�
�p ���H<g%�7�Fc'���Ѯ���3��E�|=������
G��e�$a�ƛ</�؝�֖f���2��-q�T;��LK�8VFg��؎>L}̫<E��N�rI�Z� ��f��J�#�iX5)֌WX64(����i��4<�7�l>%�O��f��}&'K�BE���z$�²�(o�_��:��'��Ŀ\���4�9޸0q�L,�E燓�1��5d;��$����r�:����Zu�a>��ZUN�Eu"O�����]�Bf�l9ޅUH�-�1�|�)9��}��-��=�Ϫb'ݦߞ:�~BPk���zY+2<�&����aө�c�y4�i���R�S�X��!�w���	{�L�n�y��`�0�Ʀ��j�8,�����5j �ɋV4�F$�"�F�o@�-�ڀ�p�=���-�S���ts8�s(ŉ&B��E(�
eE�L���zIJ���NL�dm�����ru$�_�;�{٣�zlK(�����w*�{���h�얀���4�. �C#l�8L��d�#���Br]������6��]�\�4���y�Zq�|ģ-uO$������@�	�B{&&�t�[AT8���,�O���[SG�'&Q�ؕ����j��������}��=8���[�(λ�� ���ZG�+�y,E/�h��^��Ea,-�F'����'jz.sz�k��x\+a��tt�p����{��:65�{�MN��o�5��t��Н?��a�1^gYN��9K��X�w���b�c�WW6��-�DFjg��ҟ.�C%t�M�ux�Yl������q������-1�-�y��^�$�����p\����0�3��"��%6�T��O0s-�Xh�>��iVW�Ƀ����S���Rw*��ڃ'e���o��<(�czr}�ݱ��_$��P�ۖ�������us�N�
�_L���j�)t���V��n��}Ϟ&�ȇ��Wkzѯ�> }�i�~{!n�f{���e��D���Hvw����N�
䁁��)�L�C����A��k��Q��̠�'l~W٥���&�*qML�SI����d��n#	4���9.�n��T�b�����Ʀ��Kֺ�	wB�9��{1�̚�2�W`��&,\I�y^����}$���лn�5M�=?(��`B#�+��}�7-�{LZpM6������jľ����ԇ��:h��@j�-Ni��3fK8)[4$4*O�QJ�l���o���]�dށ�����ϛ�DBSS����/?�}]�k��_�_���&wI嚸ι�ͺ��h�J�B�0LM�rL���!�:���6ƨ�c��t��ZD֯J�������	�Y�KҔ3���*D�*�T+���Ge����?�@q�|�Ձ��z2�>������{����� �֋���qc~�HY�Qڋ��ʊ.Жi�6�ZD�_�oq��p��`Y�[�j�z��Ps��PVrts�W0����V�E�?/�B�;c���}r �d8/�s( ��]O+�5��+����_����+ßx.���O,�r�� �0Z��5���>\�4�ԃ��%
�|�G!2���C]DJf����fh=hH�>|�	^�9Vˇ�7�#�z��� ��>��g�(��u�t�.�g��S���Mש��l����	��B�, ����3���Dx���>��;T�&�.�GK�`���4Ǳ�zN&^	j�������^��r����BC�v���5���
�?��~ 1���N�U�����%O�P����pq�.�t�*������o	��V�=��1������ ��pJn���z�����>�!�93���K3Խ��S�Vq��q$��I�
�6F!j�HnP�(M��g؈�x^Pf^7Lj�S�����h���r&�XJ�&�_1��`U�9���Ͻ�7�?��	��;'��m=��gvӟ�K9�����8{�G�p��˓T�>�?�^"�p�tfGK�~��������r��Jc��� ?-3���g⼬�vK[FOqV#zR,���� �ߦBx��|XM�������U���s�J�z0faj�:?�R
����M��k�l̋Bw;@��r*� M�3��d�dC�t
UF�^�֋F�J�恽ij�&w�Ӟ.H>�.E��M���PpvN<�_ʸN����OR2y�^']�!���"��̗~��7⯮��K�M����-��,�v�
������AOo VϮ�8��cUG�a�/�f &b��OS��nI���!]f3�������d�"��A)��<����\hXFB6��`�U��f�o��I��p'����V�BF5�v�Ռ{��U�1p�b��^.��x�پ����DI�����UH~4�K��@�^r�i�r9:t�"���jhE1��I3<.�q8tK�59q���X���e��Z�`�ˎ��.2����g����-`�7�zT�$3�m9�ELw�hqef|�{AO�JC��M���ZԚ�(G�5���/ �
m�����ۮQ�c�/��h^d�N�%˪ɐPÆ��璷�ГtQ%W�M�	�Qp��X�4vTCX��湯0��$[S����)��ä?^R� �HaE��?^.�x�`������7�?�L����I��ŉ?Y�p}�hiŽ��F�Uy�)6暄��N|)"�cv��rl�'7�l-�r!��E�"g{i˝�L=���/g��Iyj�YF
��l�^ƣC�;�[�Ϝ[1���%�쵲+C�J(�܅�[\kP���%I��!�c��1��L� z^Uս@'����Y���H�����.��.w�m�����	���Bar5L�^��K���G�������U��Xé��V����n���W>�d�>Z"��q�}{�2�.���KW�L�c����]� �1�O��2�7���h��nRm�e��#%^\i�;��"j�*F�_����3er��']��:w#�k#��ŅIj���@�]��S�'�������ˈds�����=K���=���D�k�Ã��{}�b���ZzyD'�ԧ%#�1P#e��R��7�q���eq���E\����UC���ջ�=��d}6�a5y�!��E��)��<��Z�\�b��zW��z� +Gt[-_W�̡ΰ��R�&��������Si�ӻ���8$���S�P"��QG�st�Hc2�>�l�uNo"C-잾޹?qĹ�>aК,�*ʎ\
Pq��P�C�6��Z`*����*1���~44]�B%@�XڠV�d ���|� !9@�!T���~���$�}�7<92I7?�zDj�tE�T?u���c� ������]��B�2��Z628O�L��q͍���Z)Y�}űT�'���l=/�~u?�Q`�eUˑ��*	�	"
�g=F�j��*	xL�����CN*d>�?��g �3�G�TZX1��i Ju��9g�͌TW�L�
<�Z�c�XOh��~�?�Q���o��O�
��{�eCp��L����'������
OGa5�7���V���»����oɤQ\�@ǉ����@���*�Bjfe%��]�(��k�QuЗ[��&�o��x�]X���jJ�_��oE��?����s,:[��
�C�רn�
���s��R!��X����=8�v�+��V�53���:�H�>2QbuV����F�|��nZ:�������N�H�~:)�p7��M:�ɥ�A��G��k�i���z�R�}q��6c��=NGRk5`��v�>_O�
i�?����L >�c���'�@ŰUY(�/�_�'1gd���g{/� ��w�)N�3xoa�.��Ң��\��*I[�{��;�{ɳ�F�(hK�J�����Fu�=
��&Ϲ���G�� �U���#����8R$�ǒ�OD�;WW9�h�J�}�h�����Vsϟb؈�J�F�0�);^J2d���X��Q&����Xl����xu�K�r���4A%��/�#ښ�5�#�iG�;<��5�ǌ��<~�]��C�kB���4 ײ�ѾT��r=��+y]���C(C7��1�����uD���r/hr��vN��߂�Ҽ�C��k�ı��ұ�"U�hg�4X'?���(/+����g؟��fo��+
��B�i���B�;���h���o���810Q$h��8�Ic����ߛU('�K�&�R�u��
�-a��f�����x<�1�ϭ3*�����Xr�� �q����ۓ~�趦O�w9d����'^��f<��A_VꝨ���>8 -p%os��K� �7����g�{�|li�&�5�8߆�^fv����;L��8�]��J�:�4z�����6�7i�ϭ�ӭrC֖��@W���� i��������}[�h�����9V�%�'B�R%�,��,��xZ.43�ħm��u���bW�dq��f��o���0�cqq���-�<��yܭ�x���ھh���F'U@�w��~��������~��{��c��wI ��g���`6��H��-������7��龺��XפH��q�Aס��������}�m�>[�X��u-5]��QR�x3���+��ef$N��z?��Erv��W���`U�D#���}��.��(� �5,r��щ	�v��d6nd�0��뾸*��/����D��B0�����Ǯ�qRIO*�	d�� �2��V�������� �U���M��)=No�1d\õV�I�Z�f�u���	��g��#tT@V!�X��T��tu5. �s��� �����R=��!�DC�9X�����'zvDQ��i|$�Q���TQ5�ܴ�����f�����py���(������[� a'�;~���;��H/�)l=�Q�� �5����v�����A8�@�.���a�������ho��ʬ񙛴{k'��SK%���a�6˅'6�����[V�f�OT�?X�"��3y��u��� �0�į�q�Q�Cܬ�)��S��.˥�.O⎵�cE��AA�{�W�&��0|�?��q�~ة�e���)���t�=�����UL��I��p��u)7�
f��vY9o�Q�;����Kы��H�5{�w��Z�W��8����y�[qG{*A�p���D��z��2%]Puk�?�,U`t����L�f�K
pEᲰT�X���dg2fh@Q<�K���T�����y��pX���=��ޑB�+�-�����?F�G����6�'�bͨF?��|���X������c���~�.�<_܌2m`�X����=D}f�R��,�7���������%�C�%⁦6H�
[��wG?�!��іE�[ �_�m���^�Wa#�E>D>uժ.���"D���NB����;�s���5���t��pB�XIb6��ؐ�wY������˖HZ$	�k��ĚT�O�pZI�e��Հ����Zk�UV��� W i���sDq�KG6�pf��	�GӀ1,9��IӦ���[_�6(�����Tۥ���Y�1!�"	6S��Ь��I�L�l�	t�4�!��1H����[�!�w��Fo�$~\�:���iZt�`N��S	�N�����Ʃ�`x�b�w� xϴΓ�K0	�y�w�M�R��ޜN�\�w�u8����k��3z{� %o��kRN����)�Q�r�5��IV�G��&3"��7t��ی �zq�k�s�����M��$5��5������*����|O�~�M���tēV�Uʈ:�J�}8<w��T&�z�&Iq-���Dr�6�_4�T���n�f�_	Ā�+���A�tGJN�Pi^6�&z��7@B�G1>yXJ��y�fu�+��������`��w�5��)^j(�[�(�4����nN�3���-3l~�߻E�� �&�aq�wW)��'�N-"ŕ�OE��7p�~Ϳ��� �5�h��B����a���L{t�Ň���}���_c����꺉�N񔔞����d1p���'%aXz�z9�$(/�=��Cb�f�<��sdR�n��7W��=Us��7x�1��Ez�P���[��e�����,W4�~hc`��%�g�IXy�ɐtr���t�x.�}-@�@�f�
��_4�lE���'����Z������k�%g�?X-�:4�9�h��}Sp��?go�V�xS���Bl*�$�?�ĮGz[��SE�Es=�]3�w�d%'���F cVb�$z�;���q: �?��$���(�r�:C�Tb��F���0���[��B.��^�4&L.��8*��J"�Ǽé���[��k���`��!�i���w��ů8��EO[�
`N�$6�����J�X��i:���`I[�������tgn�2��A x���[�Vl�>gK�f>��ֽ���X����j��"<ĝ�	oΔhwe�oLxhN���;4���'�l�%�8�f�{[W=,�:\��%,D=1�y�Ifr�e�8*#�16��݂��>5آ���Amɩ�����JpDU��s�?��'���^{݆bl����v4::]�)lq0y��"�Iml ��z�W�dT̮OI�H�xɯ��h����b1�eO�:�����FXV/�Ml�R���`'d����0�I�5T=Ig��'�͐�h�ɏ0F��3V�W�3�Fܴ_̑I�e5�tu���E��<A��w�݀����1�5��j'0�}�jVk�m[���*4�z]j,��(\Q���o\I�4�+hD_l�dY��Ex�{�h\z������SÿMQ�	j�Dv$ɤV�H������B(M���d\w�>JG5׸���z����hӤ��M��~�B�c+�j�L�� ���ކ�΄k�����$�PY.Е/E�����"���rK&UjE��=���R�?Z�����0���3�w	��ǻ;4Q	z������̥�F��s��*�]ם;�_J'����۶{湥�\B?�}^¯O ȟ� 	;w@�>�]�J�i�%QqZ�;��zl�Ӳ#��i��Er�@��x7���]
�\��܎�v˄�v_tT_��&��F�?�?nyB�?�_`oUu0A��qp�K������*$̆�Oi�R`!_�u���:��w��yb�������hyj>�?D�&�Q�#[&T��1_u�jL��,�����Z�/��%kQ�OŒ����+)U����� �a�4Al��_��S�;� ���C������Z��Y(�4��h�
���]輦N�I�?�G�;ݲ��x��I�ڒ��n��Q2��]e�����8r����H&�X����-5��敩�6S�� =�L۷I#�B9���Z�;�I?��J�`���q������M7,W_ �|mFaUl�r�� p�>@~�*��JF@Z'�U���V�ع�M�ڹ�uY���硡p�'�����%��( X�Ӎ��z��	J�C{������CE(�ާH�3�i,:㧷i	N�>i����.�l>I������}�����<�ֻ�V�X%�:?����Ɨ�u>k�3o��s������cg��tw�l���E?u�d^�j1�8�B�2Zc�V+�K�i���G:�48�|M���1��20e�i�!��� ny�ŷ��]��s���=����Y�:I`@ �d[�X�I om�z��-�=�{���G��QE�bi9� ����T�<:����������wU|sْ���ݨ��`�'�V�O�?D�� ��K��j��Ѯ��µ�l�St�T_��v�3�Bl��<���7-�v^�X���E3�Mft�,���|�6�F����*�Xu�}������~����t�;q��oT�!��r=(����R�d>v�ui���=��1w�
R[:�?��Z_���3	8h��!k7�����s������O68��L���Y��c���i��(�;w�n2��;uRG�k~ x�KU����}}�B=4j{�/D��p���>)��W�A4����I���Pۑ��r?�u�k�{��$�w�/�W=�4TVm��?g��Þ��� ��^f�1��<ö�q�ɸ��_�܎9�]�Wz�Hy�@�{Mq��6�:��T��樂���&��ς�@t�L�A>,"m*�f����{栓pH��`�C1�ܔ�}&�r<�M0���h�8!���lf�r��S�����g��ĥ�?&d�| �&�yc;��Z�-�+�?�j�l��ޓ-�Ƒpw�����w5����v����eR��p�������k`�ӑ�,2z1�\z�>m�r��M�7ڹ���p|K�^�w�%�&�{i�l+��mS7��6��<YƮ�
���u�2��j'XS ���,�I��
rI�Ǩ ��?���ĝ�&��"�w¼�i|]�y�\��h5_H+}���<�r����ӄ�W#�n"53�	M��������XK�e��}�W8��C�l��ĭ�O��'m��W���'��k�@�z^�N�E}z�Ro��`�H@MW���@.��D��7�b��om)N=��b�n���ڎ
�@�(��3dZ{�Υ�N�[\�1`j\����ه����ImB��9��ktc��e�����|�xNs��3���Bp��>�J��X����[��qE�e,�$�|��2���G��̧��y��������*�z^m2a������g	d�ߍ�m�0@uf�`�7�.�D�}��Zk8Y�f�~�2*�������L��v�������+l��#��K�4y��7O��r��ݟq��I6�	F!��9�a�;4�P!�P�U��4�!/�"�1�I:vA>�����2�a��="�	�cM��Z���1��<�]�6J
���u�Ia�n�	A�s����ccBc�ˀD�ik�Y���.S�2�Ėa�k�m�2���]�. Ζ��&RUtK��e�!��A4���\W#�ѥ���QM�P�ǔ�d�Q��
�=W�^�J՘�)�29���h���-��iV��[IƻhC�(���5`VAs�c��GyE�R� �h�ʯB*'ɯ�۷��`�4���	�[�T@�.��N[j�=p.Oϯ�Yg�O�����Ӏ<��6�|��3��<Q�Ǚ�L��^_zUg�'K�r������ʷ̾3?ole�ӥ1k��᣻%��+��*��vo�Gn�`���������m�4��O�Ņ��Iu��ig�4��/�Ex���W��I�or�Oy�|��,�������ܽ4���s��0���@T�����k)� lI�l�������)�z��$W�I�n^�-�ZM<`x� 0˽�>��dƴ�&�$@�?��b��ã�0�i�:�3Z�4�K���Hǲ��^uX�8�zi�qLQ~��c�!���/�?.��Zn~6y��+T�����~,���#?�:#A;4����@��y)j=�C�/`���N����L�������I���W{:Nd����/Ih|5e{�e��D�x��y��N��z�n{͋�D�P��h�8(V��b��BpEx�ƠDՙ/٬��8&>���OӒ�aK@�p�
��c�U��;fB��s,Ὑ[�/�U-��sP:�0G�o�V�6]���8�����!��abaZo������%���2*����䯚��纀v��Z�ߕ#1�Es�-ա>a��($���o܊��`*��ttW�1��]�g������t]�����Pס���T��h�����ſ�'����1����Z6Q�[��/�A�RX����:b�?�÷^��|찬*`D#L�Cr�4يp���n塶��/%�"v<?��K-��=y��R�k��΁�y��&=�%���4�E����t��F��s��|�O_��~�I�]�<�ݱ��������&���߲젋|J�ԏD�0��"Ao�ޤz�9*2Xs��:g�%JkQ��
�o�a�9�ݸ���^�8v���e���Kz��Jk��l�hyls�c��)S�o����OI�Q�a�XE��w�{$?�[��r2�{����ҼaBS�U(�*�������d�����+�����J�!�B������b� pU��E�.ę��R��B1T��C��m]*��2u�Dޒ�鄘u<�)���A�'R��u/t>��Փ4D����2?{k~�p�A��c� ��+˶r6<�c�?�+`Bf\����q��P+��l�F�'�q���~��.���J��6q}�'�:a�2[��&T����%�B�n�Y���<�o�1b6H]'B`�f�0��	�
�n��6������)u4���.����U[�K���kiMF�:#��v)(J���0�����m߸WzK���b�A�[f��N��]Z�����Lkz��-& \����A!1�ִ�sE@6'���~c8�|<���zmF�Ji�|���ԀE�i(M$���IAP��?99�pu��)ǋ��j���K���rh�=��J��5��O{^�T�$f�Y�#�-�c,M��������h�R���O$R+�B��C->����:�,�#g�'?�R�9R7����毿z��8e�[��A4�=���>��`�A}�Y����}PJ5�>�>�z)_s�u����}Y�+��C���;��I�}�h�����E;�M�zUb�|��ow���٦"����&�!�(u3�3��������#=�o�{�V.��ېBw��:_m�6���)c�akB��ae��~�!H��J�gԇ�fݪ(_/��e��A�$�>ke�X�${�p�6F)ծ{�=R�|燫�S�U�"��W)�_�&<�a��}����[���"�� E���W�"�{S��C��Li�@�"�p�_ ���g`���An_�j��g%�V�Α���n�*~�e?`a�~͢�*��g�U\\��Ƶ�R��e�s퍛a������!N�Ҕ�z�]|ŗzUOK�{�A�����'kG�Y��J�Y�|�~�� 6���)�ĥ!��1���[�p'9�9���RO�E9�ύjB8�ލs���<F����p���L-�a�DRd'}�#�.����Z���V���<<���^�J��ݹ���g�֟�Zڍ�Vj�,ˮ73)������4�n�5���?�h�o']��NsPB�@' �h=ϱz՝gJ(�@a�
�_��,��.fm�V�9/rz���G�Aſ��"J�;t`xG{�C�|dK���,g;'�[����5qi�[����E��,���ʗ������O?fDI��P��o␥���o��h�ẏh��F�Q�ho�A�roFNO1+ח�A������}��=�)�ڣ�K�"��Mm���<	�z�}M���2��}���񰋣�]���F��_���+���/-��ݤ�Ŧ.ld��� c6z#��w4��%�SmЌ���pW�sQ����Ȓ�o�?w��}՟6�MD�.�Z�R�e�)�F*��_���׽��kq���#%eQG�k`�O,5��|�K���p?�Q c�<Nt	<e�%M����O������������R�v^�ʇ�%�k�dm ������\�b@]��D��Nh٥R_�+�7^`��7$N����N���k�;���9�z�u}ꒊ"%�4����թ��Rb~��'cdT>w�c��Su��~b��Z���\/g�R�f�p��'Z?|R�~�B�:ʧ�4R�h$g�	VS(�|SzD#CR�.���Hs)К],��=����ް�0� jq�(k��Ե.�iFP+�	[�����#,�?�-li{�1��s�g��)i��v��0���N�<e���x�O����e\YF�h�f������Tm#7n��I?�ԭ~�=&�l)?R����KF'|�{@-�ث:[��U`7��w�T�F��,fޒ3�[ϼZ�e:#Hyh,���S �m��M?}ۈ�%t�I=�D&�������.N�=����*��+���j؏#��It�h�|���)B��ӈUŷt�ռC�(+���p��P���)���t;Q3�Kb�Ԁ�7d��,�l5�3|I���7b��׊�ƋbN����^?Jے��Gz?��}/���&�=��>���qPע��8�+�����ѭ���H��:� ���b9C���ѣX�"�[,b�,c��EE���xH����|`\0�-2�N���*�A�����a4�d0�c`"���Z?������_�3Ī<���S���@o��. ���$��7�����6V��,!�1	��pwj����4v�(N�t�h4�P�t����������F���Ra��^�tJ8�����W����]QɼN�\	�S���]�ŷ�K"�6+?$���8#�n
`���M��ݏ���-���p�� {����>�zH��.���8n�lg;��^gt�C��o�8|be���3�&����h(�����i�d��w��XĢ=)7���c8յ"O��xc�7b�^��WئU�+h�4���ԑ�����r����tn��'J���{���M��8�G>���&?:�b�xʩ���0�\�Nkק��A�<C'�Vqa��Ҵ�SH'�����O� U�D�B�u*��v������1���4.��C����;X���sQ� X��;���TP�i�<rG�RÎ��_6m����Y��LJ��ϑ��2F���2YZP	-��9;�����.b�`�(������+��3g�7b׹�?P���{����2�h���`�Ddy}���zIJ�7
*�jr�k'CrJC�(�l�U;�5��N"7R�[�������"���,SP#��$��'���z�ڜ&i!*�v�CտP:FK���Sw��(�܍Վ	F@|�4��"^�Io��e`o,)~���c����XF9:�W@�SU�RoS�.�ZJ�ի��ȼ�t0O*��Ʀ�Y��kY�}���(yZ2�z3B��=�).CM�X�a�-��=`G��n&LY�J��0�o�ձ�{!'b�5!OS�=&F��|��h|�38]"Zۖ���=������!�I��>�!L�+Z�AK+Yq�AU*� dНXT��"?�U�7�Ci�װ��.����(�wa�r�T�׶���T5�+M;Ds��X��s�X5��p�X�C_#�U�;d��",��W�t�.�����W�u�UFl ?�3�B�҆O�|�\�C�~���jz�Y,o��/n>��euׄ�g���n�1-�y��"�������-Nqt5M��L�h�^�H,��3�HYn��u+^5+^���?td���[�%c�iW4}�s���Ƶ�L>$2S�Lsڎ�Z�Q������7=E�\[͂Ŵ3��`�s�1���9��	����A �*�8�O	�P��� ]v��5J:]1��M������(���0>���Ʃ��1��+�9�a�M#��=�P�۶!��[/��p�s�E>���E���f!�Vo�d��,lo$��$��6Lj���	�|/�a��ol����}	��o)=1����Vk��i�E'��;'7b ��'�w��򚫎ZchGoRG7~��L��/��7����
9�L��\E� d�e�ny�n�Ϡe�m�A.���Y(�� �f �H�\Lj_��<o�Յ�c�x�b���r�#�yrmxF�/��K��0����lc�ִ��95������T6�a��V6�p���Vt��~��}�+�nqev��8B�@2U"<�5 U�3'b.�%���r'�r�u��"$B��2Z�J��S4=�Id$u��H̽��t��
R����s4֎(�;2Z�\����-�7E���<��0_v
�;�2��Ň"!��/��`7�
���س;���U�:�����lwC!t`M�;ƛǮ�n�Q�e���D�9oD/1��e��mh������]�|���¼4� ����`m^{�B���\[1�x���RE"�E:!L9�Wf� �'6����ɶۼ�~%�$��:�U�7&Nl��R�E6�{,�J�%�d2\���q|�W�[��j(w��ݠ�H���FW��!&ޔ�̢F
e�3�zO�d�˖_�v����Ԩ����)���U(��)4#��}R����9��`����]��}���g�S��2NE+�A�,�:0Ma~E�bHTn#'F2X�+�*,X�qnF�*�{��3�=2#��$�8�?U]rടl�+G���3�9 <b/����!�)m��ZJ�����9�py�x4g1�gz��$���
�E����,^�A0��I�C��t���3��T&�u;��h�Gw9A�����s7|��&����b9B	c`�Z>h��o~:�����m��B�C(X���[j�/-���rJ���{u�T���wa�X�/`�q[5y�M���|�le'�a�>}�f���n�`q�s�2X�*KF�� ��5�$�����ĸ�[*��F
�ϰg��� ��Mܑ�*vh!���~�Π��ʰ�IB�RTl�S���<e'Z� �k�� ����D��*��SI�����KuHW����ȳB��ns����@���)$ �y����;?�K ����ߏ�,����h�<G����襍�;\n�eA�����G�/�����v�d�7xP�[�Wm�3�yXj�����`�@V�H��]��ndH�d�7(b�V�X����K(��1n�tY@a��������=L'S+�t5�Z��S~�VUE�Ajg$3bC���L�uʌ��Dj�	kYޖj��ϝmU�<���K[�yCD���R��!��޵۸H���mFPp�r�CD�_��I~��ʃ�O�]�3!��Η/D�Mv�ej�����Cۃ�� Z/�.1RRG�NA�p���T�0��$)�Ϊ��"T�;x9��*"��-!�>eG~�/�-0�!�2%[�o?�wkUA+"lc.�aL�fx?4�
B<{SR-�sdw���W]�����p��Z��n9�y��4I%/��w��P� ��;�d�{<�u`$��2�?�֔�p�@U���9>;��nt����Sj�^?�)F��|S�}'(N�Hƾ(l��v�Y�B�A^�P��]��L�kJ>ݨ��a���V6H��48rh��> W�]5��2���w��պ|_���%J	�D*�Nf���9�s/ːx�9o3&!��T7p�}�����;p�1RD�ed$b��[����c;mvʯ*���|%�A}�2
 �km5�v�0�ǐ7���	G���o�$~����]7�)�7�����,��=�*
ٮ�pH]7��~�@�t#��7t��|�\k���[ԉ�B��
�����h|�/
}fӱ�a�2��H�)�׾�eW�j�������\S���Q����D�QB�q9ʸ��&��X_s��
�f��j=ȶ�Y;&Y���d�MX}kr?Pϒc{��%���&��WH�zK��q��/s��P6l-�Zo(ͅ����؛��T>o�\��'�"�h�i���3Й���fY:�!��O�#6����!�9�x�6�� �׵��T�ǋm^T&�u�ד�!���]���IR�k���z�i	������E���#&���M��I���d��4�}�U�k`�'*X�]�0���׹�>��8�re��=��>4g{:s'ORK[����[d ���@���(fN�:�B\u�;+d��c�����5 /J2o�N�1Du�Vԟ "���@}m�J�9Q��d����U��Z A����d��엋���܌�*�~q�MO�KbU����R�=:,G�w�Ρ씨}h	��!��4��5Z�v�Ps(I2�Z�1��a{bNw��cb�������@�[�� �`�]�;���_�k>�5�$~�v�4c���Ԧ�������;�L|%#�A C�l�I��fB�sl�f����?��(�C�2�б�m��П��e/�j
�|#�8�.�W��}C)Q���)��gQ����3�d<�ީ�F���g)~���9� �-��Ϧ�'߶>�ׯH���8������[)U*6o�.T�нzF3�QW�ڽ����N6��\t��gq�4^� s��쑭[�����g�^>���F��= �'jR]���U��^�|X��z�zR�grU����~���oŒ�s1�J�#�����Y�,������=L��6�,j7��f�E5����F�ճ����$)�1�#�p\�n�{�z�o�T�Wߍ~��J�T���ɓ�-��{$�tm���R���gZi{C�S}��S`��Ċ,a
����[ ��@�# �������l��Z��H���V��
������P؁����=��B4m�y�F����l]y��˴�==�G�j�R���b��ฦt^F���W�������G�S��zۘ<z�2c\���J�Ș[z��P%$_�BC��St�LΘ�B���4����+f�����?:� \�T|О�1ЋZ~U��¹?�[CVsm|��^������G�z"r��/ض�`AI���1s���i�	 �jF{�H]BK'WnM�֐�U�l����|]{�BNUFd�'��&yt����#��[MQ{�=��$,"m�Ϝ���w}j�ыT0��&Hd��j'^�JuF�t�o���?�`ށ\w����?��� �߿V�d�igq�d��H@����u-,�&?��
"����܄�����>Fi��y9��3X΅���J|�(X������k%a��y����e�_�_%��'�X��I�=�Dh�p�EL��7l�n�U(�@��F/���[@�~�/_�Lesy�[�K��Ѻ~&�z�I;�u|라�i_�8 2�h;I�~�QF��#o�z�R���n>vz�����	��z�"E9�Y�ƉU}n�����}�<}߲�A�6
$��z�
�W���W���j�*��@�5]v2M$��p�!r��Y�6!�(�̕�[Px}�&b�$�0�������ŚF�5���բE�v�7"�1,�d<>ĉ ��� ���m�h������#�@���9ОV$�ǡ�ȷ�"��\���/� ◹sU�	�r �n��P�	d�QQ��>`͞����>LǬ�{���)�4+oz�s���#�܋���|85r+W3�B(&u��M|�y��%*�o��q(C���k±��C�LCJ��@�J	�@�o�^�MyI�WW�8|s��B��d�pً5�)z�)�:I��ʻ�b彉��Ĥ#�Ԕ�&�-��Fx���P!���iZa��хʻ��Q�D �A���m���'���4�^xs�xM<`������rO$��;3�:�T��^�0!�͚t����UP������\Ź�� (�M�qh(����5Q#�h�^���슗fUΥv�F�Y���Ӽ���87�
�
x�-�X~�	&�voQ���O�>7�x� ��[vg%\����p�%|���M`"� m,s,�_ⷨ�z�¼�d�)	to��X��5��t�Ax�篏׾_��&e��H�qg.dq�NV,����7��l�viH`�P+R$a|5��NG'��]r��x��'��d@�Im�AjV��'� ��@�����'A�K�%L�>[2,��i��W���!|��$]a��5�5�#ͱ#6Uö�m5��Cp�~A�/���XĔ���B�Ó�z�Jx��Y*��gg�GΖC��yf�vQ۰uk�w�9�FK~	��$_�����^�BҔ~M�� >n����E���2F��E�̛�M>���W�B
��`@�����ӽSC@n'�q�w����6�c�kQ�t��5���6Pl���-��h�3�LӔVҳ�yRsΜoW=�p����µ�1���4�[���X��=+;}���H�5����l�EaxQ�4�9�Q��u/��&��rk}Rq���p]�B:1�n�v�-0_#g������x��څr����5ӱ�~��\G��s��&|��k�FM����8hQW�^\U�B'��v��A|�>�p�p��"�l� ��"1n>"�*]�|!z���:G�93\��d:���� 8�()<���4�ܣ�iT��%�]4I��_���OĆ���
#���1�I�(�oi ���#DSz�G�L��'��-	�dh@����gς��0ӧ���ȥ+��p�0��N��rvNX�v���+�0@#�}����/�Rql����74ؾ�w��<l�L��3k��"(�s^:�R+C�� uC��=��N��T;G4s�Lܓ���-�ˡ(��s2��q��/*xr�@U��߮����d+�:LB��̞(Y��в+�5�׍��(gK�]M'����L������Z�p�>o�0m��|f]�:��4ƌ)�SE�sA!��SpAK��t�)�k�=��h����?,j8pXϖ��$(kE�.��y���_ѵc0ۢ�M��A�����T+PB�r5��e5Ɲ� V��]]�kL�%{��%��U��B�G�y4��'u�C�FIB���tȳ(���
�NA�n$Y�O:y��3Z{x�q�>�QE{�R-;3��Hj=	���1�A�Qp��?���t:Ub�(5`K�� �T����U��<���m}<���Q
���ds��X���^Լ������"���,�V)�J/~M^/$R�[��Q<��#���RI�/}QC�!��
>e�M?�D�����ZC��"�͡��ۚ�	�dG3��5 =�-�- %�`�k�yW$|��{FYA�+7F�xƈ�}~.���,���lM���ʈ�}J��-���!��Td���EX�׸��q �Q��Q��r#�'��i҂^7����L@���W�F��(���NK�k(����W��:��-�)��|t��t����[?�T�.=.`~����J
�էjJ��!U��蜘i�D��D�[{`��"����EԶ[TFG�"���8�)Y5c/c9���ܟw��\�Ee𤏦�|�-&ʮ�sn�e����S;��R�f��	B�#:�e���`�F�BI�칕�!!s���d�9�a����ojX��w�|@���T����y�-�HU��4�e��&f2H8D%��=�����輔q��8��r\<��? �r�1i�LNB`]����i�<�-�wAW*F�6�l
��ʗ�`�P�+>G�M<	����uB��C@�u�
�����$��'�w%7�p3s�>���	��� ^�����@���r�p��;����0@U��H&[Q$�#p�� �E%�������
���Q����V^�q�h_b�wc����̱~�lPTSdltM�`mk��T?,�LA�m�"��g�\�%��M�RP���h�O�N���8|a��'� ��[�PyƑ�̈́�mq)���|f��s�ʨ�I��[��8��V�N��0�����{���WNmՆ�l'����b{fu�雇�S�x��H��<I�l�Wa*���B�,SfݛOB��]���MDPM��U�ӱy&J�~b��_j�󄣆�o�� �$����9wL�q�*�fB�%�㉎�Sg�m7P��ҹ��gA-�͟���d,����ߟ�/����uo�烤E��aU��~X�?�.�'��Wγ/��V�2�x�����)��Qf�_Bqc�WWN�@$������.$��7��4+d�i�Ki�v��i��^_���Yf���DGJ�7���O_bq�0��:)��"I�/?8��Ҋ�A��$w37���t�v��9fOF�h���u�l֖�8�On9aJ��'�zA����#��*ζ߫i[>h�'�K�+�V�(3$�e�f���ֺaR<��.��R٣�%��ep3���a���=�Ï��4��WϺ�a�2�h�G�'�v`�0��*���P��(�4���GIȈ���!��/�/��)�s�I(��s���<�x�[���W�V^��$���
-�U؈��w�ā*NM�f��Z���L���M	�8)�YPZ�?"P�lY�3�jw�i;�'����}|�
�[�W^�(=��Wj[�_�-8�I�DK��Y�9A�m��8nf�D������4�G��&kf,\�6���N�bb���;&�/~�."@$��7��_9��p�JI��uh%S��3c�n�A�|x7G���Uu�}@��D�q�"ʅ#^��/u�H���v���Z-��vB�Zm��'צ*7!�}�-F%:���jy�c_*=��f��{�r1��S��u`�ĺ#L�ϻ6M R��H[)�t��Sk|ԧ0�~�k������{6(� 1�>�
�W	:�M/^��at�U5�]�g��*�4�`8������naos m����8�)�|��[�g�T�{��$��� ���ߕog�K"ZI�ێ�*7$ap�L�ߍ�'}	SbͧKѦx�([#���uWɥ�|��jш��l����$n8��t*@�29�W���U��P�s氖�)�'=ȩ�P���[,�$��KIl~�;���=N����"���&��������%�6�M��cq4*�J���T�\M.4*�V����%=(v�s�����O�#�������N�A��]�a�l#++��U8����K�t?�m�f�f��7���a��h��<��6I2̔�3$%����b���E�t�,S�m�p�]R��#�,�,�֥ήMaL�����~%^e7�HEvwy��н�t`�Ll��̈��[�>Y�>� ���ϡ�yd��1dm���Ei���z�sH�&�5�Y���$��^48�<��*(b���]m�7KY�(ZD���X�������a[����	��o�AP�u�����q���!�V#���1���*Wh0\�9��'���di�����2����f}��#�k�]D�.�����{���
�[{j{ep,����Ko ��>��f��8�KA_��tkV�+�f�Tܫ����>d0pA�*b��\�x���[F���Nc˘�2�1�~�6�����]��n��6:�7�fG�"{�f#���$�StL��Y椅W ��B"�Y��%Gv��L��-�f��M���K��"}��7{��U�Aӣ�1�8��W��f�����X���E�:iѬ�8.Q��h���6�zD��K,���3�RG�"�k��E�W��ř��	�|�>{&d0o;o���!��bU>����tO�}��F�q�����\2lP�A��_#��F��ɪ�Ƚ��+do$Qr�ȶ!d�gR֓�$&n�u�����/\�b�>�Р�n�u���^z�����P#Q�P�)6n��3�ǙFuD���ޔO~.� �H�h_K��d\NJ�t8��ǆ�L:7�ו=Io�~@�iQ�Ǒx�r���J(�p�X��4����	��[r6/Q�IT]�l���7o�������Tȩfx�tև��):�V�=�9��������}��7S�b]� ��G���7�z"�b�t�����<`�@��sU�$J��Z0��%S-��'gm�[�-:%�M���J�!�V��W�9���SI��������W:��I��sY�&�V�,(e�n|]#i^C�N�89�U��g7��S��ȷ�o��ɬ�/�3�T/�N��lrhP9*��o�m5xW�.+I�����"O�����K)�f ��:������̙ܠa� /�V�W�3��1��½���dW��;٬�׹_6�.`d;��,�_�����A��!��!����$��5Eo������TN2�ɵ����?ם�ϙk��3��F[1�t�����6ɰ����q����sf�f��3$b��S�ə{;�r,�
�4�dVȶ�#��q��b]�9�MN�M�t�K�?՜M����6�4־�E*4���t�ޢ���^o&#�A��&�Ѹz֦�u$�Em�rT��t��۶J�8<��APv0�͛�n��9��
�ٿ���� �����u��m�7>��v�(��������R��`ҽ2g��-�4�֬���_�ٹ���W$y�S�����pVvt^��d�C3s��s��i��� ��qԡ�*-�Ri����i݃�"O<lګ��
�X�Cb�c:��7� �z��Xb��~'[���4Ӣ1
�X�8LY�z��rl��a��I�Hc��;���k�0��;�Yn�,-�S���	`ћö�R\xX�T���������ϠCpk���s��S�����'�T��x�i�vv0��'뻧(fq�9)�s�pЃ�ˤ^�����t��Zts8�uGF�Z^��n��V�JI��
d��������_��pq����,��(]��5��nzد�������$��@h�����KRA{�}9\x�K���F�
5���	�i�8 5����ȩ8�<����R����O϶=���T��G�~W��-��y�PO�Ŀ�|��zi������h�S,���\4�u�(ߥ��ƅ!f��L,	��\�mA!m#MW�[��+;�I'�F�6u|
V匈+tˡ�ہc�X�qN`#�N��M���&Ѳ��c���}
[����w��gn������.��:߃d�X�!����!T�����G�F�������w��w* ʽ��+��d�مnQj�6k�u͢;�g���@Ӂ"�s�Ē�Z/5�����T������s�3M�^,���p�<7��Q�����/č�*8�0qⶵ^��#F�S&�T���&�9�T�Ѓ��iV�:����n.��%g��@(ݦ��J��_����UĽA��͵8�o^Ρ��a�۟�� B�nc��gi0O�����HA�C߿��Ԏ��
���o2�N��각~���5�:t��5�H�,���@�0L�£-���Üʻ8�Dݔ�0}�؝�B�������H�U*~��]�.�h���? 8C�%�ЫE!~!Y@�K��i�@
����]��I9��y�FH`w�(ʒ�����m;��'׷s>
E�@X��&��%?>}�Oc�i���¿uI1�ƗA����n��t�Q'S���cE�!�������x�x��
Vo�X	�>s��bO6EJ�'�{>ڣ�>���GU�Ƈ�hc�'�ޏBI𛓃���q�M  �v҆Oȍ��e��&H%M�e��N���18�낻Py�	�c�a���Z8�^��Ym�ej�y���i���zJ��K����^J��zsۻ���^/-��]G6yL�B�s��ɫ�d��'�l�TۑP谂QٙUd��� ��>��Ry���<jf�9�����C�Gw�0���A��b�P���U�?�5�Yx��Eܯ���wN��]�E�삨T�u��ެb�nu�>u5w��{CM.%���hM�A篋݀،o��"8���v=�7i�>`��"d�%��c�Oԉd0�Q}�+M�QN�0�.*��"?��=��������ª�����G??��+S�׍h�{�כ'M�hc3�4r�/e�kH�f���_!�!yNS��1g�ݸ�:69䀰24m��>�X|����c2'���W� �Ơ8]8~�0�x�Bc�"��l��J�~�c�$U��v�Q����ȁۥ��P(@�"���ݑ��J*kRb��+%���ޟF޾k���*3%��]�6����3���̥�>W&U���}"�5�J��jS�m��>4�����[�̓����q-�ʍ�g�`\7+%���:k6��K������-�����n��Q�q�'a���G��D[�<yNA��"p5I� ��ҡq�X2���Y@�z��ͯ��~ġ�$9�`����- c7�����=1��Ә��
q��R̘�^���zO���q��̶�ۈ��ѻ��|��KE��1�>kv�*q�*71<��:���� �~��kT�5�@�#����ҡ8٢����K����]�:R	���I��Um.j��~`��g2�FfɌռ �A[Ԛ���,5dzs�/��~��� �e�c&��ÂԱۚz�x�t=ԥc)���W�]���2�A2����Yj��r_�"��X��u/�����+�H�8���W��K��S�IM����?H�u|���\�4ڥ�/I����nIEK�k_� �AP��V֗�.LuU!��G8'�)�cJh�,��bW�G=�ĉ2n|o��w3ͦ*��/)R]Y�U$oD$�Pg@5h) -SQǳ�����Ô����[ƨ�0d�Om�P����_ȑ�~(+ف�p�5�i���ӕo��|���i��2=�B�Y��"θ��$\���I��љ!�Z�46�%>ˣE]�ʤs���@�|��ed���/0��%Y�E�Az>�}mI���ytu�����!���R)���o�څ���w��<��0sXV!4�E�VT�7�M~�h����u���l�a�F�߷��s�$�����*.�^e�|�y����H�o��)h�+��`>��/�E;�Y�{ �{Mxx��:Th�7�<ˍHș2��Q�$V0�8�懸]��W�E�Uծ �Q��S3gft�-$�9��TJ��mw�og�?�c$d!=]�����:�wA�}�&n�����h����ѣڥ�m�6P���
��7]�⠹)�Seo�4�RhU�[c�T����������8���I�X�1iN7B�ݦ��Xn�֨����2yǍ�@�ǥA8*�~����޷7G��4z��rb�K;�4�-SM��-����#��Y6.?Z���D5L׀�f,O�}Pv`������S�C���������ت��2���.x���Gc ��+dI���S��֎����Q�n-�p�1Ң���v������,��hv�����LW(:v<��\��fql�,߄'����~gL��4k.�:� z��l���Y�ӏvGy���}��<�=|���|ɜU������Gx� Z�{�U�,�u:��",���րԷ�p�i�^��X�N$�wcj�0^�dr4�0-�ƪY�:&>(��q��2!��c-H�~G׻�3fU^�3��~�{��9|�+sj�)�PJ`�J�IK5260) �S��}
�@ۭ,v
��ts?��<3�O���M�S��7����^��M����@u�/�9s���%�+�[p��9��x �p���s��P@X	U��q�q�����H�|�{?���� [P��d��;|RZ������5�Wu{G9֠<��%F���h����܇Ds��2��8(�mz;����>*��H�=fR	F��)����ɗ�̬[+���5N?CK��5���3L]l.�6ޖ��`̶+���,�Q�Хգ	����CG�L�宐ܻdL���8iѯ������Z!��'2'��+�9���8m�L�yj#h��ڢ���ɣy!ʫ�:�K>^�:AS('���r��dpm�k��
����trx�mW�Ð���v�`̎6 q��:*_3���-ۘ=�K�&17�x�?ee���3��2��T�<(4}֓�I�?O��^��٨}b����bb� �^:������pT��u��캢��/�7��\�=˰�Ҡn>���m�Bj���17 l�����a��nT y;�1"[��Ꮼrܛ,��<u�ZK���I1վ�'���EL5z��t1lZ�,�20�93238��3sݿƥ�� 6c� ),"�1�|j��!;f��!bW�v���{�A �"Pi��,�s���\�����D���a�7.\�yR�`媝��{����x������t���H�p��������������5��߿��eS������&����ܤ0Y�-s�FR���&26q�rĬbw�9fe�+�j�[G���=�i���'��ND6�Y#���}O�H�]؏$mJq����:=�7 Cׄ��;�N�@��mS>��P�8�8J#����vFmĤo*KA���%���F��-k�9Zc.9Pu%�z�q�ri�mV�6�Me���D/�=b?&*�/����
+ s��g�0�EPC_'�et(�qC4�|+d�´�/�C]���n�p��B����h��?�~#���)���4�+(��⪚	9����q¶����K�5 J��-���Z����^{=��CS ����h ��O��=�3��J�"�3�{!�6����3����{`�#1o��$�N���Ck��HP���N݌��ϛ�_�>�kÂ�h�!u�@K?D��	�mX�@ɦ����[+��2- 
�ꗳ!&Ch\���[��ˊE�JH�=E�Id�g9��NF�-m�&y7V��n�����������[�=��nZ/�ϴ�B��C`h=�.&��1��fy�_��:FI���T�R|���$�M�#ħ�����E��������+��[�avFaّ��)a�2�1����ګA_H�#�W�X2b�б_ؐbP�Ep��dJ+���f�H V����)~�lh�]�s���Eq��H:��,�a�|}�j���td����T.�)
ؓ�M��l��jY�M�oMz>��}�������"Nv��M]�@��nT��ɰc������H���."{%+�'0N�����PC�I��g��i�*�|]T����,���L��7��L%'_O 8s}��1M9��&i��MY��q�J�bV��y��'$0���?pC gUP�c;�Q_��dg�K_V���t�	F�X7=0�cFJ_�| K��DY)_in5�:���F�-��H?�s㷽�@��Z��N�i(lS(�C��7`�� ^�?"�����P.-��������cX4ճ=<�d� V��xU���1~���(��~������E_4���I3İD!V$���w���t��X�G�<�E� �p�Ӣe�l(Q#P��D���y9j�T�:7![��)�g����l���N����L�m��F���'t]�����t+�T��Wx5�y��k?�Y�Q�s��������.��L��������S���z��Y\ �﫪�¢� �t\��9�6-�xv��$�v��zkL�h��'����Y!�ء�^�h �3w"��erf�S:e�T���fȯM(��q��oqB���f�Ty��$�3�S�u�W�)�Y�-���a�(2*ʝ!i�)V�8/ղF���T��>��`�|L�v�c�Q�[�8+��X���������MCi-\�;? ��x8�����A�0Z���ȝZ����-�H�
��U�}�ge��!��h����S�\<�g��K�o�{��`2ŕR��Gj\��}%_l��t�5g���r��x��خ��K�K^ov)�������h*�hk�b�n�<w�,&*D���.�Q��� ��q������j&MZ�@��`�������t�"��2N��8'(���Dr%�^��DR��YB��|q��D���*Q�څ:Fm?�<��$�N�|#��f�l�`���:������kY����'�`�clAS�V7Q���q�k�X�q�'qcre9�4�.	�0i�����vM}4v�dr����yX���{</�"���?�ðu��]
�rc	��&c$�v�����F"ȗ0��u�B X ���}U�l��Co��Qɰ�C�R>���O4�wɱ��WъuN�ϻ\%���H�����w���R�����ub�h��u�����?re����`>0�#����c�kl��$�n���c�W�b�aB�Y#R�NZ`�L�&wQa1%$ߢN�4���姏w��	oΔ!��+ZZ��#��%�O[,�o?�gKv 1'�<(bЅҤ�]q��X�y{�ֺ\��{�6JB�2�g����|p6�C�Kћ��
7%�Aư�Ѱ�N[䯏y�+k4&��U�חՐ�7O� 4�d�q_E2��~��q��K8�z�<�a8wq����.�z��OZ��I��FĄS����� �uG�!�td�0ܝ��bsN�� �.�^����>[7:U�m,���A�
JaS+��g�'w��t�}8�K�={��ڳkь��sUj��c?��>� �I�g�w���1�{�	;ʔ�~�
d�5o�U��`!�ι h�9������x�[)����o�H�`Fg8@�S�I^�Hy:���aSB:��6�>h�#� y��2���G����ҥ���<f7��}�cZ7����� �t���]%����.
�P�&A��;��_�e1ְ�a�8D#���H�4���$W8'ʢ�ZU�K�H�u\�:N���I����>
�"�^U���8`(h�w}��-}� ��Ϩ����2�;�P@E��%�vG�����}]�X�#��nQ�2�Q	SI���k'�̶���\��f��v����H�o=|�7o|�^�4�������
LL�,�݂�K)3���B��9c���L�uY���)���Rq8pI0 N�t6�j�0��|�%�a�s�O�i!K��V����+?�m������39��$�����%�Fp
��~{�i��Z>��b+��5�cB�8��>/���a�'n��!B��_z��ő;��S���-A!�8m"�a-��=j!�\_���p(�^��p����s b̜S{P�E���.4�͐,�؊��6���͉ˋt<�����K����i,m�m�E7�Ju	N�G`�����\��#��t�$���D�_��XB���S�P9�M�I�����i
�ׄ}����S��Dx|+"�~��N��� v$n����/�)}슐ER�F+�٫� [��YeX�H�E@;#�ߙ�v�-�_T�S��B�I����(#+� K��$N�`"�mX��9?V��<K\��E7 %6�����Ҏ����Sx���jZ��EL,��}}�i�q^��C�3��F�maN�^癑�����l�.�Pq�9n�_ۑ+B��HN[x��h��s�:�82!�����E�;	&��x9 �3����Db)q���fIH�ꋖo�Y�����������r�HK��@�p-��Z9�ֽ�8k�8��b_/��y ��� 9Q>a��ٹ6#�d�-@��H����c���.�0��=d��Pj=�2|���{�����]�]*)�n&���L�C�z��G~k�Ӧ���DX��n�8_�d�����%'�޵��C�,�K��r�$�y���k蛟�ǰD1ß�lWQ�k�Zt���0��آ<8�6X�T�P��s ��Gjҟec�}=�Ci;�

F���5HE�$��3���g�� �ly�kjq4b?m`��b5�@k��p|���:��;-Z�Oa�y��Ii"�z}Ws�U�a�"�x�c8��e�9�8�}�u��y��a���8�g�.uo.^6��H��Q��D��N�,�o�a}�7c�V�Yc��ˤ�K������oX���JV$����ɺ�v�u �mZ:�a�jz�0dZ���(����xk�2 "i]\�*�b���A&m�:W>��R`#i'�c�d�^��@�	�9�LŇ�wö��M�ϯ����V�v�����>5��Y�Lm��2��wE��AL�:��J��	Jފh� ,7����^K��y)="MSd�
�s��:�[EaO���jospS|F>� aar0���𱴁�T�k�7G�ܖ�#�^g%B��U�B���?�hÝ��I+o@{���s_�s9`��,+f0B�OÛ��@�,�(-�~�F����� �F�Z�dG�x�C�jolL	��)$�7d,z����-э*��3_�+(pe�w$���#5�]����0B>��]�B�����s���������e���=U(ݙ{��~��w��&<�>m���>�\���:�=����� �H���@�lۏ��~��՝�q"��NMa�^j
�� >dq�P�;^$���a8��siT��a�Ҋ����
O�K9��D2�����ڐ\�����l���[����������Z"��`�~Nyy���F�v\Ɓ
&�
�F�3v��SI��?��+9�;�P�ҿa�|��p�6��'� �WX�xu{�{j^ūŏ=hO�T��zI���wf��W(m���^m����}��ҽ�^��-���� ����.��%Ɵ݁D�~α���q�Έ�E٪�gl�N��P��IK�Qt]^ʴz@��y��p�Z��h��Z؊u�R7�M�	���#�$�?sRd1��	с�C�Av�h�q�_F�v��R�ҧ۶zL3�E�|�Y@.�F{@΀���w��0z��jӡ��j��=���[�����Q�I�6{_��u��n *&j��
J�d��^����w�d�j�1�E����}�U�]4E�/�u���#��t�����ւ$�0��6 ���H�n�Uʕ�޾�p�Sd�'aG^�9
�4U�������|�ق�6'����eB~C��?c�җ�[ip~�_0L$h��6t����6����9I��mǀ�L>��ly�~�ܽ�x��(l��cH���A����QZ�E���BU�M8��k��O��?�<��su��o������;ṿ3� �P g����klt�����L�u�6
�ۓ(�.��&�P|Q~ �7�q?vMP0�[o��)v���G_�9ƭ0W+N������9[�G��\`*R�z����,�"5��#?c�g���L�S���D���9�W~ܣnOБ2R�J�<w�I�,�Ծ��8��hOE���ps�N�x��I�G)5>�ҝ�N��W����	����vϲ��b�����^��~q%7�[8�
*�tSI9z.�k�������p��R;��I!�p��>j�娢/���Ɖ��lLH!nV)Ԧ�n<4��R�R�������0CR\=KP6���)"�y[he�����Cב._�<֬,�~�s�Ibj�ӵm�az�]f����SX�i���@r�g�M����̳�$(��0M2�N�l���*0�U���(#7'p-�^���iڔ��<N�u��8h��E���Qz�NY��/7a=�e�Qր�H���bV� hސ$��tK��%�x߄4Q5OO�.�.M3k�$����7���:(ŉ�Rwۏ���:��YW���)��#T�*�9�Z��K7$5m���Y�Nk�HL#dC�q� �8�9aǺ~<݉�Q>�e�������<
 ���QKsf�IV��^��^>�Fï����\�bz��S/�}4'0
��{��R��z?U@Ą�zf�̒�ʓ��H26���m�A1:DU�>����=E��U�����WFW͊E`�W]�	\����IAߖf$S`�("h��*~u��b4��M#z���:���WI�
�sHD��"����j�G���XvoB�d�8Ef�x�?��-��
�폆h��HRD�����d"}�NV�֙\~�K���q�5i֮>�����v|`��n��;a�D�A�<�k�ϻ��-�wɚ�t��
�2�8��=��u�5�Uc��Z{co䀟Cc+�߈�A�)�{9YCm�pL�*�M	��&3%���ut%��
˚�>٬4[�M�;�8��kd�΋}A�����@{���m���UH�GT95UG�Qr٤#�N ?(q,5��(tRQqo\��H�
��@)kǈn#�$T�ha;�XVJC'�@��`'�9�~�&z�IO3�>tT�g���8>�I������e;@���ε��L��j���(��~�s�uDړD��n�z^�@e[��0����j	�t��i�7���i�6/���]6�?������$� \��<Ϟh�UߺU�������8O������V٧����}<���2S�8����T��pp�0�6ɢ�����&D�K7)q(/��/T�SH�q�٠YZ���c�� �;�=�'wpY%��t
k|Vm�{/��1��/�H�ټ����B��8Ӫ^����.9�ky���nT5�zA�A���E��ɟ)E̎`0��7���i��LPh_��3UiF+�2���%-:��n�/٘��1�҅��1b�hB�[���D���2%�><�[#oE�e9qj)��fw���`�����U*�\99}X�0���$|��u����:��N���o�k�x�r�����3+���(2R#�� .��g{g�[=������N���_�	P��ٕp������zsc��!�^�{�$gu��M욚�����>"�����e��4�?�i6̴-�uO+�q4#c�KV"�]�i
��ɸ�l0Jq��pn7��/&�9�.�/{���T���t�R��{����� �
�!�(M�"��4���|cDO�]�q�� �7�T��_�|�}B�zh�;�&}S_�=	ݠ�o�`<�d
N��A&�����?r��pu�O�}��OV�_��؟B��T'�(����~���c4/�i?|�n��(l�	�p��t|��(#i��eʫM���?5vXW���V;����Ӛ��n��n�q���Y+�z��!6���dWsr4��IČ��'�e��Z�w���T�XQ�^
4�$���l�A$�f.�o�7E▵$����^��v�HHl���v�?QuX8��0�@qUk:�f슎��Oh1��6R�^]���iۮ�GH_J����?���!D4��ė�����.�H|�JKΝ'~L4����׺)��fhD��¾���<��/�~�8�1Z�9Jq��b���p�G�HgC�$�c �����CZ�cƕ_��^������ԥ�Yz��9fH]7�����A����� �����B�@<k�VHf���!��>Stv!s^멍���_�fӨ w%���� ���D2 ��p���}V��U��v����y�P풯���
�`K�@H���T�ڞ�����G)������@�a2?��c�˘d�@�q������«�/�D�p�"����u�����M۠ڈ;;������X�l�M;����X0�<���%jz*&t+n����q�%3�:m��[��נsLl��3E����>eu�X�dm��`��ԭ}�z�g:��:����d3r�'�P�49"�Wnz�=�?USJ	J���~�`�aw�T&�$#��8��?��zg^�uJ2���9`dv������s�# ��6q��qq� �j�V���ITu��7}�]�
��&A�P���f ��d@�x��}|WD�T�A�θ�s�E'����B[�W?��6�
�����O�xiddA�&�݈��I�=+�ː�0d�����PS9�(�1�~c���ܤ�g࿢ګ��H��_��qR͇����j��(�k5����2��}m�e��=��A��g���W�e&��r�iےSͷĵ�3�����ߓ��c��
�>^��q�����d��a�,9�?��)xx�s�� ��"4�h*��x�炦��U���r�R�=G#�6~��<��b��ԤK��$CB|��q�
s���ެ�˪H�>�j�-�݆�i2�STm~�-�[|�d˨1:Ԝ�IN[\H/)N�e3cf,@,���M�F:�FW8�81���"�d�����Ҏ{zQg��EO�a�a����Xxg�{3�Hd���lL`FZ���;݉v�+[�9�z+�*�?>외�Fl0�1�n-�1#NY�a��_���_<�S��9�hs'�+
%/o:��h2�dօ���Z7Y7�!��!7ie��)�'��ļ��ju��z���,b~B�7��J,r���</kF� �F��j�s6xwa��1�`qLc[�Vjψ̦�Ѷ�=)g��!'W3M�|��g�s�竢Z�v�%�Gl�}E���ջ�`���Ʈ��Mx	�@^g����g�9���6/�$���ȴw�f�N�2�D-3�]S5¥VDĆ�~c!���4�����J�,]��F� �-KC���ߍHYW-�N�?K;��蝼b�,��N�:@b�e��J�H7�^mZ����	��g�����!�(��9�tB	^\|��e�+.�\Q����9�^}�%v�lG:��&N">�,y��4]��	�����})H$7�vٝ	�k`i�4�H�a��P��4T�
#���k�%s˕��Qjh����訠
�E�@-���6n����,Hd�Uīc4���a@%���M��G,?�s�ʁ`-�쑶	��9�b�4���sޮ�kj�0A�5�7�ΦQ��+ٕ�����D>�����ǆ!Ք$g��|��"��>)��+?�9�y��T�Hj��cNj�d���u- ���5�S�t;��U�U^	&�vSxTUT��6�r�-���G�A���8�QQq!۟^���:4����KV�����e��K���G�'`��Ta@���6�]L]�G��H��۹*���QI�t�Dyk�յ�&�􂺚�/,�+ :��̺�$�<t��	����E�*�f�J�d�9�fhtLEW�m�EVU��"ˤ����Olu�F[_�K|� 4�Rbf�9!	f!(�L#��[fL�+[��t	D.n� ��u��N���LY���ﻧ��L�j���g"c�Mo�yؼR	C5�Ǭi~;#w
�B{��`[���D,0���I8����	�E��x����o�y:�l�7N��}e;98���\� �ڍh��L�ȰBTA���!j�j�ɕr��S��ea;��+��5n�q����Sj�t��Ǧҏ���6�I'�A�'�*0R
�k�#�
=XD�5%¸��ul��.ϰ0%�F����.��~��\[��6�R��m8	G)\H�%q�1��u����7"�c�Y��G�Q����F�������Q��Ԛ�0�DW���T?���5��ZJ46�I�ϳ��-�kiK�l��?��+L;p���h����?S�{+�%�h�<Q����Q ۆ����ּ�~5��S�k�í��~���Aj����9N�������z��N�8���_x�g�7��#�D��R�7cf�h�Gxkqr�D����'n���`�P�"*�jM�ݠ��v��=�`9K�Dȧ�s�N�� b�t�����@Q�'kvauwW)#�~y��ӵ�s3�8�[*.�b�.P��m���Mf�E��e��e��d�WD�J�g鐯Q�-�UaeӋ���
�$Z�4�5�l(������Ҡ<��ѵ�Á�Cݬx&+q�r1�T�l�<ꃱ�Њ��c�/rP���F���>bN�&�Jg��I�63�M�!<W�
�	�%dK����H�3��FC+�fk����1�&�n[O<�h�ىQX�3�ѻ_���C�ܜQy����U�b&6ƨ�am՚�U�%�p?����nȎ��
(�ˀ	�������^����{�����c�|��/`�la�9�+��� ��A�{����&D����������.]��Hb���i���D~�8н�D��n$T�-g��f�����2'1w�:�.30����Ab��Q���i��	d�:B�}@y��^�hq��ݩ������ri������>,�8�[F<oG�)���_�M��f���LQ�0{�oh�r�,]P�	���^�KJY�؜�?1�a�t3��@^�#��k�t�iG:8y]厀)cW���&s7���e)��#�ASC��ۛ!�� '���P+T��N�M�MO��s���%SW&�X��В�i�<�����0��W1�6���j 䪕
��x����e�M
��Ӥ����Kiـ�X_�B��`�r=����ހs>��u��ռ��h��WF��,�o���:�+��!��O#����D�؟Q6C�3�bt�� ^���E�����c�]4�3��7ql3���d�gc��P0����E+ɻ�OH�v�T�����H�c�P @�;	����/�@����A&GQ��cwU)!�1D%a9�0��/�sL����jj�����:��N˭��mq9�vܩ{2�V�0�)�!a��*�D�-dr�
��%yxXB�n`=|��JD����3�an�q����/k�5<_/�&ByO[�� V֟S0�ot�����k�����z^���&�ͼ����Gޙ���q��:2��n��B++=��Q&ƪK�� �43	�'������ �@L0��	����Rj��Ẅ�s�ih� �5�m\��i�t��O�~�p�6�]`��GQ؍վ^I��H�7����(�����v� !(�9Ǝ�� ��z��Q�,D�>���)�'���|kO��+pP�|fA� l ��
�x��8�>�"y"�nH2⎰�Ǜ��i8�z)Tځ��3�u�ȴ
k�Dzw�U6��G�W���ߟ��JQt���к��
�`9���>Z�$g���