��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|n�\&���&��:�lQy��x9�5�A6�Nv;}PiM�V���;�4�ݖ��`PrڙD��� :�Z��O��^Cw�c5c����x1����T�d��5�u�n�3QҕF�s�s�9��=��N�<�{�t���^D��<���`c�s�tg��(H���n��og�U�k',���\���Ao�|�d¼@T��6G-��L*`#�о��B���Ah�
ZpI�)��B�=�Т��`ɠ�l4��Gl�V�֎��v���'5/��e����Pi�!k_�g���s�f>å�1��e�����BRq�؂	0τ�d��	��7[m�#8j�>[�9A У�d�)R��+��r�a
]���;%͔
��Mج�n�������xk��\�с)	$h��u�E[��7�$uT���)��vߦ���2Λ���d��,�w[,Y &���D�
�X;���B.����BV���P�,k��'Ӄ��T���Z&Y��H���}��_B� ��2|0���O���^_ѩ��/4�ė��'I�HՂ"z
��d�V���e�=�f��U�^�.d[U�&V�N��xK��\���Νǫs�e�rK8������I�G�w���/���<vU�"�G���l�p��O�BX`�IB�	QRD0W��q_Y��1m&��Мc���C�#6�-�L��Y�"�X<�)��y��V�S�1��M{c��:�|��f��X�����	͇���~	`t��	�jz��p�u�;�
#�ҟ����������7��O�%�������_1��,�����\���8���E򸧶=p�M%�ʸ��Bd�8XGM�*����> ���Wcv�klwI$M���� <z֏O���X����	@@.\h���1������BT�#�?1$���P�>�$����	�e��?L�(>
�*��{}%�` ��K:%F1,·��	�7]0���'T���8J1V�a�!�kK��E�'ȁ��G�]�G+Cm�?��U�/��f� ��*s	�[=����=������s���+���[)���Z��3K&9�0U; �oH t�N�0V��J�@p05�/R�[��&��;�*o��)z�G�ZH=W���lb��`���Qʉs�T����İT=dV����_J���-y6��x�T�^S�u�^���-�2�hO�=�$]Q1���hc��^8��x���$�9�W�� A�S���|�,��5�A	y�;eo���%a}��O�I�s���H����Cj53���N� �#	%0� �DZ�4�	�'�!O�j @�0"��G3���RA�C �B>�(��^3Na����$�2?�SӮg����"V��wj�h�m��<ᓄ����AJM,�[=�u��1yȹ�|Jr�Z�������QO	fɌI%�a�C^�Qj��b��[�	�l����{��J8P�{�邳��oИ�؀��n[��']�_I53B�j����y�$G�M�=�~�l��e7�ɿT�S����6��D����h�B;��4_6X���{���
$t�ƹJ��l�Q�Y>K)=ߤaK����;0gp�Y�.�:��tY���h����I[@X��|+u� l�[�)�ڑ:E"è�,�9�7�d���H�D��6����!��:PZ�M8��eP����d��뉣yui�h��kpsV,#���"��=��U/6ꌭ�%&�2�$�����P�t�U7F�Ή�d:��[�'N_�!��<�\TwF�a#sV���/�(�cح���u"���'q���lD�'��Xow�at��)��mN9&������jE�H��P� �	r#���C�3�*�Q}�1���Y$�d�����\9ߥ?2�<���:ȥ2|�+�[ӼR�=Fڙ�}>��o�r���3_�xh� ��p��h����:�6�Ի��J'���)Q�ƢnoZ����� -�B!�w��4��SzO�	'�7���Y���e�pRם�WY�K����X�!�|W�1��3�u�)�A"wҨ��X!}��6*�:݊J��/�VH�`��q[֗���0���\D}^?tyL�#���-?����ǫ~^�N�V��M>3*����9B*fK�U;� x���	6@p�9��t�}�����[�ΐ*�D_N�\ <U� Pв��� ������n��#Ci����Y�c)��b�{T����A�Ċ���AwT�Xo+���6���t����8E�Ŏ��JXO����9�kZY�æ���L�"d��NAW4�4ŭ3W�r[
��s!��n�f��t�?8���
��^F��m�Ma�d�]7[_�8q��1V�R������-�j*�L&R����	�ȕ�L��y#i���"��GM�X�H�F��Qt�~8�[]!�?'�����x�&D���`��Qd��=�9#KP�Y՜��W+Tf��J�)(A[�	3y{ }K2~���<�IC7�ò���S�w }���4	�
�}�0�΅��&`҄^H5㤾��&�a�9�� a��#�1o��CSa�9��:GA�¥���
 �+8Ҧn[A�]���*�
|&g�8��8���k\��O�RQ���~�XXQ������T�c�Β%�AfT���ڶ��:0�H'�5O�3��@PT�,��b8Cl9:b&���4/��(y�j����u��7AW"K����*��)az�v�L�q8ԅi�p^K&Mɍ	&����{2m�;x�4Pw5����z�g��~j��Ż{��uUB���VhoQ��jVY��%P�^�h�:�&���+aݷ�(C� ���8�7b�� ���k���s����n�s'kM��~���D$Q�B��PJX���f�a"*��CKQ���ڑW.i	�U �1��j��C7b�FiXqgkm}�$V�M���&���E��o�����{Er��)�%���҈oK�DH�=ǹ�Vj��K��oP��b���� Q�Hn�9�]�D�m$�������_m٠��̈́;i��]�7�*�$g�}�7[g��׿���M�h���I�IFg����"���/�>�|�bv��f���|z�|�Z��2{�f͸�08*_n����x�v6�Ք1��t��8�(5v,�T�����4�9�8�؂��hh3�bX8Mk�K��h޿��q+�݉-��^UP� ��D��OW'���v{��4�����i�,u�hcb)ޡg8 B��������n�h�:r֝�t�����LCi�C)2��;��� �;�CN�wO&��&LD�aayaᗋ�%��T23.�l���q��M/��A�q��5kI.w�AKv���#�(��EV���B|���Y���nZr^bW��<�lP_�G"v�l�Z�)F���;��k/��l=��jS%&�rid��n�ty�S	�GD%��_(|֕1~�uz���՜t��<�:�� Tb�?-��*v�7f�Y� �f SyYS�� �U~+3��Q�^}�X^]�$NJ�&o���15Q��mܰGUTH2 :�E�,�������
i��Dya6���5�	4�&�/~���)̹9<��Y39Hp�yGH��J�Z7�@7�M��������[���6���M��C�&���L�f�/c�}���z�Rb��@@Ө��e�#��+��IzJ-gJ��e� ���An͔��$w�j��T������KÚffC��+z��9B2��l���3�4�}��B�S�ߎC7�����2�y��B���T.�.,q��>S,S�rӻ�/4�OT�chS�4a�U��gO:cW���k!��t"��H��Y���i;��3���\9��
�(��ă���E��W�=T��Xx0�qK3?��Hs�ýi�%��]��"�i
@�-[n�)�_��+yU?�_�<1V��~\��s�t�bI]+���V��?�J-n=���/�Z�0��98\�!��"Q�(��B�T+�M�ْU���xЂ�I_?e�KB���Ȣ�x���� ����ݷ�ȱ!�~f�����|��EL�Y���%Zx�u�?,�kaFcF"�[C{��$�3A������U�v� ��-;-�پ7����Z?��p�
�Y�3+��>�i�:��/��@�%��,a�vk�k���Q8HȟA	P7C"�M;��[��T�+����XpW�Hq��4���<k�w���8%�i~N�d�,4Ȉ�I�s���<�m��`�S�O����&���v;��d��d+�4;@������Ai�mHӲx��꾌��ҁ�N�B�.�\��Iĳz�0�`r���֐�V>+I���)d&�u��)�!��r�����ƛ���+�0+]��1�e]o���$�Ԧ�cm����a��i[���;֎����b�a��
�9��{�i����4�;C%����}O��[��@D΅b &��E��D���f\�є���B3�^�3Z���J��/�z_����6;��-
��Lp3>0����I�I&����I�h��J�|��Qބ�qy��8�_?|�I�P��+U=
�}U������P�2���q�O�Ү/4�Hm�ߑ�dk�l�N��#	}��Jڷ�� ʑ?�GM7�d뼲�,� Aj�W�պC�뙭�P�آ�Í�Hl���i�r�e�t�p�M�n�*���s��\J4<�?q>�������N~"�յhí���u�0#����=��a���YT>01\�b��9nAosBpq薵ADpz���zS����\����]le/�1�I	fE�(�,���r.�<�b��!ʏq���#�|�G �طr�Bt�az+DJ{}'���-�D1�Y�yR�"���`B]=L���E*�3��V��H�U�ͩ1�r�����c��K�x��G���<L"��@o������k��7�5SMmǩ3�?9��(d+y��fU�a�us2�����xX%>9����j̗��<����f`��^����K������i�۴آ�.�~g���vm���c��8��"	��)#��œ��m0�ك^�a��g�Y�&5�E��wc7^/��u猙C�E���?	ZUB'�XQ��j]�a:���;}h~x��?�������V�N�����Ic����AQ�n�S���w8Sc�)~�aB
D|��5�Ol��Z���Y���bx��0��%uSR^�59J���?�J|�}���2���ؗ���u�a������$?{}�3Si���P�'�/�|��Қ�!�%A���\.V��s)�o�}��n G�̤�l��� a���Ҡ%�dT���*�_�wIT�:�M���Y �WK�R����	xZt=r�)��t[k����C��,��UI$���YU��`����"[K=��F&��}/<�Xx����n���j:�����'���:�ry8o��*;�p��٘^��f`0����?VuF�ï��:�T���5<'yC~�ާ�t�a��C��d�����ޒO7��ҩ�f&(��V��~�ML]L��������*I��إ��M����^c^���u���"�N� 
�A��Y-�Ĳ^������2����C˗��c��f��:����@é������6�\��]n���3�������k
e���jY�OU���h'�4q�:�A�P%$�R���ꪟQk��&<��ϫ-y�P'y�E#�q�4r�$����]"u�S X�@�s��|Ѥ������-��1�:�6J�b�{c.9
��-��m���a�ε4c�!����,k��yl:>��+��e�i�Ј8��o����c3D������=gG�D���ĲBg�37�Bo�&�v̻ݭq���}�G�0�Rv�U��� ҉�B��%IRT����K�qUI��Q��ǀHq�|�����Ȭft�.�qH�%�-���C��R���pjM��82����\���(�S/�X�˛��d��t�O�,�9jQ���%���&E~u ���ϝ�i�OU9����K#�t��\���R>C�S�G�`q<Iqn'~�#8{e���yD����F1/:<��ݸ��g��Ř���7��m�8'!~%�!�e��2�����_"F�F~Al�Jx.q�"�l�9�,����ݫ6�Y�!+�a�£�$Լ�����PP1 ��O��KR��ېE��p5��&��t�|K��y0��P�y��C,1�V�z;���%o�P`��,��LX���E�13fk�t�*��%u��a��Ԛ@TY �3A�z�Li�_Ӫ��{�%r�`��L}m!�_?���r���V�}�Q�S�SK�2'�e��9��l��h|@Q���d}�UD���Jll�YҲ�ߜ�^r�+{n��Ub�e��)�{al��~�A@'���e��z�A#�`�N�{l�A�R)�� ����J�t��t�L���o%C���U�#��(��V����4�UV��Ք!Ӭ���k�Yǵ{��k����)�u+۶�N(_[8���_2��T�d�E冫���"#M�u�.�w���?E���OG�O����/I�O�^>��9��3�0tLZ��7c;u�/<p\�D��4P8i��??�_2�r�k��؜lV�h��P�����4�obD����ۆJ�b�"�p#���	�Uѥ�/��kl�r���Ac�JM��-��V=�I����W �N�����'�s�� i�U�DZbk�(:���p��\�7�,����9�1��J2����"��5i8���Bؿ��C��w��J�G]�^�&�W�~��s�ΚіTr2��o���H0�Y�y=v��bm}��\��ߜ�x]�/Vf��i��4��jO�̽)��-^��+����ۀ�@(J���������=ؠ�l��,L�g���pN�VH�9��=j�'�`[}���{"����m�(
�Ҝ��[ ��� �L�WfL����#R��	�9�-�ffHz������Zv[уj�G��U�M��(��S��Mw��g���!�5w����9l�'U)�v�|��>~̘]^�������;�y�w��<���8� U�e�c�+�*R��tW2�"�W:�S_9�zLY�p$��Al����ϊq?���&�t��Qкg��`�TԵi֠���\�Gq�g�<�)����O�$��J�S6Ԫ�#�����+������9�m��&H���8����?�W�l8G*%B�ʋKf�h��Ė�Ҟ

ug����}�F�.g߀���ǁ�`M�wt�< 8���fG�l�)�FpE��h�B������x�Q�z'�f	=�轵�D��T��l�SS6lMA����M������EQ�F������:��'�����0��>/�{O�`>jl��~!&t7e*޵��Wh2��y�5��Jl	NL�����yν�䈐C���[��<=6�ATO:j��*sf��ߗD�U3�f���o�Q�vH�\:�;��}���n�M5$�{T���A�\��=p�|pb�������,aKbP�B�o/�s �f�'P���.�s��Iv�[;��� ��!q��J=��b=ٌ�:h"�;������3�U��r3��,�G���g���"����� ��=�����U6�����8)�E�.�T1v��G���QD�P�DLy��KȎ���>q��p���/z���c�2we�ѱ����La����=p�C�����6��� Vp�>�%)�Ѻ��M@��D'zdL���`L���V���6�`O��ĉ���X�n;��i�Pe��s}���(#b;��O_� $�v����z(l't%�`�
wD���{Y�ܻ�u�O�p�/ǀ�)���2�Rך���*��By�4/raA��,�H��_�g�e������U#���x;�*�APSlR������]'ل� V��amF3�ozd"���U�c�(��Z���dr�V�i~�~��!���B�[�: �;�&%���jS�����=5���I*��"��2G�	�Y�\��cA/���L5	���o��� `�� er�\�1<��6a�J�Q���DRӁGl?�pN0T�m��-u8[���B��m�u�|�.�	3�j���/q�w�lN��eȌ�)�vq���^ �����3}��i��-$�0���!j1QO���� ��C~1�Ugx������V���`�:jF���ǋŠ��X���Ƥ���.��>�&YoD��w������h�h�ۙ�2B��Z��oV��Y�,we�Ի�yQ}��[����'P�7	�tų%�g�Q͇e[�>�Ɓ��˞��l�3)������KX%���X@��ve�~ԯ�\�,b�(ԙ�������m'݁�z$XH�~� t���:��O�Ɇ6�_s���خ�:�![?-�;ث`"���O	M oy�]��#GN�/d����x�P\!C�H���<�6(&� �Q�D�\o��t��"����w��f���¹Zn�4�OM|�Ԁ/��u�#�w�fJշ	�n���q��	�2 劘wi�\#]g	�Zo�����S��+)y��C%�t��X��Q!/d��	k�M�n�A�C�1�hĺ�_t�}V��DX��`c\�U��jL&n �/	�
`tx�;�"��B�Eo�7�@/�x@x�}���4��_�0�ڣ���R&&�@���6d�U�/��y߄aw6�k����i������2[0�4���_��\�C}����ʵ��N/�[�̰�����sx���C�!�x��E�Υ\F�9�v���>��f�TX�ln8O��_�h~K��0���+�WX�k���YP�i'�+�W��'��V�*h6��U���3���#g��*�w;e�w�s�2d���H�E��S`���@r��-KAﺇ���������E=�S��N��5517�>p���qc%f��Σ���2I�Q? vO�V���?��\�:�h�B=v +�l���ؘr����gܠѮx>�ýiNҡ���e*�����?|�3�e ��Q�� ��1�T�������B��%"m�|��ΏSb2/)�RR�
"�a`j�nQ��b�[͚��ױr��Z͋WC!:+$�O	��qE�w��xn��>`��h	�Ћ�� ��g����u�Ю��	��e���4��X���� ��	��n��[�3�Z �El�ee��u�]��������IMF�X���>X)�d)���0�-���+��È�ָ���亂8<�hB��TbB�p�o���'�.p}7�����794�C�M�VО�I�;y(�Kf�I2�W�A���a�����8����&�-��EH'�7��L��aH�����B��T(�[�r��gxɫ����ㅿ2լ_c��`	���_���ǘ�'0(֭K�"�T�$���{�k|7
�Y�������N����W��zʏ��FX��SOs��W�]��V-�g��;��_�a.t����Z�r�V���@U��aA��$���V�A^�X��]����߭�����6j���e1����m	K��$fR*���� l�ԁ�Fϴ����v��a׭�M1ߵDV��k���.!d5uV:�f��mo_�1�T[>a �f&��̹5�a�I�b�]��h~h����;�P����i�{;Is��1�r������q�״��P;/���E��I�4�<�����T���>��`qID�?kyq%���#h��ROn0\@wK+��p~Mrh_P:�ټ��a��d�/�����	���P�����`���z��C;3d������7Z_�V$�:š��D���I�!��)髥]#�a\��7�^m<��T�(7�x�E����Wb�798�Y��UZ	3�������ǰ��
���^�,����;��Uxh�E
�T�2w�v�����Rx?����i
�PE���q��}��>���	~��F��E�(m�-�F�f)W��i�����$�(v�����\!g�5����-L����&
��Z�Zv�e������чVӢ
R�g�a�ғj���C���ō���+3�vmb����yv���.��w�L5ع"[%s�CEy�H,�{�������v�����_���/�b���zk�x��`�_
��9���>�c�V�F�w"oHǊ�)2��H  z_m/���o�E�@�
�D�YzG�0���P6��5]A����|͒q8�x^Th�X�� �k�����Q<|;Ħ��#_@`�'����X��m^�3.q��������j(r�<�5�u�VY�E���u��%6�}7�p��r󠟽e��!mEC<u�i@/�Ȟ�xa=��f+����!���Ef�=J�J-��!��n�ϻO�n�r��\�T�X~:&X�RB3�����t����μ����p*#�>�9`�@�#�<��V!3��Y��1:vOc���Y��B&�鳞�c�r���w�>���;]�O=��d5��JW�8���g'�^u��~J\�V�'�h�����c[�b9�{V�G�k���B:�,���d������]ʏ��"4}Z��E=��6������������N�ڼ��Q�ʮ.�j�/��ۖ>�i�F�*]"o��B��&�&�e-��_'R+�^8Θs���Tn�cНhq,͕�Z%n"����؈�ߛ5�w�vd�ɕ�K��~k�d�!�DK�/ώ�1���<5�H��G�-��3M�
u�3w83�E���׸�owQ�t��'�K�gQ�K�QTgѕ�Cpjܪ�����Xg'4�v�H5OE枋�`�э�S��MD��7�0�A价͉���M�5{{���;d�����<tN�(��0q��ܷY�dH�T�A�/\����_(h�Rk:g7�.Va���)��[�n:�I)U�������Y)�t�e�.gnkM	4����)
U�a#���p�V:(�&��\1c_dޮU$��&7J1�����B��
Koͼ+WE9�J2Ǒ�͘�q�Yd�V}�K�c���w��]S�AA]4;�Bn�H��,�>�+�X�MNM:W$����i!���&����Wq�����):i�j6a�RNK����l��J78m�(`�tt�=wB1p���3�t抳��3t��?䱆�j_c�5�x����@��*��(�\X�{�����F��Z��� ��J�.� &�-���Ud�7J6,ezF��¬�CN������P,�	] �O}�����`Q#�̬2+�;��	��A�@���V'mMM=�Z���(09V��	
	^�V���/�����ׄ��"�$��|�Z=�DF`�T��ߍ�c���5Jx��s�g��qt2y�/�%����A��ض��l�u����p߼xi��]���h��P��I���%����䜬P�Mo�u��IrR�ؑ�R���������l�!I�N=Қ���ɣ���8��
C�0"1�f9`&3|o`��1�_��Fv ��:�/���	��ϝJ�x�1���娜r[y���rR�%�@��TB���^��M��QYDL��Zp.ٙ_#+��ML��/Ė�q�g���vFWm����ݩa�y���~ �G�$�!ѻ*^6��ی8`�4&̄>��ȳ�������F��c�[�#����?��n�ia}�&^��8��Q�T�pW�Dc��G���n0�1�?;Y��K:��c:>�NN�pݏ[�iN�4u�@<	�]���_���J�*���7�Rw�������C���&�Iz��pV�W��R�d5��r"��z�=[j�����Ne�c��Q@qxd����;�`���4�v�L������)KXI;��i�TE1ז�[��Pa&9#�ښ(���{��3W,����U�d5�B�м�{=��^�p���29q�˓�h�1��T���w}����T��B�sJ_ȓ1c�o	+��`�AĿ㪖�p������8*�H�nP����:+~dG��ez�s+��DB{�G�v�@�vIL�;l��1+�O}9���4�����߇Ń�x��lHn�A�\0(Ft����j����i��!+g��!.�XU�,���ŭ)� %� m#�r�+]v"��)oaG[�� ҃���f�#���g�n�v�ύ��.��!���ș�_�����q�����v�c믞y�;�ÿ��5��]�?ҎM��8�F��;0��c��Dt�ӂ�j2���V�\v�E�eI
1`���Lv�W&������4ᣢ;|���0a�����|��s�e�t>)G�����WC��4i0�����;A�F���1�T��'ҧ����}B�Vl���A�2?-hlx��X�G�E*hpDk����r�\η�+�$��e�x���\�$���`Y������g�����[t�M�1-����]�Ǚ�[�ڈ����c~e��J�?�	<	�Y�l���U�ȋ �\�2����L3���D��At9N�6�
���&�ݡ�.@� ng�8ӲT�tZ��-&Vr�@�w�ǒ��+�"��hn}��Xp�fD������t�~'�F��Z�l�,���1�)�-˅x�J	><�9s���Q���_z��c��$�_����<yP���_Qk�Uz�y�6�mb���^HF�$�N�K��`G��P���]ˈ��F�������bZ�w��=����O<�����;�,������JA��S��k���A������^(EY�u��8:�hE�K�A�v9 ;��B2u�3�䲃Z .��CgJ�q��n�h!�5�+r��7w�˥-��}�l��^O����X�����ک.Y�t�O]��x�5���N���E�Opj¡�;X�x��'�,�H.��}"���Y�_����OgҊA�Dh���{H�����=�z��Boʕ��@!C�HjPg�	�%��q_��-�ǩ�/����̾a�p$��]R�m�)�\C��5�����P��ľ)�j@ar�����^j�dO/������浦����3n~�1j/Y,g�4��=ӑ"��p���o� �����C"XN��8S�7��٢�|l.�Ϡؗ/���'�����n�V�.��.w�"S��B�4E"Q�� ^��E��mG�C��H]�|���G�� ���r���]�2ŭOȆg���Y�h��
��cO@���ш:����*�.���y�_�l���) �aђG�ö�c��p-�1P�X��C��\�\�qbƩ�B���Ew��}ݖdщ�=�5_p;�>�3��/pw��B�_ض����1���b:g�#��L]�n��>}��M�Sqʉ�R����/)�G�� S�Qƪ�������Z��D����ڢ������ �D�Č/�*��ۭ��C�D�30����C�0��z�9�),�{�F���ntڙ6C&rH@�����{=���1W��^�X�sv������o��^��垺	��L�剌���h"�oc���ݻ%�b)�p�;mZaH�&_�(Lft�i-����Hv�t����� f�э�H{��i:���I�7�m�G�Jnq�k�!>&�@s�F$o�T+9���-L|â�Pl�tl�����I��&Bb�q�&8IC��!Rx=]!Զʸ;x����Ɖ����>�z�8�{����ԬO9CZ1{ӛ�w��/���F�7����%OIvmSb���:-F&1QT���&��&u~�l��	|Yn�#���D]bz�j{�Eteٕ��gQ�J�l��F7��⢸�s�D�`���#t�Ⳃ!�@f��M9��ª�>^�Bp[q�Cf��I�p�t�r��砑TE죌0���"G��<��5`��޶��W��.9�Ӫ�Q�|���n�K��(���"�>��f �����5�m_�X�ˍ�x!ױRF1(�:���tx�W��'�b����(^c�aYm�yB��ս��(�g�+ _�]/�G:n#�Ĺ�������[���>o8䋠��X^X���S	���v2��%<T��s;=07�7�7�Ѽ��͠K�%��-:Z�|�$HOg����t���/bc?ϧ�٨b�a� ��]���?JR��n'w�>*O��!X�?fhOe��-_�(��)���V�5����{�u��Zj����(��n��~+p���ԗFz��e�g�������<z+.J�ET���\��彣�̂�6kU'�t�nX�te��<�i����SWrx�+�S�9�;5��W"��r��yF3д�l�oD5[��=n�5���0�,��4rJ�S�,R��OL���z2����:]0*��]F-�&��W�BtqZ/L�^��:a��X>���d�)�yX)���p��χh8d��w�v��vv�E�uqnԠ�Ə�������K���U��(��6*��yhJ����k�!��Ѱ��T�7�S��i{lUO�ŸR3�=�%�n�]��<sʌ6���s���ռfrxt��\A�J�)�l��
�R2\G�o�����5�Thmy�eO�L#I�`���C��L�`/]혙 �
LЋ�8��d�~�"3�3=��{���z
�FSo�������sP��7db��w0_Rt�v���,�0Q���1�15sK�i�Cj��i�tT�b�����b�wi��:m4S�}�v܇X�JSh�V�g?�&X�J�����7�t��;eP��tj�v_�p����?:I_Ӷ��K��z*n�J�&눊�&lA3z6N�1�);Hd�i�oؿL�JK��T� q����F]�g�� 7L�����DrV�'Β�j�w�lJ�=g�au����zI���tl��J�7�ˀzCYx��O#��@�bVL�{��x�>��ʿ�V	���h#�����4s���-���2uy�aP���7R���h�Y�Ŷ�KFvށO�����҈�6 ��g���"*Q�7yȲQ����)q0�������P�ۧѭ?���n�b��'�)z�i�K���@��M,6���4���Dt�@�����L��TvsT�����Е�M�+��)