��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�8k�)9�k���J�f ۘEN�R��>�Ug:�&�1�a4ⳉ&<h9�	�(ds�X��X�ɥ�*"Ǻ���d��f҈�1d_;|lƦ���1B�K�b�}hTK�|�Œ��՛JKF�zMLdv��#��-�r�{��Q���)�:�ӳ�Q���.&Q��[�ũRf|XB?�t0�,ɒw��I��N��!$����M4�b_�_I(������R���GE?36'��a{B��軪��U��h����x~��������D�S�����~��΍�
D�IsE��N����A'��KAZ�K�h=�)�� �XJ�������)8�PX�~0�YyYo�{�l� ����z`�t��o�(��}I�J+�t<c�oa�r��/��7��A�y��~��%��칮�+���)����u�X�\35$�~�PJ���Rp�A����*�Ц�W�ǌ��s�C*��j��J�s,|�{�d�q��d�����hΦள�E4v�rs�ۈ����2�P�NM'��o�}�Cn(�^</���5,�s�4��C{�#�
������6�"��.���M�'��`�H����T6G�R��K9(���v�ߋ(}�z-��P�|�)'��I�πp���߇v���,�X6K��/rDV����� "�@`�52��R�v7M���e��ʂB14J�]5���AO(����*{����ղ��AmrD��_�O6��ݕ�
j�ɡK;Vֻ�$M�������4���r8�?�v�T]|I��
/�˲o���������+�x�.�@[��J��l5�X+�/����u�J4˲��2'�W�3s�[���m�3�~Vd�2b��:��\���3�/������ �a� i{˿t�'��v�&9S~Ym~F����R�1�t�U������V�鷻y3T{7-8j��AcXl7B���k�u���JlX�?Q��:耍�h��H��G���Q=��_�Վi&�=��z����E=�$Z����  +i)&�M�s~%�Y���6���VV^�B�=��˺����ʱI�O7�m��yW����$^Me4c���N ��#r*oP�4���W���;5�=/$I¤N���:��HS��Q4���=��>��|���a����b�נΨ�qLtf�}����_���Y���e�1'Z��e��B�w��xϖtմ�L�˚>��'�l�w?�$�AIZ1f1��@;����XdŦΏ`�2ݑ�&84F��PZWv�\I�6¦�$
����V@Žn����#�eU��^s�{qr>�D1��2����Ql���\�X���ij�قY���צu�skwJ��ٳ����H]�i q�'5� i(k�)��9S�k J@ݼ��-������*U[������֞�6Y�O�;I�{2雀��=H��_�~�x(��I�s���A�34Z��';P��?hH5�9'��wĢ���>ZF%&}�0C�2 sxu��Fq����+���D5~^���md�*��7�� fh�V��S�kTT����)��nO)��j���Q�<�P��c4ƺݭ7�	~�"�k�#�E�]t��wX�lҐ���I`ؗ�^����H��|�,R��'�����v��>fm���g��3�饜\��þ���tmu�>`�a'��8F���/j�q��Ϥ�Zm`�����������`)�%��^I���xb��J@^OO�upt�J?hBo��V�c��þ��7�a�Mw��*�p2)N$V<��v����w���)�0U�Ks�N+�S���{s�2{�Ce ��W�h���u@%ۍ ]%-�6u�(��i��~��N�M��;�)ZS��K�:x�dm�q�\M2^��1qttd�A�x���!+�<b���x;��-4e������M�w��F��3�Q[�[Q����8�f��<��N5@�$5c�*�X�>�^Ҝ����M��l����{��td�*T1U��@6�qFO����2-z�AD����T�~���<3��$�x�E�:`_�@#Y:��}yNb.��$��uv�:yk/u��4)�����5eAA�m��,��
	[��O��М��4��2������I<�F��>�����Z�U������X����~<���W��o8c��%X�X��̝OfR�g4y<�p�Α4&Wjn"J	c��P�z�PO��!V@ul�l��ߊȾ�ᖯ'6�KTܧ�cيK,*K ����<)bb1	i4!�����^�9�	�{�Ј��7���Ҡ���t'�ۻ�"��G;�1�%wg(r_�����H5�?��w�����ޏ�IQ�O��ɹ��8X�O�&�T$�.,q���g�tr!��W3C�*�:�j��gY�-�r�����&Фb�=��W�L�
����C�zmnW)q��qD���4�(²N�Aa�M�"��H�'��?߯u+��)�z��N3��~�o��� �a��l���D�"�t�ʲ�6��q41 ���<���Kɕ	�x%~�S���
j�C�j����Q�o�B������h��y���g����oe�e�I=qN��Z��	��<A-�a�����W��z��8p���HDO���Ng@ij��R*<����Q��s�1D���R0�:9O�$���Ã����F#�2��L��Sm�d򒀟o�w֤�nk�]�@���ָd��$cC�A|��ǲ3Ix�*��d��w)p�K��j�s����oR\d���a��-v�L_�=\���4�9n۵J��/���%�^�IIQ[�H5Y�$�	�c��ߍ���)��X���b��<E���8��q�=��W@��)��	�(���O?"�)7V��0���5��I5��n[`�"�Q�S�$ ���1$�-r5�X���>kX�@	IS~��D�����g�ӵ6�s�?':X��;�w��%�*M�~��(��V�'�XI��Ck�a�ꀒۭ���Y� "�d�V�Ҙ���1����t/�ף 8��L���R�`σ��%U��s����A�-���,���B�ޫ�<re�FQj�Rh���W}Kf3�C�2��%�?���P�Ou��I���k��rp)���9�unoIp;.pM�"f���s�/�]����֛� ��lv��Sѐ���ץhZ�=��]o�d6���!D��Ѹd��� �kDط�:���֪�ɟ.�0��A]NGí�uK��*�o �6}�]�R��%�{��Tq�pE��5��c�uQ�+�͝��5�#ف�X��V_���@uc�
kA<ŖסyG����L������ݳ��%�L��,'E��7�c�p�$9�go���4`s �j�:V�Ka�m��:mJ��)���D��q�hC�ٶ�:�d��n@�fo#�ON��}�^���Fô-��s��-���y���,#kg"_����o��1҂7o��c��8�:��p��	$��/�/>��`\�cu����ؗ���i�Pdw��ڴ��h�d\������������UA��F�^| ���<�A����\��"��	�<(B���t�w�6�WT��$c��N?fP<����
^dr��"��
ǀם�4�?|�lm!� >� �J_�U�Gߘ��{R�g/跳Js
Y��~�>9�`Z���2=���]��$���ώ���� �߸ٮ�CͩTT�\�������?لh˘'�	������P��|jT��Y�"=l4,��3�,Њ�9%�}�L뫃2?{���ѶAȋD\��Y��)��J����Jܲ}�����5���xJ�
�0U���~H�A������E;th���O�Q�k���zSc�y�Q����ޒ4)vS��Q"���?2)g�^8�յQ�՞W�6lѩ�߉���y���][�,^
h�ԤƱn}-���Q����)҆��!~5����R+k]^L�sC a�'E�X���nG�����R��Rӡ���p �F��d
�	v��b���#;��'4OV:tޭ��.xr�����ju����,�u����4}�a��L�;��\�)d�Z]SLhZ���+�i����Gl����k�Hd�N���1½'	��l��Z���#���<60� �%�.��#O�(T� Q����V�iD9������J��o|=V�!-�v!�G'[$�g�3�*�K${���&�M- ЯS��O>{K��l��S"*aDX�]��.��VNvR��t4j��k�j�w��/{uxD��l�����j���W{�o��)�$���x��3�<�Q�M��ęp)/�-Z��T�)��Bb�B!�B��ܽN���e1����}?�N��7��%��j7��U�J��E�m���q�u�LR��R_�忂������P�������j��oEX�������|�������̴��2�f{�z5j6쀅��2�_l���g�^w�M�qҶJP��)���d|�	[8oX�#H3�|��:����-ǁ!�SKjps��j��H�򔫶V��� o��h��MJ6"����4��W��+��>���*�ѥ�#��gZ'�=qI?�������_<(g3'�Y�Ty�PyZ�Q�fԭ,��SP-§�˚!���_c�i5��Q�����u���mo��lm�@�F����@PD'`��i7�Ce���2�K�぀����p#��K�U�<�?��0n�ϗ~�V�;=��t���4����d�n�9[�����Q
��/-r;<$�lP��٬Df�T�;wy	��t��Z�9y�� �0 h^"�v�ét����s��"(�޾Wr���^������b�I�V3g��R{�O!I5�0���W�0)� �aԐ;�ٚ�*&h�����ۜ�k��2=�}�&	�5\,g�LҦV��F���{��7�*9"���'K�oBf);�NO�'�LM����|�<׀��ԍo��w��^ԙ�[t�o��(�}�:~������Z,�sO���u1	`N�Up:�rGc�6 U�9zn��ρ'��v�����U���oD-f>|��R�Ҟ���;l���{���Its��dM��s���/�|�3W9�g�J俁�ESL6��.[ݸ`��[���׌�\Ji]�O�p�=��o�T����Gto�%ay�=��v��[t%�+A�GoZ�\�O�w5= ��3��T��X��� ��}���5�-��3y��p��n^~���u9;� ���a��f�����@��"�;ލ*��6�ԡ��uk��'�?��&��?`N�%d/�������̓����J�K�D�Q��`>S�~늧����v��/��#�e����t9���K#�,�+��j�0�L/8zn�mZI!L�`��A�ѩ:`{~�&� ��!���p�,u��U�U������畁ޗ�)0���v�78��7,U_��Y�V/Fi��d�k6O��[i�=��!X�߿����n���l󽊼�a��Ae�L�^���d�d��f!��љ%��cp�fF��:ɀ*ة_Nl��-�h�mB�I�eq��w_sͧC�%�&)�L�q؅* �_%Ƹ+ׇ��s#-kC"P�ъ��o��^����%U�Q�c���(��p�{;,Z�.�����\_#{��R�X�?�[ِÊ�9Tv�R��/�_��X2�t�6x�aHT����<$#�լ��LW̓�G�j�"831�J�؃�?�j����9u*;г�q��w���|u�/T���v��v V�?����$����|�v�������u.��ּqWu�x�yd����+�G,��)��o!HS�/�چC�tD~ax:�Å��Y�^�:q�a�kOOAƫr�w���j�%$L+��Y�@��R5}���&2R��"v�hn��h�h��we/RM��zT읱��޽w�z�Z36n���< O�܌t�99� �� �U�Uՠ-x_,�e��������3(�MM��r�d��^��UԌd��2�)�>e�����.<��"�d�]�\+�L٠��/[��1~y�eÖ���3S&Ems��#�c5yb�J�q`]+���.����%�>&M��5*74�^��7��%��9�Ϳʏ���v���m�4�5�w�O s��8Δm��fX!'�;g.�x���U��4��*��Z�R�:���`�H~)m)i�W�s�k��ڻ1��Î����7�^bEяUAp��.�������[ܽ��+��p&�߈3<�;X�X-��z�Z̯N��Q���D�P�6��s�A�
�1�#���F���fQs]�]��,F�,6�LLt[��f?��� (x�3Lϩ�q��F�"�u��N�z���7����TW`����� �	]2���P9�e�LE�=Kȫ�*&И��B�z�"]9������F��X�	N�����f}�L����m���&]�I������G=EXeq�$`^Z����*�ĲE�x�Ap�0�R�Un/��r�eC����lA��z��{��1�q�Q8���@��u�:t���5��DOI"�����6�^�N�P	Y��.U��������xL2����
4_ 2�|f�ﰡ.�DbFQe����@�5=�^��W7���t~E�_Q��%��e� ��o�O��Id��􂷣����&�P�+����]�v�'�����c�(�Y6/��> �羽7� I�%� pUp�-g�5(�t4e��6�nL������%h�������E��%�E:�}��O�P���W�
���b����?yo_��.�ķph/Ԟ�y��+Fߑ���UpT��7"mG�F� ��\��s����_[7_vn�HX�}�jD��s�by9t(�f[���n�E��o�>u3��te�,�,#YX7����.sg�A;H�3�.C���T�!1��Sd�iyKت�c����Ŧ��/=6���j�^Bv�2V��
��o熵�X�_㛾3�2D���_s&���q�-$x�/$Nx����e/��	O��)�͌�,uKh.P�o���\z��Rѣ�l�`3~*�p��D�S��T�vkx�TqDh���f��3�K}�b8��r���
�A,c]�l�
C����}v�f�3¡R��
rA�pE�.����X���ڀ:腝���Fvʂ;#0���8��ԍE�AjC���7N��;��Ӳ"��tQ��o`Q/��9M)��r(Ϡte�Iz���TD��M�C���P9tr��8��ptpk�q͌���w(�ez�W��K�ԇ;�5r����)�8���I�Q���*���̜�՟'	r���y����xw0��N��yqM�L�gh�$��	��Ѝx�38
V�b 4��<f�@FKV���\d]C��O��=���
!�B��=x�'�*��in}[�ca��2�e}�UG�J�9s�fs�s�{"&�ϖ_����^x�GG�1qȾ�CX��.oH���_˘�b�y%���k. Di/6{q��2�,�3�z��}0�#����T.̺u)�[z�=�T	���:�L�_�{�J, ��6h뉁��i��yO�A���4-�n(&LA�ۼ��vżO]��vO#��`EL�=]� )��IP�M �'�|}~FP }y�d��|������܊@φ3�P����j�7��O�^��M�F�&S"���4�C^I��e֤L�N��h���˱��)�G�l�����#���Zx#g�� ,� ;��qpUX$4-2����ޚ�L�9m�xLoJ��e�3���ڒq�x9N�H�Jn��ȕ��z=�� é�L��߆���/���2�^z��;�b
#��������S��ШΩ��D��x�D6�pJc4t־�R<&�����"aTc-yT��,����-�T��m��q� o���o�����"*��4	w;�6F垠��X�wt���m���h[A�#��ǭ��D�f}۹�������RI���a��7q��-�9^�X1�/���Ј2�UJ���E\@��͂u�H��5�����v�ԒZ�t��V�P�$w4}1vH�����a�`q�aI�uH6�
g��+$á%4���P`�1�Q�<Wِ�eo�	�3�`����'܁*툣Zn}�*�7��,�$�Z��wPj���IeK���=[2ɮ[��G��%&v̙
���abJ�,z�se�ǭS���(ڤ]��\jq�Ne�,Y�Z\!%ӞS�ϛv���eI>ʛ�X�}�J��&�W\oG޻�h6��e!m����LO�}�1)w
�s閏�ɽ��(�Q<�*�kN`�#�cqO`1��e�r�=�r]�K��K�o���Ȥ��������'�p;"3�g�%�{�3�s�/Ơ���(���� �g�W�W6q/p�iG���g��7� vm �.����?��z��>�6�쉱����A� =*�亾-\�-�\��k�;F��	xY?y�wDw�1��\/�W�U+D��V�G�lB����o�#pa�A��.5wS�?D�/�nsZ�����u��di0��u��,H�ۜ^�������ͷЄ8�)a�����ί�2[I�30d��g�>W����U��岼� �;鼩;�\�x#��X</�E?���2"ƃ��Ǒ�[�@ �G&�%c�G���C�C!j�YH���3�~o�)�������)��q����9	�}?��Wng��� �Ϟ���-�X'�zߊ����B�h�P�W���kB���>Pi�)͇�J��.�A���/����3vF>	���ůcq?���'B��%���h�?4�(��ˆ�uC��/�9P�js�4C.���g�#�N&�l��l�!��r&�h7�w�1��`��?� �dk��W�63�$9�k#В_�\�nŒ-�#�%��'�u;�1og,��oo4z�s�T:0_ �h�ٿ�՗e� �3���� �|G���^�ldz�3�r����]�vc���\�w`�VK?��=��Z��Pr��2���0$j?y�^}�z��Ԫ9>O�TJ�b�1����\JFB��6�����脿�ȴS�[�����m��O��L_�B���|�1��G���&7�z$�m[=(�1�|c�F��{#aX/��F�d��U[u*���cBb�}�
9�a'HZ|V^��A�0�B����P�8��Aq��r�er� �/T\>s�)}e�a���EJ���ֵ/�l����4���i���n�g��|���-!�B����B#Y��e���C�_���x���&=�W�'Y�c²��#�� �CRX���A�侎�P��v�$>��;I}U�7`�tG@(D���3�`|�h��v��Q�O�p�h̜�;�Y_s�M��e@@�!��ʂd��hTt�4 +��y�ӬY��S�<K�6~�?};��C���t�R� ��-��2��c�;�F����p��@��}���Txɔ���?x
��k�	�ӥ&�~���űPh����nO-��`SX�,LNk�6}L!*ŗ�v����t�ǂ���H�x���;�p2[�f���UZi���WƁ\D�2̝�*1��� ���@e�����ц��:��P��`���d:n�����+[)�z]n�ݝ�"�~����+��`�D�=:]����f��P�g`yj.D^z��F�nMv�cg���XM�E�'\�g ����<��7�*��}�R��Ã+F��%6�,���pdE<>V�:�3�&y^�ח.��i�6?^�Κ+��>.���.(��ؤZ�k.���C<̹���@� 3�E�Ȏ�?,%�L��]j�����j�"� ll��#ٵ�݀��.(4*��!��b%��VX0W��lv��)9Б�t��)&�H-ˋ����n�j��>@����)��>N �]���>�ꅴ��d��hVO�~^a	����9K���F�+K�Zy�^)�^���ᷘ��A)O��%���p���A��jh��)��֔�����R��q*�B��B�=��m��uNBQ5�c�Y�~;G�Ւ4fb�t��s�'�	k��.*̍����*9�넥���ٱ��itbT?�\[��q���k��Њ���rֆ�!j�pП'6����{,"[n��F�!t��T�
��0�i:fZA�v���W��,��+,%{[ѽ3Jyt§��|���"�]�(�w��k	��,��*��<[2{`�;2��;���{�5A\<���+Ȥ��Հ�����C�|d@J��0�����Q�b��堧ɤL��3hɓS�C�@�2���]ȅ����M^N3�m󌈤8�̷?��3���C�i2���1�n��E�%�S��1NKؼE�{�T�+Y?X�n��|�k�P(jΰd}SH�ƞ���n���b���ŏ	mc �7����${��l�V7������'�O���1���:$\�2��6P�A���pwd9O�
m���	�>��1���'`v9R�Z�\aw�jdA-Ņ�0d_��h�"1ۢiB�eNZ��@ ��g��/�5�N�#�������@i��bԮE� ��&jemxQ:�ၤΖ�>��&��T� :)v9ԗ�$�Zf(������r`e�s�v�K�Y�Vl:T�4h���%DZ�g<�9��R�8��t�j+wA���u�Jҗ�]v0;�V��w���mn��F�� @�%�i&����;d�<f#��.�=U���
�h���)�u~#�����MD�eJ!o��	�o6V���1����3��X����!�|�� l�l��>�N|��i]�n��B2�0Ap��2�^�Pn�pfɬ7�oo���b�������ڦj�.�m���d�^����f�Hu.��s2+Z�T�3�YmfU%����=����@�x�5x���'s�!��h��I��T��%��,���,�/�Ď���×�:Ow�.A Z�c����o ��D�<9����v�����o��6JY��ɑ1�����-5���qݣ������N`wi��d\��x����o2��/��N�\����tՁ}=l�x�w"��r�����x:���%���X�T����uAPo(#_¬�p���i$�;��R|zC^��m���t�� Կ(�7.��*:f��'Tj�H��8܅9���Q���O^wg��Z��ߨ��w�����%����?� rcM�$���u�~�1�dx������0�� Ղ��#O:�ֈ�'T�S�3�C�SM
�e�܄?/&���zDV�Ӟ+����x�}����{bJ��Aŋ9��m��|�FC_<�MI=)�	"W���*�!�褚Y%]5nڶ�*����2B9w6��N��aJyC�W5�ֱ�x�k�~uG���bY��d�$s� l_-�D���7�޶ou������s���������� ��j_�O�G����c�4b(�PB#H������E/7�^,J����B�ӱ�]l�f.ʒ|�
�+E+��ի+�tǗt1Y���\�8����ۻ�	$�6X��_4����"�����{�1j�w�C���7�Ola�`�� ɾ'M�)���]ܣA�yd���9Œ6�6��3�QJ&�Z���"A�X<h�8�����f�u�mc.yn�(�iig����ý��j��ܞv� ��R���;I�US`�N�Ҕ4���U���%�db$��6��Ϸ���̗�/v��$���#���l�������k	~A�!��^OD��i��V��4Ξŭ�b;��	c�R^��G3&��+`pվOے�4��sb��eVQ��H]��b�ʛV��b�����0��ND����Xܾ6G�:7�Dc\̜y|M
}��'}�� ��U�(�[B�R��Hu�����eݕrqT^^l��&���]�Þ�iߜOisT�����t?��"��P��M\�zO'R�Z���u�,��Ê�؜ o�M��d�ǥ�M*r�����L#�rM9�`�]�N���&�t������H$�ߦ�>����+C����i��Q���LXr�.5�ee�mY9���:�{6�}Cs�z�8�j�gW]��k�`�r mzj��%��e�%%;������	�ְJ���c[�[ � !���~�,��$z������#�d�~~��>�)\��j��q��:R�	��\��G@��M��GV��3�
���z��"2�l��M�-N�Nq|�_[�B(��X�!�c4����Ǽe�a��X��������Xt=�ĩ!�Ѹ���ŝ����u`�E��\�e�����a���9����ûc8ǻ:T��Q�����>�z@�u���A7�G�j��f{�)��m��V��~��ȏ~3���Lɓ� �Gi� �fl*c����e�a���?�T4����?�@^UB�(/�F�v鬗�1�I�Ӑ˝�I d�?��@�� �[fW~|{ر��]�h��W��/@�#���_&7�ĭ�uq��[�GT�f��'�
�T&>. x��7I�g��xw}��%�9+&'����1���12��Z�΍�(͎'�Bf�){�c0��"8=S�C��w�:NĂ�x� ��������Qe@��^�2��p�c�]wW��h��ֵv��iE	��tΌ��S�֦b�<�]��
��U?W9;Ϝ\A$�*d�溘�4$�Iet=k�Yk�l��`r��K'�[��q� �>�'���p^�[��E�w�!�(&YI]���<��*��0��B���8+�shQ�J-yΒ��m2��>�Uls�g�n�w�w�҈V{TK�M��i���Hb ʛ�[�����e�lz�e/>!�Ϗ���Fb�|lz3�����!���	��u�!dmrs���Qǳ�����Gm�N���-�'�%LK�[���t��&�s����y&=U$�7Mh[�+���a�}�f\��c��>"����W��8}x#�{�턣��T�F����MG��	,³-7�f�9��$�xC5�PC�r�������g�~u\J��.�Dó���Zǭ��%�xԝg��@y��ԃ���w�Z�vL��ȫ�xÙ�ԠY��˹ϡ6q��2��:�N�L�De�O1݆Z��RJ��L[�0t�Z}3�����]��1���(��$5��9����Y,����,�e;��cG�B���s��l7ViRM���@x�K7�9(,qud]����PY@4Fo��oy$R��~��x�V��Gjί"����Y+Ջ]yyh5��ɹ$c�)��9�1�j�e�_��Lo�P1@j�#���j��)�z7z���h�b���G���P��*q��)��I_�8#�d�^�A�1�S��Qm_�G#"��Ed&��_ܒx2J�5���P����|`�ln�	`����OQ͊Sh\đ>��8"����辉7�<pV��c0����e���7p�9�{�zɕcՐ��ovk��XR���'ȍ�ہ���d�h.��Eg4os"��	ݟ>�i9<�6�W������rԑ��l�aG;���2��-&L�l	�`��A���+��Ǐ��2����u�S�vN�R���>Ѫ�����ԝ��R�d������;��!���{�y"z� ����т\�捎��A�:�j�5�olH����@H��E�>� ��ћF��;:D؊h���UL�n�O�gꥍ�)z���Ĳ��iؑ"	8�K�6�=ſ$�0v��
i���R�
�[��I<���Pz��O��
K��-����]ǎ�����G�ɇ���:��A���x�axy������j��0vp��O��B�����r Z+�om� �ҶZ��'�t@(�6|ş��jF�q%8�b�>�%����?�㵇'���Ga���Gc����Aވ�V1%�Y��u�,���jx/��W%5&t(�����o�m�
E���S�"ZBL�6;�b�f�FW��-D9|�j�
j!;�e���=��=��lI�\�Q�ᣝ/����n����aŚn}�>����=g �"#��y��l��̡�#��'����8GE��<���N�w�5P��/T��>(� "m�%�z��2���χ2����h� �@�w.m�/�@1����
Oh�ԑ��B$ �rʿ ��/µ��� ��@W+;�Rc��a�4#�;e��:d�Jğ5�-hc�nLH%D�!�����Q�B��	=Y�bVr�yE�����re�֡F��w_�)V���Xs&��Ԇ��@L9"���ec�U[٨&�kl2�28���RLp�v��u�=�^z�-��'� ���F�q�Ɯ��4�e����J[p��̶�u2�����#;}Ω�����u��=$;�r��=Ȱ0�N�<�_+2�*j����')�!�1kQ?NG�9�x@4%�L��n�f�% ������h� �]h_�ڼ-/*9�K�!�_ Ŕ�6��B�ؘ�T�m�x�������I8����,/;���5k|�μM$�k}Sе\���(~�Y��o��B�{� ��PҼk��¤�O3��ȃ���A������`v�q}6�H�H�~�s���P�vY#��@4���L�[�!�_�6���Diӷ�Y�1�k�4Q��~���$vK�Z���D���ϡ��@�i��
Y��`�{���-¸yh���Eaȭ/�˻��7�8�y���H)r�h�s�cW%����P��'�6���Jˮ��,�ٚl��}�����i5��#i�K�(?¬m�hzX��=;�B��'n*oӖxc�����Hi�	�ֆf�Z,x33H�%�nik���pRo�<��9��ƫ �t�/����?��v�uk�>S�>���g���\|z��܏:Dd�p��-/���Ŏ�Mٛj���\' �xND� �$!b)�btq��>`W��̟��m+��O�a��Y�g�X^Ⱥ1�Q�JMX7N�D��|"�Yì_��c�Z���J��a�$-���+[���]����F���-�����'���x�IvK�1��H���U�l����I�O�1s#�уA>U����\ھ$j����U©H�~�Xʼ��'���/��Yq8����KV��3�,��mW 3>'_p�qk5&��e����=I���H "�5,88�������a��W؏����w�ȱVR6ث]0�`���'�9�V�ٲ����ֵC�����j��Al�)�]���w5�s����B"�T%�<�Q<W;�M�7�QF��z�vq�.~&���sE�!i_��Vع�'0����)a< ��RK���K�S�ݫ�=O��a���Gd���L�5���7ґM��Qorj?� y3A�V�UM��?1|����-B��KaFMW�;��<���`c��4C��;��;��v%-��j���N��ꠘ��ߖ�gD�	��J��ѿ�f��Uj~$g�ߦ�O�������� �CF��!��߼�j�/.R&[�2N�j̥r��Om31G�Y����r�k�H|����U�7n��ߛ8��5�
A�
^�;�v��<�]�OZϴ�M�E'���ͱs/,S���+~�q�/<G6����X��P !)fxt�2����5�RH2�67�i�$SK�f�����&9?U��*�v:���B��e��-�m�=ĻWl�!����iu>��7�9 Cyh+FqK�'�̊��ՙ�_�Fw/��c�t��|R����=�상��(HC��9�*��g�������(�J	��c��K�.�L��οF�k�5�k��I�#,w9�j��D[o\D���`��g�$!�0:�mh�����-'Ԡ2`���q� 2:f\��+h힖�"ͣ���bƨ*��:������_�y��?���8�%}K�5���}������TsTC�Z�'��U�N�\��;���)Q�΂gʰf�YO�������ğQ��T�0�'<������y��w�C�ޑN��v�OIus&�b
�..��U������R[�h�a��j+�Xր�sQt�c}D�Ĝ���jm�wH�P��7�V��.&����]X�i*6�z�tj���5x�~_��Nhy����a�9n�JY����|��������o�n�Ϸp���#���sA�>�l�&-ME՚�g��Ͷ�[�8�5T]�nM)�e�}�n� ��v���7N������|����R�O�}���[��;��l�C�/�j��n�<wjz��of�V��wz%z2}�kbYAZg��M��sº+��y�H�f!֭��R�(g��9gm�*`����*8;r�`�ZR[[�54~r�����������~�T2c��n�:����Ⱥ��>w:k����B����_�3�Ľ�qT�m��e�-wNv*zU��Іcz��ּ�n��zF�����(l�G��3��Ȃ`B�e�{�zI�.���RyN�xN����<+�j`�N0�ߺE���>�0�N~O��qR}?��� фed�F���(�9mn"��]�չߗST9֕��f$u$�H��ۺ��3�߶v�ZOE�uJ������\��v�"��Q���(�O��k��x�* !Дފ1eee�v�>�i�O�ު8��B��U�%��.�( �A��܎��˟���WP>P&����3A������{g>�ږ�GƏ�z�`T��$��E�t����ϴYJ���$����A�p#��V��.�n���(m�ܲ�N��Ig2K�6�^>/m%��?�p�r�*[x��"�qʄ��rA�ʋ bu0\�f�aA��>��LA��7
-�{O��� @�k����;g!U��u���^�5�RM�������Z�_��N:k��S(�X�NLB+� �Vy������-�t�fP}���[�y=�1Sr�)�5�ϐ�y����NުcŨ��@�0<z�U,�CY��2$�~��.�$'��꣆no+���lW���kM^����F��D�lG-�+N"���s�Þ+@�Ǒ��Ҧ�A��d̩J�q7�ৼ]��Gx���_�/�w����b����ʹ�#�ZԯZ��2�/iVR%���4���h�Ty��l�UuE�����M���Y4�Ť�aV���j�����F[� �.]�)t�ō�@56ɶ��F�ߓ6r�`�e۵�z��A��1sy_sU��ڵx�E@�Ѽ�s��D��K#�9�ͰG�6�^��<���c���̩D���m!_��l>�g��5���Ŵ�J�445����kf�fjH�Q1��C�D�)��󻩣$y�P����+"�6�6��~�E蓼���0���.� �T�$���+�o�ֈ�<c����Oi���,��hh�`b����t���#��|]�+��{LÙ%�x�ك9�H�	���)�.)��ô �+�mI�!Fc��/	P��^�
]R,�uh��m*�X��R�
;� M������'�d�H9�����, %�!`��)h12�pZ-`�zA$kV�H���*^�\Gq�20D���;�k�x�����F��q��D�6�B�p>����E���
u�Y%EfX�����K+S�E\C�'�Uv�6���.?n#E��W~��)����/P?���a\r�8��ӨZ����L���.Fـ�<_��Cud�%��qL�F�#p"[�ٻ�4�+&�|��W���-�����
�ȹ�!�ۅ3*�`��ߖ�m�ڕ�*�X֗�d��C��3�	��p� ��Y�%s��ܙ(}�:��H���e.���
�p�gr�������@Nmx�5����l�T"�|U~��������}]2[����T궥�&D`�`�o��s��v�����*6h������C��,�L�dC���J�ˈ�FX@���5I�2�;b7��p4����V��A��ݫ��}��;��_�ɮU��������P�%����	��ybBi�e�R����4-{��F8]X�͌~k,S��r���q{�Ck�`��� ���+�'1�_��[އ.���� ݏs�\��#<NȑRz�{�"U>ӆ��J�
�,�E0��E>̫6I���՝$i)�Pf���5e�z�=E���]���""��nS�	+�B�/��_9�Z��iq�^c���SG��ǻ�Y(�"���m�r�M�E	ǘ_;n=ʿ�u�1=%��7(tW�jMf��_�/�|�4[w�ae�/���$����{L>���1�QjK~���fӻ��M|�t��eʬ�l��q{�6�:����xF�1R7���u{����[�ᳩr!ٹ�y�,Z�$I$N�b�1���M�U�wΚR�BL��R�1hc�����Պu�"@K����dJu�=����^��ew+^�.^�s�Wk�+�ټ�xSW��M�������sU���[R��v����
QE4�}	%ƕ��dTSa�t��<m(���{��R�j�ds��cq��
PH��s��ؾ=!C�����)�ƝlF9:;�azA�s�9J�l�8�I��y]�,�(��\�%����_�y��� �ԳV��RA��φx�6�k/;���z��R:B�5I�&sfՒpt�Ezļ�+�u����lM��)����(Ij!S�G��FAe��W��]��8� ��UD��U)V�:��?L��G6.F��l�Fg�^���)�>��Z`So�0G�B��x��rO$������c�78�������p�ķ&���1�<n�<��a]N�h8��ڱ^��s��N�0��&�z��^6���4��nE@�(�S/�8�٠޺���}�m�~F�V��9daK���D���l�w`�����ʃʩrkR��Q��w&BM�;.�Å�N�������{�Z�򓫿P�N3�"$7�nR�=��"Q��&6�dF}���*��b_i�ǣ}:�@�%���Ho�@*����L�F'.���X�`������"uo/��w��N�Z�!�	�B� 0���]n�P���0�.�i�4� ��NC��m�n��dbFW��ϔ���)��=)&x58��tG�#��=�x���NJ'H���Pq�.�h=�$4&�Z�Or	.����U���c����u��_g4�t7G��t�Fgb�+#��I:=)rX�d�0gtۓ{5�߆F�0���7��B���u���z�i�V�	9�o��p�hL=ь���u���^��q�4��:�^�,|n�3%�ǒ;�H\U��2�/��
�y���@����}Q�-6��8G�-�H��i�����t���{P���������C��r7w���
��O,^se)o�7��éӣ^���yAc���Į�<]���I�5���#?e�c2�cCT���Xc1r-_S�,\e�C�w��0j5V#�pK�`��?jt��$���@��J5����|�	�u{l�*S3��s���C�!v�Ci���w�9�_�DևvL���/�pY�$����P�!p�����kږՙ q�	�.� ��,~��4_xU��ԓG�\]���WO��r�\�t*-�ժ���k���I����;.� 4��J�+�@����5��=��AY����g�� ����
�gZm�E3�ck
>,5 ��,�/w?��b���)رGR�2ͳ��s�x;>`�o��;�$U;V���SRj�! �� q�F�6P�51Q(8��|۠۾��=�:wL�k}C 1N��,D��*U����<1nD0=}�e0�_���7�	�kI�?�9�F3�'�N"��(�e��[����u���Xsa���]js�݆A��ܹN�^����ۼ�P,�3�|�ͧ�Ueo�dR��U-��^����ə���D&�ׄby���$�b���ޢ ��F�c@{�RV�w����s]����*���Q)��nQT�.�i�c	��6�Y|��L{��ʻd��4���y������Qҕ�p���L�	MӬ�����#���	��}1D������ �k	�n�ִ�f�[�a�nG|N�ҍĿ�=y����v��:C�g��J�0-"�Š ��O�M��E��U=V�����]a-�#ؘ|8��W����{�����X�,�BՒU���B$�Fx��WfŬ���T_�0_�d�� @حɤ�}p�9�O�}�h�m�h���,-`�A�	������樒o�,k!����G�【���VX����Dn�(V%� P�dwn�Ӕ�y��(|ꪼ�U�!`�̪��%s�n��='�����۾j���*�}�r�/�q�5���cp����c�����>��{Ww�) ,c[�Zg�i����W��zhS{g�B�	�r�|^��� qx�f�m ~e�KF��!�[MB\�1>�{U��+�0	�E�V�sb�.z��d��+��^�-jI�{��i�O�X��8�gr+����e�C�i�������[��j+n.D�XG�ЀŝְaQ���R�r"Ij-/�6L��h8�ʷޯ�kɟ�d���D<���ߣ}$�Q�QF�+z>�F��bv����<և��\Oɓ���z�~��VN��P�3�xW�� >]9���o�)�,���qg\�u�#0��q�V1W��~��_���#~��{���q��+���Վ�(��;�3�;Li��Ӷ�6�8!�����}��k��!�M�rx�����q�~h4r?��W�B�X/^,�jF-�`��d��pgRC^f��y����",Ce	L���t����+�seU�2����Y�r�p�I�~]
K9{�*��<�����<jx�)�����l�P���s\��oW]���{F�Gg4�x7��b�uu!�:�n�s����\O���:`�O^m�n��QOt/X+�t����Уkk�D�p�׌��O8�u��ޅ�R͵�%�s��q�B�t�	�F�V��9�4����c���T)'�;���������&�;��<3Sok���%oM�
��#��4,"+K�`ӅD�/�4���O$㰫���}"����� ߮_�|���~�xt������uX�N��^�	J�P��߅�!=�[�Q��H��G�\��g4�9E/�������ޑ��.�����M���k��dc���,���E�
6sZvf�D&P��+�EZ�`7&ԋ즐����H�s'L�@�������O�4�D}�zY~G�L���D-�գ�ˀpIMO�I{���8�|+ ��M�ȱl�7Cq��kE�|1�k/�p8cG4)DG�FƗ��	H�\b�U�y��^{�~����˧�u�99�':o�nQ%�;ɪ̇��B�;ː�]�ۧ4��l����caT�ь1��춫�4r���.��@1��2?�F�W�t�H|�@��2&u�g�ql�h&:ߑ%���@,@�f�@�*�����C���!�P���`fk������� �)yZVm�l�&^����4%���N�7�q,�e����V��M�	K:��y�0��=�������A�0�k�d=�������V�P�D��<�;���Q�(ɐB��\ܺB�u��ν��NR�l�̼cdv��K��c�5�8�&����0�Z �ɿ��2T�eW��m^�����4+n��	w����-�� hn7#-H+�_�{���vV�K-~��|7��dA��I�'�"w@��`�g��D�����-��p[,4���n2���VS�VB�)��,WH����}�k7�wD�/�h3���͑$W��~�"�ܩx��|��*ʨ�W�^�r�+�>�v���G���$��VL�o�_���ur��& �^��%h[ �5>(��aݟ�Ƿ���4}�=�C�V��7�T*Ȩ�:@�b}�A��y�]��XO`P^����,ᤴ[������Q�T�-3a�{#�;ҵGH���J`�W�����dyX��H��c��:��/��>q%:����<��Z����~72s��1����aK���21'IF1(	�����,�X������3�Յ%�������d��E�� Jߟ�F�B�q�*C��ItIO�̸m�?�բ]�؃�+�ڃ��_�lĹ�N�z���#��*�C$.� A;� ��B�]�b���*�(��e���߇r�0Y�V����C���D��ms�$I�Q�?��{z�6��n$b�6��=�r���{�p�&��^P=���6+J�!�7J�~=�y�3-����/-5�fSѻ�H�k�agD����;�jÒeM>{?��-p�Xf)��(�����1Gl�X�	�qG��r�Y�������b��2V��]���{[W�γ�=�Vu"g�ק�A?\���炲�����Nl��OG\�tՔ1�s����|8#�G��ȯ�N�y>�i��aY���)�Mc-�
�P*6��"ɸL�{�EYA�"GC�����ӡ���ۏUL�f���'ˀ�=*��� �<�_�	NC�\��0$�!��!�GG����|g�~�"�p쒫|��_]0���Cp%�ZXCJ�u���M��hw`o�n^Ҟ=ky�r�
�kww���	��d�T-d��M*�͖� 9d��y���_S�XF�aԡ�m�`�U��h }0���i|B|!h�gndB.d3վ���s�U��Gm�g5��⸅�x	�d=߃ �T�h��ST��M;8�@v��Ĭ���y0�WuYa��>A�φ��~PH%�-�}���&�R\�X�q����;#��sN���#TYy�vQ��a)\M��Ȝ�bM�Հ�jkVT�%��!9���M����=�폧�Q�Nf�s�+����?J̑k�g����}�&�%Vg�mz(~�g*��%qd	&0Amb�VQG���vw��{��
c?7��?&��?[r\�.��T_�Y~Xj�kψ�{-�qb�5˦`$KUF� 	!V��mט��o�?�(ׅ�DU{&�o;�K>�qߜ��(C�y�H뢾�WK;]=
t��	� 7����� d�V�	H�aI*��d�Q����S7��/��O�7�9����{�&��f�����t�tK�/:�����2������^�����X^��D�ti�����Ip���v>�^�l�3��c�g�s�V�C�����N_�C�C�J��d�F�7�W>Ǐ��}���?���3)*�:�e�/�X�C�A�E�gr� �>qn\n���k�$�~Ax5��n�&9i&=���l�wgse�n4�w,��$���y��f&��~'˰��uB�y%���u�j�eB>wd��I��d����e|��H��4}���P�X�t���Cmq�7&5�[`/���nm]1��<�'�j�XD5? �XX�}�.���L���^�/?��O �>XpD��L����*��{rx�8h*�)�N����pa�kF�����L���$�p�T��`6qt�[��:GKw�>�>�R���|(S
��#d%q�`H�j`���[=�,�t��lG��J![�
��6���_nP�w���{x���I�����M~�{{��	˔we�K�R��m��⼅�0/�s(7UN����PC��1��/e��'R��h,ۤ�₴h���6=��]�.>M���0;K����h3��y��|C�n�7֫��>��H��Mn��H�X�ݢWe��>��x�8.3�[V��YE��0L����n�ؑp�]����X��?�d�!�؋�*�a*�j52=�KH��+�vl�F$i���K�l?u$0k��[.ك���1�r0[�(�4�˩;�y��2��/��v(Z��=w��喹U[�s������_o�jVŗ�@%7#�흡��ɦ�jlO�I�JYz ,l���+����~H	{� ��"���/���S�1�*��/8g���,��
����F_oXD�1��o��4�f8%�hEKOʭ��a�~����'
u�a�=�M��
5�X�����\�xY.�˩E��8սe{�,�
T)��]֣��#�x�4�!���[K��CfFvmKx�>TP�+��(�?۽�;܋��grp�OX�=5Տ'j� [&H�.]l!�2�7±?�m���Ƕ0ּ����<x}�S��O�3A�4Czr�U���Qqc@z�ޙ8��~/Trb5�t1$�io!��\Y��^K�E]��J.2�*�bY�uZI���d�Ԍp��Ba���c���W�����7��a)���pB�����3m�������1!��l���F�m���Vos!q�a;m.;�߉��
)S$�V�Њ� B�WN��9|��dRu�sr�+�tO����{�鰅�T��|�f�����4:3�"����+�@��䎨�*����v����N��m��L�4�;���+��-���k����rཝ���t�����ޝs����i�r���| �<��%c����w_����`gBɕ܆��<�<��R��G�����%�����	+�R�����9\C3Z)\'}u��#�كa�$��'�sJ+=��O��F,�	1J�5�#7����T���)^�­�jC+�i�^d���o�{Q�g��K��Z�\z��Hg���6��)���KQ�6+h���]�km�i�7�Ϟ����ܛ�=O�����S���gz��U��@%:]md�:¬m�Ё;��6!�W�����ul܊��*�Dg
b�:��d�`X&�#�e�)�(<�	Շ��������g�U5׃����}�g��������3��̜��޼D�J1RtN ���;��t}D(e��>�P�;�5�\��В��^Q��8I<�A�����Qg|�y�AU���)K���nn�&.F �9��:NЍN�J��KA�Ps=�씏�B�*7�=~��+������N<���M3X�^�W��u&���CrӉ�p*���a�A,�8g+ecn��k��#ǠC�0�M0�Bnk�В.��!����)[�6�ɍ�0�~Zt:ɛ��`N�/������V �1-��/��Ow2��n6�W~��9�Q4O]o��&�;�Ə�2�![���cV}pfG�[]	��U��j�������]�	��b�z��E�M�S��5�P�eq�����P��)�H�eg������0ˉ��ŝ9	@*�
���k�'7F��`8�'�T�ڕ|�2LJ���嚰��M�u0s�s�s�`�gp'c�v��C���}KÎ�Y�S��z���_�S���(fl63C�N���n��C�mo�t�=h�]g~�&� �8��rPҀ�(����I�4Dj�l:>M�R�T�.D���S�����f�D}e��Y�U�_�E6=��_�!dJ�n��"��q���T!����y���;9,��yY�ݽ��o��[�39�������}��h^ Ix^{Pb@��>��jE5�,�H�!�.�·~����>ל�����^�@6���&�'�B�l��z��r�����,����H��H�7�\��}�
�6�S�-����Gql��"��[#]�@���կJ�w�mtx�|�3����.c���֩� �n�4��N�W��H����NDs_W67xv���|�zF*(Э���v9�ۿL�e�وY�����'��4u��l���M�<�����8��=q��q��F�Щay�=oؖ� Smp|�
'ŝ�]^s�y~��X]���t/��ʒ�|^זּ��"��B�1�e�ƕ�=��	�8ߺ�y�8DH/���h,m�c�W�mDʸ�<��C��P+
�)%��>e�t�eɰVN�gD�(?"2�v����+U:�0��B����tg�\��X?�����\w��ҳs;>�bE[GE��{<o���t�5A�:�Cب��	fOY]X(�%*�[K��IE�<��~�D<���rͭe����6�~�#�
RJ�!��ݱU��T�,Xz`��&����\W��&&}���hoպ���<�_��1�M%��u�S�=�m1��-�@� �`��9z��8=Ǜ�i	zE��KÃ3�����_>ߎ���!�k��e��3����H��D�{OJǂ���Z��mǅ���m�X�xG�^V��𤙂�r΢��,���۔ļ3�B�[��-��ȔlvW����_$�sI�j��̢�*���{���b�F�N\�#��(�I8�V�\Ȭy��km�KZ��lɣ��W��wɃ�T$�iBDGY`�=u�0b��� RH����9�ap|P��a�H�]���Mw��h�h�2p"���=����d+�S;M�Ϳ*��̇yD=����B"�U�~ t�K#�cW��j&4𚝘�;e}���4��r�jy��u���|-�)4�7k��RB<����`V�%Nt�>{�p��L	���[4 ��F�W
�GU�ҡh��D|Ps��c<�ͨĔ�c�wv�~�$�E�ndz�9Е�Q2��g6�S]�NB j��t�ϑ)͜�9�%��F&Y�Zd�̽���/�k�9�4�}�h|W����V���}
<As�Q9�H4,&�}���Lm�i���j�%����\iٽ1\�)�:�p؟qp��ꠓ3\e�����^nT_rH�ƹB���3���L� n����(R��p+��s?���ٺ	�����.�_E����2�\�ۀu��O����@�$�������D_�D[�譽j ���%4�R����?V��q��Wѫ���K�0�ӣ�8~a�n�����u�*x��+�ٛ*�`DR?o���0�أI&
DW&I�o�]�|���N�*w��2BTi�F
�$W��l�k- h́�� !G�����]�7_�����Ǖvc=FB�T��T�2Gu����������������O8�&gVe?�j)�1w0<�V��|��J�/���m_�>��堩�m(�p�0��߱�U��P�l��w����x���o�7���L��$C����K)�5ϖz���!4���`�ez�7C$e �Ǔ��]������� �Ͱ�U#�g8l�����Iz�I)��YY9��qI���9���ox��M�X�һM{��a�����Aмy�P?{��oj�(̛�>D�.U�.�&�����埵�`����u���4�"B�TP0(n�� 18.��=Wl�bDˁ�K9����G�5]E��D���F3�r���"^�����4��������q�2����e�1Ũ<֑,PJ����bzY��<��Ï̓�lNt0�k�２��bJ��`վO\���T��\����~��+��nB�׻p+�M{��Q�x�w*�I�se�ݒ�3헦I���ט����Z��X�pyX:������ �>3݁�Ϫc݂Ӥ~c��|n�.�����ne��t���_`�����e�������� ]�+�	N_%Uts�����1���Z�	&?|�!�:+�eM�2�q���	��='�n�N���3J�������X��/
qԙ@�R��s;��]?�R;�4��%vG��T]�I6]j -�H'm�t���^F�~K����#МyN�+˿
0�y�sZUE���k*��À��[]D�65wJ���=�ss�W�V��s[N�ɬ�wN-͏��p�~�?4��.}���ٰ���_|�.�Ew������8�HŌ�u�����t��ϭZs-Nn��;�b]��k1o��uoQ�H�q;����5�&reyp$�o�:$]�mP���v��{!�n²H�(�B%y]��$���B���� Y�yRqt�,!��3�s���2D��p�����U(ڞLM����9�o�^*.��"$�v�s���*):X��i ����ΩQ�-��K�ky�=���_s5��+k�/sj��Qpz"�����_�ϩն�V���=ˢ�D��y=�R �}�ΰ4v�K��@�r�m�C��b�H��NN���Yݾ ?����e�폒�V#�H����=��,h~�6Ώf�����cA�7��̙��P��acA�kl*���w/���uW�e��n�+���f,�DM�<6�{�+�_ی��TvI{�M�ʻhB �0Ÿ�����ɧ�x�0=���6*��f�2>��Rt��;9��ItE�I~~b�	y�|�!�}m�	�?AOT����|nه�;�_�������zg��lP�N���y�#�Qr����X�~)!��L �%����U�ҏ�=/�"؈�Q��vu���\j��r�BN�5Q��(�lڣ�x�'�Çv]�X�g +E>������q�ڮ��=`�"~V���o~�\:x5����mn�c�+�ӵ��[<dF��]�X_�)V.�&�b�]��^u��+����"I)�j�G�[�5��4>�J�w����6'�L �o���O��1tqđ���!f�$o�А��{|
���]�h�Z�T�a�r,�ڜ�DQ�z��D��G�%<��ٝ7(�W���ƌ�&��YS�i�d���a�G]}^���'�JA�sF��I�ˌa��Q]�f[���ds<����֔�YP�=�q������}o�1�����%5��U��_t*|g�Z��{*��a��d厳��`2���!w*6~�!���x�D�Q�W65��f�|i*Ë�����"@���l=��~Y�*f��\��q�V�,�!r`#��֬.o�1��z$1��3GT�8ց�L��ߞ�nzUeC��['v��x.DVZbi''����1�}���Cb�9�;v����q�ɢ~M�%��.���uI��߷�X4��O�K����O�DDY�s�8�:����$�uM&i����XY�l9$.Qg
���`	�# �el��#��Ŵ�]���N��j�)�-n	M*=?�L<�n�R[5Z�U/n6&ۈ�+����!ɴr�<�`�+7Ks�@��z-;=k~����c�1���E1��Y��x��K�&�����ǃc���5�[��'Ƴ�V6�ӈF��(��XRi=;��@�f�����j���LX� zd���@��#4�,�q�^���9W��|U]������kR��Kk�I���*A��!d�vV=���)�$?+�w�'k75y��cn\.�l�������#��f-|0����%9𲷖>�3��h$iV/����҃@��+-e �W�R3{�^B%���F��}!�V�?�S�����P����P]��I���YCZ�WݿR.��lپ|XxV�\��wx;R�~�_&�EV�fkF�|eR �)
���>\>B{� W2}������pٳZ��dvG�u�q~�p�XeXM�K�Mj��ᱳu8�&ν;3f_	�Ze�brxJi�{*(|�4��\wh�qpD�-�匐�1`��P�Z�
x-@��?}n{ڒ�gJ��B4׮hާc�%KK�Gk8�vm��bf���4�:
�-ు���f���#�k�jBBC�s����vz�����
�>�ą�P�.�7�+�!A�f5ۆ,ѯH���#��y��n�\�� =�htZߠg䥗@����ٮ$�-r��p��Y�sZ[n��	����p��J�fE��_0�
 |RL���q�2�3!˒�;�ҺK��x:��(���1Nu����u��H��=i�k�T�>�Z=ecU�I���cz��pz'W���~^�A�Ptq�髍s0^P���#�W��y)f��5B��償��Ȑ����� �W��̨��f�60%
[���y�Ý��Ep���b��<�����#���+.�]i$ŕ������_�KF6���DR�ş�x�^�*��u�U�q��b�KA�6��<� �X�)8���gH�}��񂐯&��w=��=L��e���|`�He&��Y}}��O@����G[�B؋߈���a2Y��m�0@�l�0�?�Z ��o��g�I�{#ܼ����өI��4��M���7rh��m>����k_���,)9��<>
u` o��2z�E�\W�ŃmO�m��@�ͨĽ�v�� كԔ�A��i�^�T�XBJ�w�̾ZJ�&��j�R�6�#�V���V�񩊛E�o�ǭv�-�$�T��Feg���A��
�F��o-��7㥷���"�CdA;�A���-�\��!{�QR���T�!d�qߌҖ�{p^�>$��$EgФ5ea�ڛ���#`s�A7����k3��c����2��d�,#��Q�ok��})B�������K���;��������0v	e��
��VY��Dj����L�S����,	��'>��:���y�a�`	�"L��$�1���au�q5)T�ah�PD#�EKL}��9�j��B�:n�OkN�"����%q�~�`�r����l�]c\?�7���ƍ�:Q���J�B�>P�b���l��/wB�Ck���Vlh}C��G�pD���r����S���g�c����s���ݏlq'A.�� � ���ᩴ��BHX{��w:}Ξ7��)�J
E�g�1�Q���w���fwE��"��m�_�*��[.,.��e�Q������J�E,���9�+Lm��(������ �苞	i�ĳ�)�����]�GJ��^G#,��,H����]pJ�kЩ��|o2��bC�����"C����e7p7L���t��%�.�Sq����ȓ6�zbn�������Q��m�%��Ѧ�#�!_vy�QI��@�3F��yѹ*�wD����b�.4�R���}�e0}S�A�Q��A������½����}u�� �r�Owh/+��H���ן5!����L�V=YEx��ˬ&@�_8%�E�4Q��$W��+1��@��kv���`�每�I|@I(4�˦;���	=��dKN`c�[���W\:@h�QQ&�T'gᬱ҄}({Q�sA��h���Y��Q[�t�@O|�1?��b��h��G�#R}Xe���~8-g���뜂��W�>|��Y��@�2�=g�����' _|�pҖ�`E*߭�L�.d"&��"�����L�.OZz,�[r�V,�>	�o[������X����OQ<a�L.6bOQ'�nYv�
�K�zՁ�����s��v����0�v��OH�, 45
m_]��f5#IB�)0��uW��a�Z�Qz�`�yVn�93I�L/����㝛N�y?}I��u�[On-�9ӝ��޹�\���\o��3���T�U/�`+�j�J�Յ�B���&����Sࠧj��Rw$��)�XHw�>��t!�[��{�˯.�}�mEJ�[����3p?7�ŝ6&�BA�ȥ߻���{Ȫ-��J�TZ:�E�C),��v,h�d����/͛�j�*n ���V;�
�3���Z�	H(�-��̓.�&Y��u�.�:��4�Q�>�9��1Dn�����%����!�hy^�(��Wc��D���XQy&)���C���(��j�N+z��)����弙�M�<���@|/�[r-I���|�x|���U(���ls@1����n>�^	h*/z�\l���|s�ݠ��=��8f�O�-L,E	A)�L��4v�G#7��a�4t�q��rY.��#��0V��H\�o�|��aB��T�}`�Y�O"�Q/@�x:��:��u.S�&�0k%;	d�Ʈ��#��_0��鸦��d�g�����(4�M��Z{S8
�N{E�.���1�>JF���A���l1
ҳ �^�:��͛�*�_Z�]�X���7݆��Hs7� ��Q��[�fR,�0�-(KiRi�H����{�
ѺN�~�A�k���`L�G�Vrå ��hhT�~y��T���>0��j����T�>���Q��X9�5-�zlg&bՀ��,�~;�v!���[T�&i9 �0cѱ�Z s�؎�X1�?[�����۸�Y�Y��r��z�@5x���������Ǭ�d��d�} RW���l��~'�(����2����U�#�z�>3u�N�~���ѽ
���I%�Q�0{���oJi�9΂T��˅���+zu6*�w��p�����n��QE�ba���8�$w���%�d��u�`��u�9�P�Y�6;[Y;�[��۲�͈��Gې���um>�ja7�����-n��y��x�s�ؼ����T���|�|ы	��꠨�?��X!�Ba������>�*��a'3�7����ܛ2\�G�o�Ch,v�-�	U����l)��z����B�iq�4�������6��,�$z9-�� 2]���|���""Q��:�y����D����3x��韵N xe�	�W�+�qb�{,��i�	�Ӌk���_�$\��8bzcf��O'�=��=������>�F'}ݔJ�6X��ޓa�[|�J�:q��n�����D+@�W6�w���u�7���Sj�&{ڝ�uN� ��0�����Gb�%մ��?��;���sKĊ2���!����p/��=�2(��S��KU�\�V�Ȅ�����J�	 �>/�S�Ӌ���9b�%�s3�ad�Ar;nz���d��ܞEw_C�������.'YxQ��ra�H�G��!D'�s(9�;Z>^���~�X1<{"���1�w0KY9a�+�	��}�f=���c �֨��?%%T��)����IA�G�o�VS��)�Ҳ;v\�~^�_��7}�J��#(�_�Y%�l1�����Y�!l
�f�u���C"M�vߔ��9yt�sjHaת?"ᚤ��n���7�&�\�S����N#@����%U���1Ʊ�v����>�!G��
��D��w����F��e�=���]B�zcPZvq��Z�2��6�c��/徵/�}�J!P0m�W$�Qp�6�t�O�xX��Ӓ�Ge�ʎ
�-�^��%6�o�'0iP��c��k��S�ٳ�V.�rƠ�6amrK��J-}�h����]O���'�:�1���,ߜ)�+��N�­�6h�-X�Ơn�*W�׃��)>�$(����Օ�_�'��l�7q�\�e��m5��_�w/H�Suo�wn1��L^4H,�n�ٛ�B&�K����J��l�R�}?\?s2�C�$0c�ɨ���.���=�U��#��w�Z�
S7�ړ7�;�-�2��DW�k��^�B���@��Aϙ`ڻ���İ�K�{B3�t�G�{�?P�}Пz���*�Xj��":G�Zc�!�O�����?� [�dyҍP�@���w[4h�%ƨT����9p�.1�1I`�d���,s�h�C2R�(���w����,�_j���GhY��3��_���)����}$����Q�����4 Q���4�ѳm�x9��Ԋ/�M�d^�S�m�="8��A��%u�ݝ(E�FCg.���d�7 _ʊPk�9�!1���%ۢT7�B^�0�بCx� ��,��ΝEZ����zQ�LbSr��S��*6����	�"�w�3urfa	 >�0��NJ��	,C���Q\�Q�����9z��F=oB.��](IȬ����T���B%z6β	.���6�*�;�$ٱ+�����i|: v(B<a�Ak�^�C�T[j2�\�;K����KK^A�w�/�������/��W����[uZc�����˰��K�h��< ����T�/�j�U��t	svw����x���d������#��c��cs7����F�����S��@�p՛�3ӫ0N���ؘ"�E2��$F����{Iז���r4u��C7�g9�3��:OtRD_p�v��{����s�Pj`�N&����`��V{����v�g�73[>!��K_x��sv�#I�*S9���.�u����;4}�	���(c�>��������5�$?��0z��h[���I�n�剡P�*�NE�Ȋ^�$X�d*l��s�y�7KN�������$��D#d෻�޴� I�+�
O���c(m��\"�(}�<������"+$o�	�QG�x�cY��ze�B6�|�Z���>��e濢[r��줜���z�GKb���-��-;eS�X�Q[�6�K�^ėVNG j\K����C|��P��˜���cO$[�����V�Wm�Rw�u=��GsV"�fs�[ʅroSO_4�۾�e-Z-�a�������솚��������	4"C�,/��i�5��dX6	s��f7��A����/���h)P���v���vnY�v�cd�Aշl������L'5n�4�=&7i^�mŻ�6��/��	D�����6L1ݗ$C�i������&*����Y�쭣����מ��M���¸?�/t;�56����4��7s漞b>l�U�/�#�A��B9��
4.X<��/��pˏf��9�	�������3UR��F���ć-��h��Ƨ�H�Ήf����e$�����'E�{zh.}����$�9���U�s	w�d(I?�
��fZ�ޭ�d��<��;N�t7=���ا�������xӮ�2��ؓ��L2�NP�����h�Q���p� �4������$��y7��̀���2C���<�gi�j�(�3��A�k�9���+���/��X�H���F���C=�q$��i�o����t�L�LC����H�3< �SF�J��ǲ�07A+?�O(	O%&?jU��p��'g��
���&�Z�h�p��H/�����y���/{�׵Ը?�HN�7�s}q����Q\�����?�9��6n��� 3��zM�&c��}�$���و������BʍF�ޜ�i��KW��j�������a�_�D3t�b���Bpi�H#����b�����&�((�2����T'������D(¬p� |4�d� �T��/��[B2������FF�������9�t��)�����\$e��T��l�&��!�RD#��z�'�u{�e->����nu��՞NE��)J��OH?�%�@Bԙ���c�x��=�2��R���&q�Q>��(�<_bt��U6�q�j��������N�H���p�I0��"�����%=!�X��^��X��[eF�TO�C�7�۵���]�Xp���I*��9�g���cޭ���|�֐��:�w�PG;��u�C]"�Չ�響]�.���0,&�WZ�; �Ԛ�6ÿ-$ 
��������[��d���$x����������;�lm�����#�"���Z�y�M�	�O��(��H�ۋ�5���9�T^T���.��8C60�ȝ=��
T���3\m���=ҥZ�-�nN��y��b�0<��%���Q���Y~@��ɖ)x��*��3�5�ԜF4x�7�!l[���`���FP���K�-d�F�A��v���0�{���n�a��+�E�#%�a��|An�|�b�,O�A��~vo(�<�����L���!$�G#���F	��H5���dy��5�����v�spg�M�C�:\^��&�N�pU��n6�Ȯ4�v����=��΁��Q9�OS:�9����r\�����<u�R,�9\*#�0J���(�^d$�&�����'���U}�r��'Q�-j͇��u�X�*DE��R�\��_�.�x��.3HN@z�X�6t�5��0�>p R9l&���}��Q�#0�6�����ݬ@�U��EP.�gsF�"�c�y��j��1KnA4�7�߬�v-��$����q�?���(_��ڜ\N�X������`�X��-��v椎7�W&�̽>ШR�ĮpsZ� � ��4����j#TZ��	~�.-�$��?�˔p?�􀓃j�{X�����k{�����F�n��XO�+v�����x�S�/*��b��B)�UX~9���s�(�9�fO��A�)�Йy��j]�����F;~��0�t��K�Y��^:�I�[�D���ҁ3���
{�O�pmg�M!"~�rP�KKσo�NZ8Dr�ܭA�g�侜��ɂ�[_ w�x>����Vő�JDm�'���H�E����	��`���I*]���ԍ%��J�y5{��!�P��z8N�ڸ��Sj4o�!�Y�qe����nY��w�y"����h/���+� �7߼
mހyЗ�#edLy�}�d�:�S%�Q�r�`���de��D��y�.|_;7�l�;�I�c�Gnl�����2x���X��B�Y'�. %a����ZTV���(.�{i�p�8�ʲ*���֊ٮ��9�:��L;�lt ���uT�v"����H�M���TZ���΄��&�'1�eV��H?ѐ_}�Qs̡�JjV���Д9;+S�Ee�.p��=�O��w��	Qj8F���5`x~[�$㨘p�`�Ob�61Y�숓�N�^l��n�7խ�'Z�����Y�(���j���/!2^ڭ�/�0,����V��җf¦%�v��lfn��y��O=�.|],ET�ɭzh��G��Yn�B[BU@�j� X��a��U�d:��P���!K&�`�!/e���x\i�v�*���4_�'��y�) �us�~�A�FڵC�� ]�9[��b?����tE?�1�-��k�[n(��������փ��X��p")&���C���1
�� �����i�?��p�b�j�}��-�<^�L%,+
V:�b�"�8�ldo:�A|�g_���C��׺M,��B��g�ʩD�:�;�P�y&������#�]��z��:#� �cI�5�����M1��J���3pKp��H��k����\l�5) Glf%˟W3*�(v����, ����}){H.�������P
0Ttc)Z��EY�װ��0.����o��,u����D�����VK�eH��@��n��)�)�ԶOb�{J	OQ�)[�4�mJ���I9R���	��ֵH�1��������������~uא'����a����h��+�IF"�N"ѺiBj���b��M ����jǰ�?8���q�oo���Ru*��fɿ�`��{�W`L�H5^;�F�5�������a�����,2u�G����'8�kQ!��+��4,X�PQ�>���뤍ϧ��ؽA��7�B'C����c�Z��v�d���+D��E��;�Y�G ���j$k|y�g����<��u��*�Z�'��D�Q��D5wh]�1;�2�hN���P��{0Ƨ����V�#EAnR۪�7� �K%���c�Xc���hs��15�~�����?!V�e|c�'�f>�?�c��!`#1��K-�_��Go���Eo��==��J���wd��H�j0g�#þ�� �>]��7�-�̓�10�$��J�����$��(�䍝�#C��_4KK����~��_w��"�W"%3&��o�~K�t�ex�a�(�E�Y�h������K�#M�cI#V>�O��C�>-!�V=�Eђg��(=:#\n&�S
�e�'��J�I��"
���r.R����Y��cýv7㬵9�,IМ+o�Xb�:���JuM�v^#�L��9x��P�iuF���<� !������B�����b�u�46V��\"+0�nm�U��>d�`���+�{�D~�|G&U� ��pr�_ ��Y�
M�Rg��m@���H�s������$�]Dv~�Y�L��HZMW��f��B#�R���P�x�  *��wDz��m�+�}��©��r�i��<Mx�>2��XhP5[R�SUͻ*��lU,�8[��� FЏ��P��xy��9��B�B�BR1G�g����1���|`*�Q��E��$W%;E�~={�ϧ9�!��G&�|���6}��έc�;�JdvbNV.�|���(�|�E~���D�� >��D������AX��eH�#��fݴ�T<&�t��r���z��RU�S'��x�Ա��m��/
�&1rFb�,.��}��2t@�O�R?��p���,ݒ��[׈�e�{��w������"A\�����@hl;¨'o�N#�m_S�'ۙ����=�ޜ���#���ى��>�l�
�XH:'�1�^��V�p:D
�Λ��Дb���0���P��u��/Q"�.H��Ka+�9��ߓ˺�90{�c�ˏ�(����2u��Vd��A �O/����R�'��9:8qGM�᝭Y�lʁ�Pz��k�G���~��$�a�-J�?�?�W�S���������L����q�Eh��w�mr����!>�77��ɂ�����&z�j��Ĺ�a�m�oW���t���{p��H��,��s/7��b�����30�$ǅ��p� �w�$�mH%�����3D�Y�o �"-�Q)�E�i7�������]��w<��5&������Q����<�iI�Ȓ�b�k�o������I�ϟ�me{���{�y�&��>�c>Rq����z�s.��4���76̈́�gZL0�b'��� J2�^��bF�	���_�(X�a[��<*�O��	e.w3��[!�hǳ�&����e��R�]�[9æ)9������O��ĭ�C��):)3"h�m��}��ͮu[��v��aK�ZS�^_��{R�ff��!o<�� AnpPE)�PL���[�3;rXtw��6�L�iw
F�+���gnL�]��U
��@�v��p�AA�H�l��~󪗤f��T���}p�I2܎�`<���<_�q5��A�sm�꾁ڬܟ�����;\�m���]qy!W5w!*��(I��v�"���*�f��z\�� >2џe���|�t%3�\n*h.�E�Em,I�4���k��II��̋U��zD �5Ð�D?a�V7�Ŷ��BC|�U=`��Q�:�@¶�	Fs�;�^Q�h�5��=SEpK�J�MJ�	b������2��< (���,����[��`�"��XҢc�w���L�g�;&Y}o�~,[᱇0�7���V[��l]����$�vKr'͑�x.$����	0"w��Y�BT�cAc_xګ��� oX�!�|��ӏ�&�����������ˬ!�͙&I���vgB�A�m�R��U!�3t^j,)�����������,�K-s�ˑ�`H0c���&~���.�h�C\#��B�ߧ�x�����j�i��j�Mw�Ask��mE�u�mG#9���'T+'���-d �&�	S��8��ykQjfK�G�_��_�B8u�N"8���O]��E9g�z����w�?`�N`rƙ�V21ڔz������i��C�K��l�����:��bL�_P���$��O(�>��R�s�ؾ����J��j���޹����%�ƒFvpw�_���ґ��g��㜮�"�[���~�4���pl'�V�ĺgyΌ__&�3��ߓ��ڣ�"qu�O�v��
yo����3|������O��ӈ���7���:u�s����%���>o�^/�������o�)������
���bQ,a��%�r�Q6A�0��_�X�QE��`�GFvq�u͆�F�9h167?�?`�$=ȏ^��k�t�-�6$����!��bD�'�|I|�N��%���v�Y�"Ց��:;l<;m�"� ���D%�Ѳ���[i;��70P�ȩ	�L/8�l�DX��@My��[:�9�~�+��G����W~�	����~YT�ڽiz��,����%��8@v����d���C텁W`���|^D8ֺ���..��,$�Y�!Y"&W܈�䒛�5/�2Wh���u�F�`	b0�B��s�
Ŭ8e@_��3:P���t́|㐱���[
�!���Jx:��su�/���E�\��d#��k
UZ�?ݥrIH�����
�T;�����em7�ݕ��hI�4׈�C�Dؙ��m�񺲤�A���az��x�����c��N�B��0o���1�U�ш�ڐ���X���j��<��{>����L�f�t� *�D�c��S���U�R��T��R\��6���bI=^Sh�N{0޲6�DW'띹\V�6���DvU�؊�!y0Y���nMg��۠�9;t��0԰��{Y+�6��%�}R5�F�
[��"Bʼ��b(��t��@�&���ms��E�� ��U�{Yt#k4��1$G���Șy"D{7F\Cm�tB_����F�YO>��}����3��c�rmE�4��2�{���y��vI0�K���
�Ƽj�"��9������6+����R������ E���޶�+sjߤm��ƭ��j�x�y0 ������s9ҥң���帆���CCIl�>����3�O}���@�X#����8�*��-�eg�,�Q�X�Q �$�a>#�x�Pze��ut�Q
d�-~�<��x;��+�a�|᧽+�ZOi�K�#���HT�l���t�u.'�����zڏ���O�����;�j���Mӄ�_,/�� {�`��T�ЀF�Z��L��O�xm�^�Xq!�����hV��j�������T�'��^#byū͢%T���?a@sNq�y:���O��9�;{(���4�x@�Q�y�ծ��b'�1|��Hߧ��q��)�8�[|��NUO&
 �.^f�E˰�/�l5��hԟ��9��{  �]�\��g�RP��$�Yz7¶?x�$�:^��W�g��%�E.�Qʤ�yӫ�X������N�J�1$K�����E6�V��o���"z@��ƧP>�u�"�z�����J��xW��Ǎm�.tԑH�z
Y�h��v����^C⡃�O[��LD�s�F��%��7��4;�N�sI���C	������y��7Q���0k�����b�Bj�����o�J�:�&��꟤IF�LyQ�_5d^�M�Ͼ[}�R}/
ƉiљHc��T&����p[aI{`�t���$���;���n�{�K?��`;�jG�o�ݏ	�	4m��?�V�����fO�vp���Q�)�Qq��� �;p�ڬYA��/,�'O�@�B&8�غ����%@g�����ݲO2�i��r ��t���mҰ������)~���a�
^��6�g��QCи��4�wf�C=;���C�P�WqB����-�Faڽ�ۉ`�!eZs���7����Is��KQ�9_��|S�ÌR�牃C~"������&'�?�Z&0*��&`p[�k�և3����ָU�>*H��H�A��X��:�.�eۖj��K�ɳB�8l�қ�]���A��0K4�9i���nTp�5��f�?,�DZ<�;.��S���^}��q��F��A.��Pg��¨�^������?im]R�.�REDV+�SY��?�p��@��!Tqē���TM�W�!Y��h0P\��0�d{�F"EpŐ�ʓ�Hh�j
�'�t��� �3r���V�zC��sb͌��RikJ��NUh�T�-����hE,:@ �A�=�J�k�U�_B}�/)*T��d�@�J�%������F|�]�+
�#S�^��k�L>Z�T�k���p����*��/%�	1�e�Rh��'���ǜ����
�m���jݞn�Y��]vB�h�����7^�!}�҈ၵ�E�VD�4>n��9�層��"�-0���su��*u#��mQ����G�����% ��~`�Vbc�f��s�׀A7&}$P.U�I?|_'��Pµ\�qh�]��L�p��)D=8P__���qΪ;آ��1�����`��Y�d���;{Έ�YC�k��4��c�Ȣ�� "qU�d�e������|��G7��&��B_Y&}��	���{V7�,�V���AX# �����!�F¹$ƍ�	$}x��&`{σဉ#�{NՌ�W54�h��0&���{��*�!੓�?���Ih����	�4ha ]؛��/~�mw���(&���Y�-���Ja��;/P�~�oO^nUQN�Ȫ�y��ڨ�u� 1W!�v�Y���� yx�A�h��f_�u���K��n���u¥�z�u��KƁ���':Vl�ꢄ�Xԋ���8m�61��j!��0��,a���E��]���.��4Ik�D���Q��.��JO�w:���%��UN�� �2��~��!��w}�����z�
4��z%דn�vJwT��8l�bx4u	�y�N�dLl��F��۔c�2� �Vp-�uK��*&TK)TI���=�z+��3���rKTM���a�Aʷ��5HR:��g��!��G�>�j�)�F�¦�%�1�OI�%���=|�Y;�ĺL�Ҕ������m�{���~��_��}��H���@�}�������9u�,9Ă�����c���Eèp��W�3�EH��Q�8ƺn+����k���Ѯ�N@`���[p�ع+cD���Q��s�G�8�#�V�t�m�-�l�U������&�)O�wj��sD~��Kk��S<n�.�m�ɩV�^�"��,�Dn�^�T7�����ZB�]m�kL�D��]��?��	�õ�٫$�)��t�E9 ���,���wu��+����r��{+C����6��q&#:����x����Ab�B	bxz	?�6��?�N(��p�Gq~��e���f.��(z�e}��k�|s.u|XB{7I (W�X�'آ|d:H��/o<a�����ٖ��?��&@��C�I�,�Ĥ��[�LTOTj1����1��`X
�>�^c�KB�� �3�.�2�����Ҽ�@o=���e�����+� �r=�����7Ū��r�1��	�hÈ�G�7���Vfy��W��X�U3ck qi�Kd.�Gv�n�{�n)��^��HM9����/�sdO
�$	 {Nv�_�X�z�ed��
GZ|�d����[��Ty���C�C*��:󲽙V��RfQى�̈���&:ou�MF]'���ZK���u;F�Fi?Z���/���ڥ������l��3P����1�̭�ۖX'gI~��d�o7�N�3����T-e�8���Qn��&S���;E��s0��0Yh~�����H
����]pb�I�^j
�40���]yʊ��4,pj�����#��z�{��C�qCH�J�����G�{�]��U1���-Ͽ˝�k�l]D�������aV����p�X��d�c+qt ��ħ��{��*UA,��D9�h�n��smE?�<�D�}�)�"t���R�Ґ�Gވӈ�-pOVQ��a>�b�%Ȉ=�W�_��*��3?�n��%S]�ml���S�9�y��
��fʁ9��/ft��r�l@ �{s�f����p��q����I� p�ML� �rgn���su4+��� {�qj���4�89?��6.@QW�!��[g����Mp�K"�2la�H;��n���w�����=]y������KT)��Bկ�[���.	�A:���,���%Px������F����h��P]���kA��ړʓ��غ�t&��[���0mŧL���\yϣ#�X*������Ve ���:�[�?(	��AA�ǙU%�(��-�ܙs��9�Ɋ?�8��M����s�����gx����=v��_~�)�p����Xx���gۭ�n�)����u���N�Q&k4�m���-������l�k�J�	;���P�,Uj�cq�������Q�e����z<���	\=
���l�5 h�.(߸i���D��t�7�ԥ'� �$�>*�w�2[�d�y<.���y,T�}]̟��SHJ�~���>���9D�pآ��Y3g��e��������Y��x|v`.����%v9�X��B��<��H�hc�S8��j�B�k����!�Cp���l6gnrB��V��^H&p�ST\z��Q�˰d�kĽ��&�ϰ�~� ,�0uc��K��<�����w�W�Y����~[A�L�v�Cv��X"�_��H����o�c:'T�G��q�*�|����B'��J�U�&���RB0)p �s����$��\뗸y�5qI�j3��Ք�	���U�d��qZ(����w�Rg�q�dwN�f�G�WL���~�s�x���.e�d��a&�N9�A����!�����C���X�R����+ZUr�}R������B�uL׀Rd�gF �-�j���Nn�����Jb{�ˡ�N�r&O��)U��Ī�j�m�����jhǸ݃��ցd3N�aN�z�:���̆��ɭ�O���5o~��,�
Qrsx�]>��mn*ہr�as4d�O��V��A�nWXo�*:��vU݃-����#(*�9.����x�����+f�V��l�8����+���7���v!z����ͳ����#��9�,�G0�Ƚ���jf���%�m[c�]�_���T~�$o-A������..ɡt�8�%d� �0��l�z�(1��Ø�e��x�����v?z�I�,����G6{��"M�a��$F{��F��n��"#9��g2�
������������O�$���U�x�l�
d<b_f��+`�4A�%�2>�a��j��[4 ���q�re��I>W����Y0�lDDi@]	��9<����5��&��)"f-h��!l��3_�>q�)�띧-�|�]ۃ�\f��Cb��G�������B�͟��-m��9� �b3[��KL���fF-1�w������+Ԍd�������t8ʓPf�U�n��f���M$�Q�Ls%�'!�0W1�=���W��bA�Ơ�%��ޏ�s>_��Q�ʋ���Y��W�=΀G�E���g��{��r5:o-��|v#�>8�f�ƒ���@r-�5	׭������yǘ]C� l|<jWף1������[]SCTv�l�^X홳 ���x�$rv:nI�����H�MHƜ�](�$O>��/J���U�`{jC�]�f��L����8}���%���Ґ�&��_�k�E�B�l�;#��JQ�E=����k򂊺�ؗ�y��e�/F!��:���<5௕&��i~���c�|��NB\���L��o��SJl٘g���IZ�ף����R��	f��y��_�;ܱX
�9�Y'��Cn_��)�S�^�R�_@����,����/�$>WN+����嚁�a�~*�'���UX���g-~M�n��b���f���
"ʑk���K�x���(Q �e�� ��3�=�P$՟A�Aμ�:�?�$`�/��ϟk � l3�d�We��#��@�f�s�&QnN��[�}�o�#Y������ej��	vtt~�:���X����1����qmX3�񵯺���P��'GJf(~����8C�=?bDS����J�sc��L������B]>����(����>��Su���mj��$��s2[�:4.��2�AA����+�ZzKDD����`�G�'�1�b�_�:�Q�I�����:��Ny���ұ6Y�k��juOY��L��j4�I�>��a�;jEf,�עy	,�����߬��v���;�3���R1M=9f��6��u�W�j���8�v�eUS������X;��Q��5\i�y��bJ�����43�����۝WH�l{C���BZ�К7ƹI?�]���YU�L��NV6�	<?h�� >7	l��SZ����H-SO�,!Aj����=��;�2a�'�,dDHYk1���D��M�N%���g�cG�ԓ�2�ʏ�Ǔ��$�KY]4���+�\�./XU��k���1(d�	}h��'I��>�<�3�$Ȧ&�l�͕r��Ѽ��<�q-��u�MR�_�q.�U�z��<K��[F��8��sN����(��6���3:���pwV��PY)�N�-�NU^ ;��AS�	�������Ƕ9�)%�D��/H'!��<z�����ڐ�V*P$����Hd�͡��Q��U�@��"2�L�&^��0J����Q�#`gzf�kw-��D���g�_���DDG4��Kd�xk���{vW�}T��M��K�����U�$�?��0�������Hr2F)�]m�zQ�h�aS���H�u�� �Z�'N�A���|St�!]��&�*o�ıD�2*<�����`r�v6ܡ�ށ���b$ۗ�)�}v�j�:�UЅ��0��^�E:h�l,��X�Rn�� �U[scNlBGV^�f���K�S��GQ3{ �?��v?Z��2�F����=^��p)�^^xҮ�A�"D�5��e!��ߋ���@!S��S�2m�ҝS��8�*�2�prX7�a�	P�Hd��a�cKH���Z������j���	��.K�*Y����En�2�1.�$�'$���,�܀�(&�@C�a���[*���[�����k?�_ς�+��N��\W@��SX���UP웣����#;��P�br1��yh�yu��`�&�3KvSjݎt~�؄����ԟ$���v��k�f�0�*�c[�
�O�ZOة���� }Yk�] ��F�m��ݙga�7&N���&yv��� S\��z@㥂�T? DëM���S��w�g�������eٓ� :�K�Y�t�E�JM��qQ��Vz�W��M;[�|5��i�P���\r�c�E%�W�#l�<�)r������\�n��/���}��^�N%�>�m��$f��ύ�s���4%N#4�����8?��P���4�wS��@���&V�p�!_�ŕƶn��)���$ZK�ň�Y�:����.����?P)W��cx��)��G���z�X�*�si+$�Ю����Өy��b���8�1j��z���s&�)��>��>��	����7�\� g���Yp¤�_]G��`��`n�w��p�hyeo�&ĵ5�*W��{�9��H�tk��R��uN�,��ҿS.T������&
(MTw��~ZŇ���;]��nb�p���&��/qBl.���bh���d� hG���	�`R¿�y�ѡ�ڶGA �.�i�R�8�[m� ��8@��Q����
�8pƑ�������C�X������Caӊ��l��_j�������3ز��]��t>?��������ͱaeM#	m�%^C_k��b��T5�,�+��RM}��.@ �F��s�ؑCr�4@zEt�8J�MX�voO[|�k��5�� ���x�������� �����v�~F��9d�%��E�פ�D�t����"���R��K�9�]���[j���o��Y7/L���{{)��O�/QA\d�~�_#��)6~6/{�7�R�Ɲ��E��^%i�zb�x�"a��HW����@�qڛ��ա}9�$�� \���$�
��u��H���M|"�r�F)��s_;%���n�F!��	LT��p������g�7=�7 m��v(
&�U�#���bL�fޮ����s!Z��*]5�m���D��3���K�ڿ�N s�y@����9��p��ϺÞ��cE�ɪ ���O�6~Q�f���qМvW����d��2����_����;U���	*��
d:��a��>���l 	wp8	�<1^��f)}փlܐnֹ�K�j9��U6��(Tlo)+Y�����`���iv��1�<��HW�~�ۃ��=~h+%�ܝ3|�;b����\7/N�B"FO����G>}�!��d�Vec
�EPH���.�xYZ���2���BzY�XY�*Q>��	A����N��i�l��.�o�KC`���K
�?��d����i�����3�]n����v�����S�o��Mk����� c�4�����В;���5� ]��2}X��!�\��.�&�ë_��.U��'�E|6���ϣ�.;���Z`�0��>=iȥLи��]B��_�kvPT,1ڶi�R�O:]��3��:U@�"�:�!���'Lg0�ken�tqf?���2)'�u8_oV��Q��cad��0P��g�mX]�w���Ǒ��G�
]�q�\�*�N_'�/�����,w�6.ԧk��Pr�v�1U����T�?%��gV9?̸�"����}Ή�⚣r�S[���Z��t�.�T����/��n�����SOgr�d��H�)���	�tGPK�O�{.B���	�`�k���9B���	T�+I��50[
3��B���|��3�^-}����I=�2G�C|up&�	x ҝ%A��?�q��*W�J=�#{4� [~2 93�FX�A��V�IA/9%* 0Zܤ��B��hU�jV��&�c��#�c2��d�G���Xeqe�)�|���ė��|��_��`�z��j��19�q�i���p2��^��F	ה�����uCS�F̢���ו�-��nc���n�*���;�A�g0��Z�7����}�����P�V%�7*)W�BQ6�@=�ĕ��۠�4c�j$��ov�C���d�4۩J�d\��q뇜hjv��|��2R�C�R\y��!q��I�Ip�/ԶH��Y���K*E﫝�G�eJ���)b�Nb�'g$�	l�XN��@�� �` Nc��g��U�:��%i�H_��F��h
�����I��+x���H'��(��O/*O��bT�!�oK5�_
8�R�|�'P:l��[���r��C�b���z�M#%�&_$ ���mz�\(���������]6�a���`pM9�! 8�ާ]P?�>�|ͦ�wr��aD��T��v�9
o��Z�B�H&�}5QF),JN�dI:f<޵_�|�v��Kg$=�L�p���p�Rq�CY�gnټ��!eDS|�J���|��?%l�Q7����"BJ���֭�٪�U��j�5�E�7��坳�D���B�ur�6��ff����2ζ[q�N� '��2��"q�H=�?BZ��@�兗3�z�@*�[��U>��<{�wn1PY�:<��чa�"uܣ�^Q�T�л�@�n��2O�A����/�/�~���.�Tտ|�W�퓇��D��?����b�Y��!#�)��\6�3o�~VAA�s�i�M%��=����e�lȪ���.AGP�;hٚm[^�@���aM ̄I,�����E��(l��؞�@�㗐�\�!/����p�ֵ����g�
��;&k��C�k/@�s%������� �/V��|�@�Ӌ�}Ŏfb�92���+/�:��^o���̓n��ɐ��lP�����*����s�������U�-m�o����Z�'�{6��r6Z����4��(�i�/��R��L�Ɠ�٘2��fE6�~�T��{}77d�+�_@@�{���LRzg�[Ra��<�qY�.�giV���GQ���h��U��K�@5��9�F�E�@��>���ՆK����SCB�!A�&܂�߿���J���	��%�e>��X��U���y����2 �rf�*�.�t{Y�rN��cYQBׯ�[����릠I��"a�]���k3`n5<0+����fh�����)]�ؤ�+�����w���x.�G��E�6��0z�&F��jt��Ћ�D�k*�f�R��_������G��] �N��ѮP+�8����uZɫ�=%/F$Q���kk. ���8���LQif���Tl��һ}ү�\Wt�f�"���!S+�t�Jw��o��I*!_��2J��@D��0�u��y��ͨ&x���\���.Ƌ���Q��E|fN�j_q��	EOC�y���:˺F����_2r��"���ʙ<c�4�n�1+�s�R&���{�|�C�&(T��LW�}D3� � �
�����C��a�P��݄G���(j���5`�³�^��gn��')Il�F],�0���VZc�Z0sFr UV���,Z�z{/֬8�ke�L����>n�X]��i�U<*R��5CY#E�[ O�2�$�0��Fm�2����9JPU���'8����7Z��r�wt3��$>��Q����wv��x$߮�Dj	�r��e��;P���9I�sՔS��0��$�O}��<0-w�\ΊIG���C`��&U��D]�2�0]�S�����m=��t�η����{f�y~�����^T��C�W���0�6݇��H\^��Y����ǡ�o[���
�������_o�L	�:��U&i���O5R�Fī��j֜�@ɍ�:eghQ�Km�@�B�"��FL���$k֚�,�)[e�O��=	o��A>���=�Dq�w��a����_�)C{2ѻ�)���6vJ���]���b����=I�Z�?��1����S��H����-�vLغ�,�k��vf�=��R@f�n�����a�u���D��&eY9���{�3��)ʒΚ�,l����m��	t�h���@u�W-��5˓�ǚ[��B��'_=6#���1�®`UnE�2;opG�Yc϶�H�ţ�W���vm��7������`p��>�=X'�Pd߻t�h���6�do��b#\-�Ak�~�f'��ИSxU]�/�B�Q=��)�A���p;��ը[Bbo�i�������4e�ݸ
-��$^�:�#/��х{0�j��8Ũ�<P��?��@�r��nDz[yKk�o�6 i�x�/��SU����x����x�@�A"��,�1�;K�L�_�|}U��!�w_m�G���\�m�<�U�� "�i]v�'�����m��l�2ϣ7g5���.c绌��cJ��7p����W��q����^�� 0�V������@�P%�S�$m0��_��՞mg����Ə2'�+E�Ÿf�^��i��5�iڵo�~BK!�F)�C��R�ݦ�J]��q���g3���H�uY�nB����3�&��%�o 3e�Β/���\u�"�M ����!X_�r�������p�U����՗�&�DF�+j�b���&�ΊH z��,f�\Q^:�X�A#���0��D��⫟�=J
�c�{ ��GX��c�P�԰!�g0��i�zA�o�����+�wĊA�K��n�6wD_�'�u���Zck�@9�v,�GH��&>�K�sd��b�q��������L�t����#)���mp�'n�?�H��	�]���ir��*�eݪ��I��{_#�Lʧ8qd�c]!3��گbF�m[�#�Ҳ�>��e�l#�[
x��\zj%&e���*��|�����3�xE���6����b/;�g��"�Qq>û/$%U��]���H����60�{Q?�Qj�K�W��m[,>���g$wJX���2��Q�2��Ql0�?V|A>[<�u6��&�ff&��;��^��Y탎!�70���UIo���L��`�!��p%\N��GRU���\�������4)�� �;�+���#��օd	�9V̆���
5�eD�����,3$���o~�.�|�?�I����~L��/��VK�6t%\�T;Y{�BQF�#C���*%?JO�����$L=�@��'��5|�A-��e�߉I=��`�y!t����ԥj�����S�8�El�����N#I��T�ǟ��H�8&�OKӆW8���y�E����j�*�b��'v�9��KI�M��)u9���<)A� �緹o�����iTl)/����(�!�+d�U� "�c�b�Ic�s�#�h��@��q��� �t�Y$��T��p�e��l���O�&����k��M�6������BQ���T��+M�7�\���n?���$��|�
S��#�`1`.�C�hy�D��5���:���}�S]l���R��c�%_��⠲���ъ��54�kR�e$�\+hI��%K�24����7���e� S\(���`�I��z5��u��Wj���qF���|��;h�ֱ���8�|��^���nN	IM���#�a�a�]�o�9nP�Mӗ�UƤrR��_V�K�O\���4�/E;��
�����u4}�5iN�02À�I]��x>��B-P��9�7*Ѽ>-q�=��~4��%f�낚º�ǃ����ZO��_K�S*��f�+���λN��_�)�AOJ�b�����?��l���M	�g�&0��[f�F&�9�ϔ��9n��q� &�����8����W����c��>P�}مJ���Ƀ�SQ:�&:�~��7��h�s��)�H����� �Zm'7��n{�鼬^e�8�׫h�u<����k&�W�ɿ��B�Ϩ�7f��(��� {,.��;NJ�PN�mgo�1��o(j�m��Ռ�ܮ�����k�.�G_���ad�0�XW��\"zX��T;�Z�'�a�l��/2��!�s�� >�M��5�)��P� �%�!�(�rڔRwE��Xǥ�O�o�����fx
l��ފO>{�OsC�ق�c�+�N8�?=K!~�7�j��o���jw�ǌ�5k�6���d^i�-�,A^~N����~���j�WE����յ}���
aR�0a�ƶM2O�č�w�whoʠa��z�X��~���!��%u��j��F����˖i1T%"�b �����l��J��H�BZ�bj�f��j�L�8/R�q�i��������d�gN�}�
C>�<�'��K/���g}��2�S&^�ђnt�\�pɂ�]��rɐ�6	D�\#�=��#��P�~`e�u�ؒ�;p��:���<��-��z�hu�:8M i�.��U��������g)�1�MT�����^`�B�7����;H#��(�]K�%��S9�DFP���	��������W���r!��<�ݍ�B��D6�Oɐ~6��#����S7>�f��՚#�8�)gD�w��a<�G\��U��+CTz��!r��X��_<>%���ub��"��v��>8��ڱt��d˪�y�/��]�h�.j���>-����Syp�4���Ke��T��ം9�/?�CL"z�V����Z0'�Mm.v� <�	)x�J�s��	vZ?O��&B%v��ȼ���#�L}k�H��:����r�[��?Y,�� �{�OF�������P36iqPr�Jv��"��N#���F��Ys�vׯxj��)*A��cF7���y�Kv�NK^'���=@��Rzߩ����#�^����W�8ApǮ\��s�|Ku�<]�L�9�f �c���J�p�'7`e���4%f�n�4�`�;8�ջ����b�pҒ;���RE��?^��������A鍂�#��"G�|���mD˵����0J�U#�H�G)�v�^/�0A�ˎ�ü�e�]�G7cx���P
5�"*P"��1���K��,�6�V���<��D����P��,�� �t�Y��#%d�bi����L[��耧�D\��Í��$�Hv~��o�����>B+��~!��0�:Fx)��KSm�cj�mF��A(IX�)p�K��$=��J�sp�gF�tMjo��� �4���wwg#��"H,��W<�3��o�rI&�W�E�:��Uwo�g�>�~!�RUD��G��D��V�5�\�N^-Y?��J�r.�e��)L�&��#�]N���c���[�O"����@u�lE���Fr.\�F��,a[�k��Q-��GJ����y�e"�sl����Ş���,OQ֊��S��.��K�k԰mi�D'��������r����0EA��m�C����8kj[�������m�g7�F{$q��\��o&���y�����E�lL�Ss8�����^� �J������?B�ݝ6Tߘ#�&z��~,g�J���a��䡽c�(�0�v�'�'��
�S#�����n:�+�n�$�L��W[�@��|͚-~�i(�6݄I���w_��iUXt��T��G|�}��� <j:a���?��k�f$��þ�W\��O�8���n�;����8�t�!b�yhL�;�'�4���/4r<��[����#P����C�9'/���b�D���S^ϡ�3�6k�ZS;
*.j1l�ZG��	�� �kN>e���AIl��B���Μ��� �,Z�xe�Y�L�J*� 0�8e�ʥ4^Ҁ?����	.�i�	96�H���P��f�r''u{�X� 0<���Z�0�i\���\��������>s)�j?E#�e��Ҍ�EH�J��#G߳�zI{��rp���"$�F �>X]HK��͞C��d��d���V��0�~�8��%ā�'�x(���8#��Nv;��P_'�C�����o(!X���L�u�j�ׇ<�~u�|�Q7��@��Xs�_�� Z=Y99b�1F�M��8�`ɕ�-d9AjPk�&�f��E��]�= �����e�ȧ=�M���>��)����m��9�#$<��'�@A��s"�@|�Um���/��ꀖ�fu"�Q�ˮQ#�\[�{���CN�'�d���0�il_ɰ�Cp8\k������F�+$�4�J���;Y o�OpS�Ȱ���[�ULI�J��JL�]�1�!�9���2��#�������?�����M!���&����`��r�`��9(��$N��''eX9[V9���N*��O0�=�K�ؖ]�澂!8�R�&vd��"g����z�}0�<�x@�֬S �>�-D�N��I�M��ȯJ�:=�DJFˏx�����\Sc�D�QA܌�G��"��C*�^��QEt��}Y���+�k�{�"����r�:d�Vڲh�6n	N��2�s��'k���^��P�:]��(�3-�����w=T�0��W�D8<q�`�
o������:9�@5��r$���p�w�m *�����Tf��T�5H6����ho|d���3&w�g�HTНj�T���a�l��GD&ң��]r�@�������:�R�����u9.>�u�Q�5z��J@�����B��]óoe �K/�;`��X��P���h��ayי�K�M`D{�i'��Z�ט��f4� � ��@R�1�#�U�s������J�x$� E�?�����!p���2ݞ[F�G�v*W -'[��y%,�R�DT=u����y����[�iX��D��z�e����;=������Q�g�H��!�+�ţ���C��xU����Q���o��dӂ�(�=p��}�Z���k	>,��w D�i��]e7��b<7�f��\��]Ax��[)$)�D�?�� cA���[���R+T���\p�E*�,{�
"��ʃ1�����4'�^S�WC%j�Ʊ�3H��"�ֿϦ�����b�[�H����o>� ���e7}�הJ��y*#Z�Sb"�~c�����=(����%4	H�&��^�"m'�<#�JW�xN��kH� ��{���Ը�j��p��wV�xx�Y��s�>1�\��7����_�]�jH���������"��b3��jW��ha��LN��`'yfp�$ַ�3�kCk�A%\�ǹ��<���d�]cia��"S?��I�'(�q��ψ��e��R��猥��K�Ky|�M®� v�ce\��o�wm2'����=I��+$`��dD�~QVb�Mg�ܿ��Lk-e=�a��uA�~/kj�<
ŰH�_)��	-*V5�UQ��k9b�A����r�\/��᛭���r��)�	8�Z�Z��!�&KG��B�� ���nl1��.b��x`�9���*�^�����;Á���r�������t_��Dk׸��7�.Vm0��y�qH��oC�#�)t9�r���@�"�A�)��n���ua�vO�٘��{�u�Km~�7Jt�r���9]���]��*	�5��l�vR	t�qWq��4+��
��u�W]Pe�l�'��d�������A/� JwzUx=�_�v��R�c^�X�2��يz@�o7�L��2�������N�+b_Š:f��_�&��E�I�,�I���q�o0�g�w���]4�.�2�q�fN�v�{�'e퇱��ʶ��/Y��X�`��|N;������'7�!�o������)?j�� �쭨�a���u��$۞z�H4�'��J�(�nh�{���~�o,�3r��[L��>Wm�I���K{s	c����H>?�*�N$�m�;�}�q&俞��ނ{c�L�#n��!V�J�Xfe2�����f�D�C�'�n<.+�R�ܡ\W��rY���RF��e�x�zJ��p��`� ����[��5b�l<�e%�܄(8�.�!��;.��|�K�9�(So���rJtM�z�ȣ��9�u4P0�q"6,P��w����o}����g@��q��7.L*PB;0�-��2ͯ��F�(/ �M�����U�'Ϫf.Q GRmD�Unf��q�f+���:0�`��>cd��^$ �%qskg�?`���������.�!]r�{����4���|��|�%�� U�puvN�˾ؘ����+�&��:��=�W�;�l�Cl�v�(�s�����u��"� 0�7���N;�O�!^���S�,��"^4���g��`��=@�u	<�q�S�&�$�v�qR҂(�Y��^洌�����o���=`kI듘aO�F����YpK�LQ�����PA(Y��-��	B�0e�{Y�,�(��=A�(�L��@�]1��̜�"B���7��I�^��2A���RO'p��&
��@/��2n��n�z�wQ�J�L�87��"�SV�[�Yg�4	ϙ�cgw����������y�'��N�l�VL�ר��9g"o;���\ﾞ_��׺B���[��r��xb�����=�Ra'���$�/E����Q#��i��*Q��`}�J�Ό�)�{������p���+��T���{�;��yüs��A"��|��L����Ā�X�Zzb8���G/xzJ��s@�D8����|ν��g`��"8���v��ʴ{�JY���+����r��5��C"%w���"�ؿSs�sWd�ĬA`qh]���7^������p��J��&��\����'}[��2;�Ei�2[k��g%�:t��v]'<|�-���
o;�\F���j���������qݸVۣp}~<�/H�^�xZ,Gu]��@��wU�����uo�v ߅7��rg��c�[�*�Na+Gh��X[R�r����oÄR�ޮ1G��;R��!�p�(���qF�3Y��5j�_,�eF���e�l�A�>��M�0��U'9�h������/ן��d��ҝ�H�H���
W��b\��e���ş1�����������`�&)�G^���&&^�v�z�m ��GS��HA�d�ԝ���Vq��W
�ְ�?��H/�W:�lG׍�Z:bL��g�e7�Z�$ڥ��-hI�(��J�~ٺ�a<Y7�~��ǳ�~W,K�aɆH�2蠜�
�9����6�p��M#<�;i�$|$�� sq��%ᡠ��j!�W��	�+��ȥK�E�]V�.��-���	�[�H��S�տ�ow���ׂj%��^��1��fD �w3f���恴��,I�C�԰Y���6P�h8���6��:j:��J�５���>��d��:l	�б��F��iR1���ɦ��4UĤ�a���y�LYĬ��S�Lt�],����.��z���j��ًN	b��j��Z���Zigr��v���
5��uC�i����B�H��}��:�(7عd��e�JZ��E���,'�Ǣ���G6����&�T� @)𣧙9���1C�?�<M�%���,�Y�������t�Ȥ�<@�RM�8��ZS�U�B�I0'6�B�>9^.v�H�t�r�t�_�b��J���K���n��^ne��A� ={���ʂ=�{��8F��70�ɗ ��դY��k�x�A�^?��}y���qvŁg���9}�5|����b���7�T/cB_�8?���R��T>�V��ȎG� t�y5Cu����H��Mg�Œ�]~(���K	���C�����`n�8!4��+�������q?���@\��Qf&0lތfth�i�������HU�:�3�V�R���߲bl�R�^-D��kZL��ߘ�.��x�>�h��,�W�E�Y�䨍����0-�m��{�
�(�m��{֛�m�4�k�Gm�p_��`�}`tt�My� �a�o���%���.��>j��Ww{��׋o~�X-�}�ܙץ���,��OI��I�� V�L��ķ����0\�-�<�3�Gi�4�8�L����ܕ�� ۯ����j���$������Sl@�"�[l�
���pH����Mv�8wm[ڐ1�Ft�����Q��h�,/ytl>�%BL>�����ϴ q>Pu�c�5��=\h3jHq��$[1` 9�A�7?NJ~�+M#���2t`.�3�j��4]L,7J��0��ȭ٩fHٸG�����	�Ӯ{�-�Ǫrh���6a�ܼ�y�!lb���R+
���%31S~��@���+�o`���	z �[�4<��@��V��v��xi�w��#v�<�5�qKP�9���$�������ó�zF{OU�LQ�RƯ-1�-�z1d�6�1��P��U��	1BV�ލ��4����ƭ-���M���}��n�J+�V�������J�������d!+���'�FPF��f�>lH���R��=�H�ڬ[:��Bc>��':؅ҽ�]���o^���bJ��;���]��R��v
�Yup	����e:(���($+?�\@˩2k$�~9E���0ƨ Z s��"L�x����VuO���d�'�sX��tG)�na�j��I�r�Det��[Dy@��v|.�`�Z�|G��ʆ ����2�c��1�dwo���m�~g�±��z��jo����5�[�)n��.$?����?(�@�C���4��A��8�ׂkn�xm� �~<3|��H�~��+Oe]fǀ�0� Ɣ�N�Tez�q^0�䧕/{|J�,���u,ݮ�U�`��I5W?8%�+~l;�{���Y���%d�q@;��t���M�7%VMrÎ��޺���ޝ@�/�Yխ��#"4�H��܉����6����n5�E�
��s'4]�:��>7f'3JD�DB�T!�܎�ɉ\��O��m���8P�K�?�G��ё� u�?�]r���$�s����N����+^����,���D��Y�P{�똯���0:� �n���^��M�w�)	@������}U"�Z��(���� ��)�ub�[&)�����<�C8�}���}4
����������t���%���<�=h��{�Β��.��^sCE��v������<E���`s�����0����`�fg��S�)����o������WKHQY�SQ�(���Ĕ34�tCZ�ne_������9��D󕡸��I�9Ev�Xa/D׫����.�2�#R��8YZ��Y�B]��N�!$_��2�w���1FBy2n�rmq��̾���h7���%����s���)ǭ����N=!DlU�襌�`2r�� β���'�!��<t�����Xj�G�� �r�(�0�2���@�eF!�e�+(m����O0�R�]Ղ���Q7��Z)��CQO5���Y#�N�9F^�y�&Qӭ��~��B�T��j��ϻ�v3�����8Pg5�z/5�P����z�E�E-`��ݳ��o:9�:�N���`�EQ�;CC,���g���,?�L�á�y� ۗ+�hB�ꑏ�v��mN�˨��,����;�Cj�B���4��
N��M.c!2�o��0W�-�(2�^�cG��ZWh���ң0�m�)��)����l\A��(�scy��R+�C 9bC���WC@�<��ǁd5���X�;��Q'�>F'�|�[0�J��f�m����~0��0� �� S�/;�<mٝ�S���(�>�J���6,�Am^5环(��|M+��7�2�y�{nR�3�O�2���x�tP�m�/ϸ�����k�*[���Y<�p�[dAv�H��~���J�Ǒ߰QZ"o7�*��Ҍ�I���/'Ea5W�emTo��q�<,�����I�cڗ�=�)&���}��]OU;�x�N�����7X1 >��,Jv���>>c��O`hGx8�/�I���	O}�Ҙ��"B4�Z�����~Q�ݷ��v�ӹlg��I�+�L�U^�� ��WC����.��x��E���ӥ���D�~|߲�rAH{�}� ..�]�R��Բph&n��uۈ^ I�n ^���a������wD��yl�� ��l��U!Ŕ��1�$\q�>*�[w����Ǳv Bɝ
Ȑ�ڨ�Jѭ�0��2�#���H�#� a�o6��-)t�2ғL>ӧ<���χb:D5b�h�w�� (��z�8�o�;�>C�Ō#�k���̂�
 �O�O���3�v��������ƞP����V`�e�F��ce�1������ep�\���ޚ��ஸ�}�.�G�K�R9�������	���}��%����U
hh�- M"�S��?\����+������7?�	�$��v%TKk�W`(�M� :7�fN�����W�|A3��((�{�o`��q�zsP�jfΏ���$������T�"�e#�]�4�[P���JϽ|������'ruBx4���<׋`C/G����Z�4y�lN�_�Ôo���-"=�[Rܠ'/w���lz����WX�#y���儤Zh�L:�F�S�B�@>8̗�ˢ�r����s�������7EZ�j֕Vú};v#F]j��!2+��@S�c����_���� ��v����G�4f�VH:l��1�����1_�腢(����vC�T���A�#�w���6���D.�.X��f��0�Q?�����0��JV����7�����Z6%��i!NPQ6l6�5��#�׬=�5
G�Gu�N�޵Yc�[�A`Nw^L��_�5��"��q�̧�H�;��ZB�Ԃ�!��w�
��ß5.|����9y}m|���+fa���T�	8/��Z�|��
K0�wg	e��t�U��Aw:�ͣ��5��U~����9�`�\��L�����8�w� �_|���<u\7Y����Px&obDf��	X^}�6\�+!�&�*��ю�}�L&aQ�Xr�������}��	,�:�Z���1�
���=_y��e6���o��4�7�"��i�qQX�2����A|��L����eN`��0��27��^�_yYZ�{��&���zs����%�:H�����/�(�pS�q��� j�j��߼�U)��^e��~Y�J��ObvX��e��8�i��ܬ\���ɾ�%�h==1��ԆeT�s�VuS�^���c�Kz��o�a>N���Z�����HKHP��kͱ��B���T���w~��D���^Y��O�hR=����ǱK�}��i}k�g�r�@�O<rPc���9�U,�UyT�́2lku�UЬ�w�]��휂4�ۖ��8�d���A�O�����;?�.��(o���cX�c�Uy��֓4��)z!��6�]n[�4��]s/���;��rV3�ރvC� 	觽�R�s�;-�N��~J5�$w,7`zy�l�;{��`�16<�x����nk'�1�W���-�xd�E������0}�|{=����.Pa�*����n�?�hJ9��14r�g%ǨV6�(�f$(¤0%�X�o:����U��c��@.�ꌻ�k��7m�'�5;X�'���g͔��� 	�a ��ҧ�}wuw"V�i6}�@��Rm�B��x�{��:�R��i�k��mIȬ0G2Gw�`GM�8��X�jv���',�5
�W�EO����=M�k:��5�+�oE-����22?+�u0���S��JA����H�"�Y�~���#��a�zq�����M��Ɉ�66�4�s�Q��_��H*�!Q�[���P����3@ ��*"hͭƓ��ٱ9?������5y;�	Z-��nm~�^]˗s�A����e�ʾ~U�IT�����nYhw	A�1r�W0X�J��m]S;�S)� Fn.��[@�❬�Oz0�T�q���܃k+�|���Ԩ���E����� ���Vy�U���#R���#�Ɋ��wS����r���%"ձ��i����z 8�����u�=�h��B{L`=���\i�V[E�	'}%�P0P9_��Rw����"���T��y���$
��\Q���j=p��n2�J��Ka����<��U,��7�8���=p�M��z��ˍH������.?�)�za{���o�m齹�h��ޏ�(?>�\�B�^��`�"��gx#�4�Q���wf�>�q���s�Ddu�q줫�_,��|9E@��Ս�=���;;�
��|�u�����lԟ�V���ç�V��o� 	`�Ϝ��]�4m3��#���g��6��y�08���������֩@ֳQV)�s���{ռsL�AJ�\�t��l@�\Dvjͧ�)�`&��	AC�S2Q۷P)�����l{�$�m����k1�9n��n������'�9��E�BsI�^��\I���
t-@���%/>s���&&�P��O�,�{QЫ'Ad�8<�ۤZj3e.;p*�h�c��ގST!߽��@S�7ZwS2�0CM�*M�����~�|:墬�k7NC��0H�y��lp�W/�铓aF����]�&����3�@�#�yĄdZ�4��1����ZI+V�����qAd��I+�Wd�А*�m����8�<�S�A��!�E�6�����[��!�_p;����׶��C	2�%��L�GrY���8B��e��y#���w1mg���g��2���'���օv�.����"�����3Q��U��<�J�?,h+B"�0�XN!��;���'���L�2;��++�|�d�;�-�^��z�����V�a-�m�L2��1�އ�&�����9v��6�T�P?`���*2<�¸��U&[���r�������ܲ@M�E��s��R��Ϭ?�e�q����<C���J�yܷ��`'o�j��C<:��&�ی����O�8�=���a��5]Y涩�[�O4z�ʑ��Dm9�][b��Z�5�
h��EH���[)���1X�S�li��b2�Xd�G"��[6U�������6#� �g$�ǩ����X~'v89H�"�W(�����wqɨ~Dї���4��I����f6i���� uH�fzy��yϞ��qZWD<j�t\J����Ȯ1������ӱ&�;��@ko�z�'�
6%��5{F�)W�w�7�\�^��1ա독l��0�N�h a�����7���ۧ�!��UO��*[PV�7�Ӛ�HH�|,��8@ P�CI�`�����C���9�����݊H�����sB�ȥ޲E� �Ӎ�[$T��-߉o2���{^�/{�\�B�B7���ܫl��?uFT�f�e4�;g�����JGi*>��qb�q�š��;xE�e���֤=�pN˷��d�ŵ�[ � �]{&촚�J;K�pJм�zl�����K��j�5O��~���噆�L����xQ<�|/c�
�����fx�SU'��-�C��륗�d{�.�p��@�0J$A�P�#�c������I�(8�N��Z�ʙyfp_H�+iVT��M��R`�L`c]�5�o�J�(V�v)����hL����#�<&B�j�x4
m&�R�=y/���� �|��)gG!AK.��,������#���32H3	a$<׌�D�?s3��	�ů��Sak�:3��[�����XH<��j� ����C�3��S��$2Bh��Ðw�F�
� ��QPP�vH.%Ǹ��ٚ���ˌ98�Yr��{1�p}K�x�X������3H�[\����f0P���z�*H��J�2��e���-t�&k���L�bm���U�Y��=0�{N<M�*���Ś9�قi�)�$]3����1?�,7���+��'�\+�ms�y�?�V�Us �e�s�!~�KF(�*^���� >NFf�)@�M-��U�ß>K��S����ʥs�3��<��F�u���h�(k��.��k���Y��Ʃ'T����	����+y�h��%`�bk���_M(�>N�a/7&��r�UW�?rcگ����V3��U�����\�VM��i�_*ӛd�-/5@�]� ߽�̿xH�W6�X �z�z��9z/"3��ih�m
/n�c��y��������<�𳵝�-���N4^��ai�vĹ����`�#
��;j�H����bh���������l^3��?�x�].�˜{=!���I�f3Ù�w�G$�IA��~>���#���^]���}@R�B�]�~)$G_PU=mx<��� �J�?�mm�%��Ev ��h�&	G��6WSEr���h!�O*�ކ��+v%������N۴PX������%�Tx,���U��Ks�>[�z/�aE������z�A�?K��x�����eW�׶�]]��!�R�� �T��kr�4�k���uf8$̸��L��*nB�+}��6@�ؖT��]��J���Y�q.�v���d����D����Y�8Î�0�G���ew�N���n�;�g59
����ǥI,u�[TƂ��/��2S��Di��������r�X�-qh�+y�@�\�\y�|H��㭬��T�L�@��+<�i�9�BT`7-��r�y��3#�p����/��l��� R��ڲ��d&��7�5P���Af�hp־�~��H���	���-*�-a�����=.N�u�d+|�5��g�u�F�>+�pq#�R����b�ޡ��^w�U��t��G^�����	�7�Lt�� ��*M0s�;Ȧ;(Q�6����G��{�igҞ���lW��*��;�M������ b[$�;�>9<Z�zL�!����ۚulD�������5�ж�.��������xHn[�$�Q;�%�[͐MAM�8as����)	�//����]���o��������Ԕ�4��e�'�E������o N�)���� k�òF���&�(��-�`fb�d ψ���J�&��˧�[����H٩\�?΋U(���Y���뫛th�������xCHp�	pj��9�N͹���O��G;��I���W8�υ$�#n�b����Z=�ET��B�j�`Jz�Η�ɲV�E;�s-^Η���1E���s�pp�L��g�=��?��0w�E�`�9��vdzXd5�s�Mb!2VoOԣ��#��g	Q7�|���B>�2��>!P-�O��Aݶ\�9��>y�E��*b�vc��	*���ĭ��{�����G2���H�Sٛ�rr4�M<�Hi�/���A�g@����_�5S�k�9�L	�d���x,����	���D1��կ��h���7`��ƽ�5��C�^n����"r�M�sC/P�k2����Db�YX���x�i�϶��[�IB��r�+�u���`�"�C���W�55+�LI`��\
R9�4	�Ka	_�Np�wi �X�Hx�k�M\T�.B�+������6��
�������U�0���Zb�	�܌�W_��c�x>������r�0b� ��x4����sK����m\�A�+�b�"���q��P*I�Oq��D��ӆ��Q��("��J�!֜?9�&�)��ݖ����b��O@��|����F����0E���ר�?0В�3�~h�ύp3�����'�Ȁ��%�Uu�Y�=#�T<��I<Vg�	�Ƨ�O�G�.m�� ���U�,��@|�h�2�R�D�O���Q"���-)��A��6�����r���X	���M�R6�gQ�=-�c��l`�A[����͕k���W�<�$YA��l���LR�n2���k�l~'%�������z�v֩��-�nE}���C�\���ꙎV�0��ݾC��36�q6P�Ǯx!$j�w��z2 %J�/g1B�`K�<�Ѫ�՞'�F����@�Pm���(!.���C{�ԲIL�f��葒��X�V����N̘GQsp1�)X"��^k�S��N�� ,�����M����;���J��v�ڻ�d)~�H |��|$kg4:��� �=T�N~Am��Q�vՊ�m���-��%R$��>{��4�ȣܕ�(#�ڬ0b�g��8���%�9nJ	4�Z{�;J�ΐW�4r�1��'6@�Đ��_W�d���#,2�6��PD��u"�1=�[��/�y˸ ���I��܄v�P�^�]�?������FxM����^�ƣKp ��7.Z��� �|��"{Xg������ybw%������T����J�2��𖔙Wgj�r���7�!$yq��0������(�㞥L-��1��K"�~�=�������������m�O��_fZ�-![n�Y�c�F�w�QS�	��m��g�E��n���4���/���s��#�GB��?)�X1L�`��Q�oJ�Ǻ���àDj}7������E٭I���^�Y� �<���-®6�F��m�8>1=*O�-�pޕ���L� �|�lu�(ƨ�K5lf�-y�A��V�!' �/����l�c�쾐���3q�0��K��a.ZF]�sM39�>e�����ta��Mt�,@�y�+As�Q��9���'�6~��u9,�̚9��畸�P2��F�
�޳9`�YDXDOS3؂s'�Ց$~x�Ύ
w /�"�j딦��}�����E9d�t���eZ|��Gݵ�n�5�N+�>Ī�B?����%U��HgV��[u�eC�>۞��r+4���&���-��d��;�ߏWȚa㪅e�#����B�\˪�5�>p?M�ee���D����t+oX�����t�7$��?2�"�Oת���~�gu[�� |ٳ��q����VC#��H �D����w_,�%-����J^��n>ӑ��(p��(Qx�:�E��{y՚T\̈V;z��X!�T�C�}�U.�ҍͤ���oS(����&sA�k<��sAI�)�s��ʼ��f�� �Ѕ����#�]4���쫞��K��Jm�T��{�o�N�j��ʡ8`Ux��B��'��˫[�����K�=���I%��Rl��`�ҋ6�ocW1{z�շ��?s�NN]���3�ƅ�����F���m/{>M=�,�E�î>�/�0 C�Zلs�� �f�F�8�����1�H
���uQ2�C-�g	�r��I(Q���|{
��Ӧ��������e�%�l��q�s]Y_	��uv��d�c�Aw�� ��yZ���z�'���$��v�j���s��-�5�:#6���έ��Q�}((6`���a��57(��7K�b���h%�vjV���&ǨA�r_OH�B���d��P�L�'�y�O��^B��]�bs:Ǯ@5���6[���rƶ#~�U�����/r2��`��А�wy�1[���ï�2�luF�v�f���q큻I���R�5��Nk�^�*t�QOǢ���lܐ��JnUZR�l5�S?D���Z��	6�qY�w~r�
��Xf��Z+����"���R ��)���9V�O�/���`��G(dn��	�,֝���ԩ�0Q�p3�����	��NDT^�@)$�P� <�>CD9?z
K������XbvQٕ+���5@���Iu���s޼52�5	������{�j��~08o�����^����=�q<GD]��N��L���X��)Ǖsb)t_�ڕ�K��@�I�^F�@�ܶBY�PlY�d	��%��~R�|!x�	�P��m.��(��߶�Nb�-�K��#���|�{��>���Y��}{�͛�^�5���J�z"�{c�K�v��-�L�b"�ce������������^�f3+�������5j]��ձ�%���:�(Z鵺�	���ORB\�n�+¢�c�����'��4D���7G��51�G.��Iƶ�H����u��]��l8-�9Qj����#��
���T�`h2�?�~]��ݜ� �"��<��r$�`�|�=�v��W��B܏E�f��66ߪ��l�Nfv��t����n��fz���$���Λ��tk��}�i��n^�Åm�����)x�b�׾�����T�k'���e
$ͤ��g�N�������*gPIB�(���mU/[�������h�0q���u輐��2z�!���v�C�5'��K�$?,�?Ɲ�ݍ0�0�����B���ܙ�l�=l�>.>��[�����v�^��;W�X�Wgpb�Ԟu��Tn��R-���"�'"/�)s�j��� W���]�^�?ačpf?Dٛ �O=Λh�:���4���WVm%�>Ԭ�9�nh��UG��L�db?!��n	n;/^�=�*�8fj���uV"Tb1������;���������SU}f�vM���mht�	�K��f�4R��0�TY���+qׁ�=��J_3�PB'V�NqFfB�&9;-l��7w����٪bs&���ϓ��3���X�٧�#!R,��$$H�����>lo�ju'1�]��a�(����6��P}�=���]	�A����\����}�5P���~�����yO{�w�_�}�ǀ���L.����4�٨:�Ц�t�9��\���Bb�oh���L���6'�Fg!R	��-�F�o1~��4�X��@�`�ݍ��1��n�B�m%V���Z���[�;�aH�O:T���ba<�+�����小8@}to���c��G��N�Q����Qz��ɝ�-o/'�Q�Q;j�W����а�`��a*���m01_�ny+��Ԙ$�{YY�I�-p��#Z��w:��9̽ḿ�x"�}�����N3>�S��1��"4��ݕs����p#e	0�T,ț���vY�fL�.�}�،$��ӫuh� H~_�X�6�ۘJW�CD��q��%�>�?�
�ό~2��r��'�2�&�nt��@?}S��X2;�������ۮDn��~��ɥ*Oꪡ��:W��ay;�JR*W���:#��,����_r�]=�ЂJ$Pu`wɩE��v	E��.�d�ȯ�rr\���`j��!eF���&<W�Pǡ-)�����D)1VҘ��|�UvP�6���!7�Z��^ˀ.iF&u������{�{�9;]`*.���N��F攪�(
WR�$9�%''-C%�Tg��ā��(�-�NWBK�ps�iO�F��0�"5k��G;�Tt��_��7������ȸ@&+D�W���� �>Oj�C�Ȼ�OA����9:��Im�� ?+�Tժm���;A|���0,(�ɢ4^�; �t��
6e�q�t*F{�n���r�q�Je���+/ �+D��9��n	[�9dD ﾉ�������L�+d�<���l9P6��#�;Q���*}����H��먪��L��eDe�3;��p	�ш���ػ� �@P:�ڼ��9:fɌ�KF&�V9G������#O��ŋU	���L�2������Y�ө�%�h�������p3#���5D�#��=�f�d��VD�{kh2sS���;W�|5�^�?��eܩ\#�ή�,'r��B+�q�?g�=2n[1������U��<fOG��c�>a7Ѻ6�n ��<�>$d�����e�1|Y���f-��~1L9i֖z�@�0ehٝq5�7��h�Jg[��q�#�ު�r<�� �H^X�1��#��wB��`��PX�ɫ��^�ӂ!�e���.o��}�[�ᠰ��@}k��\��?�ε~w/r�^ʏ���c�(�O۫cSd�v�3�*NU�J��y}�X[���E����/uɎfT�3?5���Cl��Hy}5avw.z��3JF���ݥ'��qGbu��k]A�A��8��P�l{��t|���l�9EN ��t ���@����7�H-���q�`0��l����:��fÑ���Ǎ��v�h����#�x,��#��C{�B�Ln	��P!��5�Z.�Hu�u�+���[_B�Qj��i<�ĆA��ٯ����a�~�%&Ï\v�yG�Gr΅��_+�|V�B��ګ��
�̇D^F��!�^"�.볧S� ��J'��T�N����v-���z!�&&�P_m�.1�4�0�Qy�8d�M�f� -�]%� ��)��9)�Q�X)|<�-p;/��o::��0 ܶ�����m�fQw�X�zS#G/o4NI��2�0�i٤B�L��qnԮ��1xr�}�MG�ZK!R�|�3wS�d|����5�db�Ud��|	� �V�Gٗ���{���Z,&]�|�<�����	���~�$�[����w���V�6:���18�0��@�����u��<o.=sY�K��DN�C]$"���J�̟����G]g��V������ה-�i��Ǵ_ˮ+���+�����!�cY�1
e6��U�VZޖ] t�����Qw����a�R����i�r���Shx�*����X�%���5�g1=}�[��1G~P�*1��|�)�]�f�_��'��Y$�Gv��pv;m��:��˸�<�1�n���6~%��k�3��E��0�ێ����t���S�taK�gW�049�Ҡ��j��/�Ź�gF>����	VpH���֤E �>�2��9,;�X���Ѱ�������+'��<�h#���['y�k�����#
�C?-�5��S,[�H����j�H�j!�cڥ	�dTٓ9����B���¥��"�Z;��(H=�'tT�ᘚ�]�K���{���5���K��m�s�܋U��a���c�t�)B���jUN����O~)w�Y�+:���'=�G��%����� MBps4�W���4o�-nOͲ8?.�lY)��>ˡ�͙�
�i̻�з$����|]�Sp¢�!�Bڅ��*���je,L��q� �:H��)d^�pz�'�[G4��/�E�8}�y%k����{zh�K��i�wk,���pl"d�x�Ѐ��l��S��WMQbv�S��8��d6����k�fUS.����v���c�lF4��W����*.�݀U &�c�ӧ���i�����R����N;0�[�3Kɾ���3=�����ᅍ`�����|��w�r������d��Q,�sË+���Yu����Uah��,ofc�!^�?<�����X���Ls���Huc���%$F��C4�?^-�韫��^=�hMp����#��f:�������l7�s�E�_��r�)���i^�	\� ����c�0:����2`��h�\S�?�R����'xTfBu��ŧ!���K�Be��]�u�5�G�i���u�����$G���T��鱞� ��'�N]�H"��V*k��:�����RBRGի��Nu�d��}N��!K�������rԤ͏��VCB}�'�j�J�	�,��Em�yx�:���"�k؁������6�q�,��w��%��<H��±�Uh����!�ZY�{�lW"+Ns�:*ː�v�J\5��� C1e?A��[�U�c3ީ��A����{�,��9rHxA�h���J-Xr5���߻1��M�Җf1�_^oxD�מ��s�Ɣz�ǌ�k�8��v^ \����)�7
�V��;Eb�]�G��(]�(醗����V�=�>12R7:��:T��&-`bq�o�lQXUo8�V�[Ő�]2	�'ʫw~� s�1Lh�N�6u�
�B��x�d؝��n������^�n�a�^oZ&�<?�_��کe�>�} a�����\��/,Ͳq�a�W�i��q�����cיt/���Z�����$'�Kzf)����L�� S9����kۨh��+޶����]Bj4�~��+��o1�����z}��`(q�t���-Zb{*��N�]E0	Z�����&����׬$vTb3/>�N`5�����V�9#c��_�����0X�Q��$������9Xӹxt��a��*)(��7-'-��zt+��"n�F]&��-)�<M��,�|��H�-����s��%��}-��Q_B�J���b�B�6����3�����E�Y�Q�#��kT���Re���_*䫡C��S٤�軀£�Ct�>.�8���%��mu�&}���"g�e�����_��. ����F ��R�镎�7̩�3f0��Os��ɖ�as=�Yd�a!��<�n�6$wX9�Ym3 kr�Ǳ�A�7f��3���ǭ�TE��$�ؼC�o��2�	�F榦���FT�5��׆Rl-ۇ������4�d�ux�4~�ڣC۫]�c��y�7�^!N���\l���^�= %W��$G���N�3T�aO��"���']>�5Ӝ1;f̎$4i�7{U��ʓ)�r@���A��	L�R�:�Oi����Xsk��#C���\�\H��,�~�Yz���`lA�w(�+��/x�rxi�6;;o�_g2�x��]4��{ ����t;m	x�3g&��W���]"�<d	ք���/����Gu�ŉE�[H�"�D�D9����(��3b_E�͉�W���� �[�n4�!̯����ԝ4Ț�f�D�����P��k���*�-�aB��s��^�4l填�^Z��!�=�ؖ�֕����Ɵ ��D�n�^�FSW5;/��`䟥�V,2��-�n�I���+�0g-y4m�����{�`s�R�t0�$�y�]�T�����5��j�����4�nO�B���f�r�2�}H��� ��d[B@����<��룓�YZ�1�9;2�.b3v���i��E�m�-�%T�$xė��w��g��7�@�4��̱ׄ�����pt'��+�8s���,} �t*zW�ųٴ~��3�!�M��#$	�I��Hh2�aY| �Γ���x��b�~��*�ϗ�J�|�ej�=@�9	k�Y J���le�j.�>��졅{�{�1cw�&��#9,bٔn9$�L��CҚ}G� c
��Z��������t�:��G���q�#|!ê�k�ރl�/?9,O&�%��I������"���3���q�wW���w�Dg?F#���a���P��G{_��Q6m����[��I!��@t���:���Y�C�/�7��H9{�ȇ�=%�%Z�L@���t%)M���(�53|:�-�#�Wύh�o��YR�᳆|���%���¬˻f��V�Q�I%' ���]���A��4��8Sexb�g���(7���������O��)��t=G��/��,���L�־:��u�!q�Ww���;��FR���:�@���<K�YA�7�(�dG�F��oK5���>u�%	(�[�u��S9;�8�Zx�}��L��Fu�'�� yG%7�1�}fU�w������>��YG�t^�6�O�`���A�Y� �4�R
�u��uf��n��D��bYK8�ۢT}�{�<���#����K+]��ox��;(:�/Z駐��'R�Ʀ�:�bC�bA�8��#�����a(k�F/]z6?��<�H��;z{6sG�Z)�_�wHb1@X"��>��(�xʙ6�R8a���W������ׅIk�O��k��Y�ŋN�^����S��WrA�ă�T�>)��fe�b���"]���Y����5kKN�M(C�ꉲNU	N�q�oUhXMBG&�u��jњ��vl�@Ye����UO�'U���U��W\��N�h��kữ��k׬?.��n�b�T��������R�`5��,�w�t�&;��Y<l<Bb�e�/��k�n�$���]ߌ��T�c���V�6���;�Y����Tn��`���K�j���L��E?�6M��u9	�`�K/����Эuͱ��fQ�#�$$N7�2����U�Q�5�h����Y�����	���PM3��O⇤���{�^[�|b��3.�׷��A׮���_�G ��z�o��������L�qE+�"(c�\��Y�g��c"LX�	��~3���Z����.�W��HH����}�vc��3.	ō��f�{�Y�m�x��L��Tq�/>ݵ��˒+G@���M|�R|�w�@�a9_�>`JP���j(^��c�Ƙ��_�EaP��0Xk\BƴOB����K�R��^޻����=�[��"�6G�IqP�r5�3�[*�T������������H}̥�٪���e3���\�b1��Iغ�I����4�+��F��']ȧ�5LI�����I�4R��B������*�=����'@�������~��=�&A�x�3s�w5=T�f�s�w�2�3�\�qzr�F~ZM�.�2�3#���OSm�J��})�����|VOq�罷����2�4���i@p5�F��{~�\�I���B��C	�W��'���Jś�w�d���m�z����1�^���k�*kf��e�qM ��U/�Lk�+��Q N������}O�R^���=7��������L8��R2 i2�Z=���O�S{�F����$�}���Rb]nܟ�.�6��l�\�8;x�϶.�2�D��]ͻ��)L�N�^���ن(�%��L�?w9g9ͯ��s�
{�w
�b��]���3屒�G���$�}�\C� �e�UTH�����V8L:;H�i$=��s���B��:��6�S�Cw�0uyը�{����>B��K���8�`�Y	��!��?�#��Q�S%�C�I��H��/b6�'���jX�Z�U�n	�w��=O9g��5Eg�E��ú�X���lc�Õ>4��x�/�A}X�[�o�qÜ�ip[�g�����"�����$�Ϥ�e�Qi�-	Ml�DǏv�Is��^1P^4��m�z"q�8�*���3�;���&4_��^��̚Ch��
�\�f����,<���|��R���\��ڛ�"�}���߇F�.z���u_3�9]1��Sk't��E�����P@bMf����Ο�	A�A_&��Q�i����XP��{�6�4���՞�s�tr�A���㝷��}`W�$��	�m��������q���f�T���Fnf��Lrb��@���f�#�� f��a(>�%�sf��;J� �,����fL�L�E��v����mY1:m�6&��䣑Վ�Ηa���mut����z��<:SR�*�y;~ׇ<[����<�T)�m1�Z�\��+�nX�%�x����8�N5)?), ���d�	��AY�'[���z�V����1�O[�5�����jD,�5>��($�с�&��}תY9�4��p#���9�k�jFn�p�����H�͔C�1|]U��[<�;��Rǭr5l�0�*�rO�i0F�U���!�He�?�DK{��<�b�&�^HnL�'ʞ����y�~�����H��4V��N���kq�mCq~\�@2��Zl`],�tsT&���":S��Q��L�E��L��:��0Ocu�K��]����L�H�m.w�#u��֝���Ã���+�8��*n��0���+����3��j5��><E���c�i���i�������K}�=��{�b��3�����J�X%�}���t4 N�0�A�8Jg�^H�|͛��	_��vm=
���ȇ+�f�^Ϥ?פ�9k{�gR�<�!�F�#���-�,��q{o��Ԋ��?Tn�6d����~i�EIy�[چ�?c�J��Vv�T��`�Ȍ�éN��+�;���IuФ �C����n._��C����y�b`�D��;��j��+����;ǽ�8��\V�QͶ�V.pn�^!�"/[���q5���j��~�Q`ݾ������N�%4�\��,��M+�|�[�_���:�0��mL���Y�bFѴG�ą�m:w���N��ir���|O
bm�*����6[�?Y
�RBm�!Z���y�l�d�ue�Yc�GZ*n�yˮ^9W/��k�O� �Y�n�gf��#����D7 N%��h��>�V�S3�0��S�&(7�추T-�-)`5U�(�3+e1��zNf�^�k�+��D���3a(<�����t��T�ϴ�pv�B�V.�^�u�R�V�"�+(��m�Ѷ)�NJ���)�pPL6��kY��e>F�|�V�ΎT��Zќ�!�g�肦F��σk|iE/t�oR�s��Ջ�d�m>c��`��<W�����B�`����v�^�BE�pT�Ք�_\	�~�m/��b��d���d^ȥ{w�������[�h[I8�\`d#��߱e�9�f*|��Rs��"2�\��A-���1���gifU�=���	�Z'��Gy}�A~�i�`�W[m˜�v�����sռK.$=�2�|О����6���t|�fZ��j++�o�`{�>���*
_�D�e���Z�r4pf̓�z�?գ��T�O�a��\,���`V��d;��-��r��i�V�ϝ�[Z3��㵎��g��z��g_HU�M��qM����XUƼ��f��}v���Gև�4�p),m�x����O��u�_"���i5Bs���&O����>�͵�*.�cj�������ŉے�ԭ�Y��H]0A&�D��^�� C@��~�?�B�E�9�	?�'����ZA���Z�����܃�R��>�U�;>~�k�ۛ"�N���~��z�9��KF�A����~�]�<_���x�d��o��~�����N[��+g��?�s�����>���y�S���T��w"�>��O#v^�N�rj��s14B<\
]�Zr����GxE/�=3�`R�?z�N�n&�����nT��R��}�z�V�
�[T�NKo�&�%�{%���Ʌ�粌5�I��b+����˻\�x�?-��/xvaE�����X�L�+�)51Q�I>5�=��a�%g���N?^SF	��:Gf'�#"�x�L,�l2Rƀk�љ�B�/��3=��v,���b�Z��|g]������d���lSU3��U�y�Ġy|������c ���!:l����.�'0)X*H�$p�B��[<�L8FDI3�c_%gm�Ӹ�t���cXD�V��[ϣ�38|�, [�d>O}�3����������V����z��ģX�ͽ3�OA�ڲ�o�2F>����D[�Ǹ�A�a���X�.;^�;�$b�'qdyŏIQE�Dx!�vٸ�-���(U�������jLE�`�Mع��=�*b�#�z�P��B��نxEsbg�O�t���S�Tb���S��j�B����֮V��G�j�IE�C�k ��9��^"��f4�/���b'��5�S>z�;2'��y�5���T��ES�#ݏ��_��W�0��"�aєƝ��F��_O@-m���-8w�e��~�XՌ�����������;\#
pg"lo����-8�	WSE�i���-�b��0��v>Z��q����о���C�<��
:��i�dA�N�Y_�c��\���)m�Ҵ���X�E�p���;?S�z�$t!����]��k�T��~�~W[�{�ˑ�-e%s�a�5H�s�'���Ģ�ݨ;u�w�}�τ�e�h�.q�,�Ԉ�W���?#��yDo�*g���|ı=�4'@k�5����X6)3��vb�_,9r��TY@V*��=��ה��u\�²*�I���A
�6<����i�(�J��VR綟�\ްK�9���1.Y7�M��&i��壠�_���2U�=����<'f9�I�W��f�V�w/�׳� [�<׀H��߅E/����&$���ET�m?�.*��w�)z>Z��qX/&�(v+.˩��N��	��wS̚���cy��NjG$�*�rL%�gU	���I����e%�a[��W>8|\dp�L���ބ��c!�(�'aopK����p@�b
�n�ka��:hM�zp����ѵdt���s^16&�KH� b��y��m��C0S��鞂�Q�����v;������=�p��4情XN�ݠ@�]������D.�C��b������^�ȓgk�Ǭ��K��<��'�Jߺ�S��TF�9j��H&)9Ԫc�)��s�
��_uE���#��:�?��QWH[�����W�̝�7����$WO3k썱�{��S=5��3�����ۘNS�����=f�-�
��T����mEF��D����>޻7Ϛ�׹�*U�*���pX��K��+�NS�J*��h���ػAϏ�9�ؽ�x4�8n=%��}��\�!2��],Z+{MQZ<mʤP,����N�����Cķ�j�D�^��ڡ�*F����)IQ�Y�ë�� )��m�/X��{��&��d���zFg����a�8�ؙ)����X�x"V8������7t�Z+c��N�zQםE���mF�`��LG��=4s�L���3I6�w�Fצ54�Ǹ�HAb�K}�z�Ǖ�`�
*��H�,�����[u�v��V�����6o2i�A]�wǫ������-�(�wUY���i�K����;�yMcr,]�� 0�Y�( ���A�ia���Ǘ9l��Ƣ�-�{u�u�b�dd�@V�-�"�Z��&q%�)����Ѓ��٘�A6���C$��,�3�:]�b��V�=ns�--��Ӗ����@��Rh��/�rk��t�� ���7ќW3x��.
+� ����Q"��F�q����ądd�}ք�G�c��J�5���eЯ��h%�!���O#�BԈI�hI/�8"�)yӰT���u4�����J�� o��"��љ'I���R�W��unu��������+mz�-�-~��T�B�(:����ҵ���<<ߩ\�&5<�;�n����g��z�MJ�2-ٗW��&8[	����n����$��]5�0��5� ��鿳�h�I�E(X�xL��Yz��R�R�ba*��A�J��Lb],�{h�Dx�g2� wQ�4��'�I**آ�I�rP�)�J��j}2���t�c�,�Vc<�ky^lȢ��ğ~�İ��$��qY��R9�i���t!��ڼ��%���&�#D��A<(�G;]ޖ�r��:�~;wv#�5la*qr8&r̸Կ��Y��b��qʜu������w7mGN3�j/g�.�����/2���(�pK��;�[����HݼT�*���w�.uh�&�"C3ᖚ�6U��D�}Y�@�eJ2a�ܡ�����͊�r��$�?�u�9)µrӹ��i�Nݽ<�t�3?(ٱe.����=(�̀������ ��Lɜ?Kz��AM*g��-��P�������7d��\c����P¶����*�[�R宭����H�@�����k�]g^mm6g��y�U�a�yw$L�ō8#)��6����PPn�O�Z��o�$Ī3�l�ӑ�ӹ�]��5�0��rJ.9.�m�um�\�D���1F
�H+�dg,	��C�6��z��^d�ɺ��$��y���PBlt9�RY�G��uD�݆bVPFe�����O����˝"^�!$��/WZZ�+��5͓���1��v���tQf}��R\��[*��l�S�)��
�
5�0m�(+�Aӂ�|�K�P}�����5C����� ��vsڙ�k���</���WZ�GB���eL�O츽{sw�Oݺ����T�- �����?[9��C����=�%�[X�[�	P!��%�k�9g�	Q���'�����h��L7�����子G'_U��a���V%��C.��	c9�Dbmz���4�/�]	"���n����:�xX`R'�E� Oa�[x�X��6�vUL�s�3��B2k J�	I$�&V�������y�%���m��w�����Xr��,(+3t}�ų���*U������lٜ>��Y�b9*!	�aF$9� 4�ym>7��L��+j����`3c��J\��@7X^�U3��j	)u=�YƫI�g8��0��	�FV=3{�G����m���>կ����#�E�B���
�gL���n?��wź�n9�E��g��]we���隖������f"$g�~�k�1eY�3ښ����s����ݲ�$Q,,�����٭���A$_�Ӕ� �(�؆�I_�Ed���T�9�]�!E��ɯ�]�&�q��P[��2NHʜBPhn�q�j��u��n��,#��b@S3橵:�֛��#�h�sl?v�~v�[ϻ������N�b0nv�Z;�=i���?�²���w� ��tF�X6z�$hV����[�
(���!� ?O$���rq���^!���L�0���=Ï��*����W�j7�hA���I �N�H�F�L�������UcxO��
0����U�y�)�I�dbn���8�����Qp�8��h�t�N���4C�|��&�o���Ϩ�gh��h������J5����m����q�$g�`!	�?�l�ل�CAp�c�T��e�5ʢX�+�����/˓���ev���X����:8)�v�m�-�`K,�T�v^����Dq������R?I^��dg �I����c��S��u"�m�*��2Þ�.���1�
�L�]ۖ�h���PH��A�YYk�!���5��~��,�у_��`g���CAҽ�/c��(m�wh��3��@���X_��yD�v�7��RXjPߡ�Ht��Lz��4�5��f8�oߨ������f��Ŷ�������j���N�b���x=[>��������Ŵ2����nJM��=-�*�{,j3 �K�w��+i}����E;�LV��̪�7(�s(��N����^3D��]Yv4����;���Ч��]R��܃�܌+��e�B���w���ԟ��e[�~�(=g�%g|rNS���B���C���[����
���I�F�@��ǁ�v�&K$�6<���U��1�����v�k��*hy����{މ�=U2'��/�y��>��Df��p�3��#��n��\i��wtL�b�P�&�SN���7�Zj�nw��������4R�<�*{�Y$��;�l�}��5%	���gt<_��"L]4*����Y�	�h#���=���%3JL�s��J�ܸ�|�ə<�,�	�����=c}-�"-J��f2�l<�r�ǔ���9*�1Yh~���\2>��������7H�=�X��c��$7�	���m�!5����_������|�U1����?1NP]�'"�	�8�XY��H�j�s�D��D�gL�	D��HB�PS�U���=��4�������k�?0�bNܧ�5d#�����W�U�?�~3�$���յ1�� ���V[I�R	�c�=TD��Fe���j�%�@5�th���w!�Ѥ���Ǆ� V����x��Y��ރ�8tC�2�X��� ���<���_2�/�Sdf!-m����z��H$*R��NB����h�����e��� �e��H������rs����0�8j��v㫯��w[�u��}��7~z�pL���<"��+��g��7C熒���VZ>��^?�7�����>�����tA����6�!�4U"iL��'&t�TM�s/Z�I�*'$bRy����Ճ��x
ϭ
���`1G�ąy��L��&i}�8�,1%vaG��#����)����n\�U��x�J��@k�.��� ��J��Я�N�ᶅ����(�ʃX���!�'y��ϻ�%X�P�|iD%�#rM���m�K��dAp#pF�[#[ҫ��!e(5D�"���wDp~�+�p:jC|_�2�?���S{B�w��rc E]�ɛ�tP��c*���f�dȻ�N��̜�8��z�T���Ow��gꆋ�9��9���E���`>�N��$o�������M���R�ۮ͂�ʼ�RS�ޯߕ�0 �9�����3Re8���p��6j�p�����Ò'Ts�3�c4k{a/k#DP�����Og�N�uNHrW���Me��|}�Ү�nIF���t�G�i�c�����+L^�x�x	��	7���f�"���:�*+i���ND��H����Lf��E��K=�� �x+|��a}V����W�tBP;x&�1�VUBg�J3����
��{�>Ӳ���]`��*��f����A�O�)��C�5��K�ü��ww{�9{ic��a����8+�N�2|�Q��S;���!z��3^� -�^6c�j��:;� [����<I����fϚ�4_�2Aۄ��!��00%Z�`PZ�N(����/���f/�zH �![��KW�F��S��U�l�8tQ��Nq���S=����ƴ_�H�#ȵ�i�񭝱d�l���;x� \ ue���&��|�TO��rÞ�����Pr��VռUP��0i����Cy���D9����2��Zg���gL�1�e�� k,����|Q�K]��|X��2ٽWwf��C�����h�X�q���洘�*�o5�cU�M�tS�ho����"R*���/j-kr!۟��ӼI�'�k�%�������w�����^�Q<�����'(E3�(���%�o"��^C�����R�����:��b��Y}m�9H_�=0t ���$���%Jz��/`);�W�
[��(�K�}y�)�=����'
���~�c�Ƽ⟚�48��2��]S'Q��W�O(�����w����f��5��ӨK��O��������X��s�՚G�x��^X'�uJ{�Q1ɷ�ݥt��W���<�����3�::��ځR�"�X��?��(Q�,��P7&*c�t�N�!rjy^;���ow�zr2c��$<�{6d�Ϋ��+]@�O@�XD�<Z�r���h�}Ѝ�<7+&�E[z.�n��#rR޼t�_����{��Do$�[ �br�:�����N���F�����\zu�d��ȼ١eh��CG@�e6�0�����'>èt��$�Ͳl�����qZ`]��ڽ���f@E
�g}K�oo��y��<���]�dw��Y/"\�
TPx, wb�!\���A��$R�cpڌlGþ��SkmK��+R0�9��;J�~�M�t{�/l�%��l_&{�]�D+���61��Rn��n((F#<C}+9'��j��ߩ�F>`��*@�7#�����d�����e����f��/��DS5� ��v�#>�������TV�����H�\/nѯ��%����)�r�*%��A ��(�v�r��"�[����Y	6���@�-��J��oΪe�H�p��)(��%MԬ��������)� ����-�p٭�50�V��^�����hr�� n�.������ƬB���<��EY2Ad�A���U4�`�
kG��j�$�����t���{����=�q�I7��',�);�@Z0;�[v�o޵T��ͨ�ѓml�?�c"w��qH��H�q7�q�8�yZ�l��DYbaj �%DR�;�q��`6 N�g�v�m-� Y����n�|+'�e����Fl�Yj�"S�*}��2R�o�5Ӎ��yC�G�E2���w���C�
Q�[k4%0 T"k1 &�EJ�`�*�*|��"�u��%�v�u^�𯻅����[?�:D�8�: ���~�p��s1��.
�)ߨ�m��d�:�SA�
�ΆO^��&$�*&�6�|ʏ�0U&��AF�ͩn[V�P�������"D��'_��R�����_`�sО�57g݅�ymj����t��?Q�ܱA�ͨ�Bn'˾�,F:�O�Pu]Gq�T.rJ^yc{So��xx�(u�k����A����d2����1-���fb�KN�hF�j���1S�{�����d��q��K! �Qyq���v�d��F�^�@ �uuҘ�/1�ٌ���ʑ��d[�>��a}H�JϺ���'�����. �pz
T|��ga|���\w�����F
��f[�ymQ�-Yu �r��[4�q+�%Ds��pό�P�J�Ըg�.8W�3���ǳ{4i�"�܆V��d�\/�+G7�MQ�Zto@�D ��d���o=���BÅ] !\'�*�#���z�b�>wm�^{Ew��Z�@0�5,��`Pg����s�����z�`9�m�7�٭�,,�5e�%��~tO&ǮR�h�vq����Z����8���u��i`���x'�{}3ѐ�= ��J3W�%#��Oy���VoD�[@I���r��v�����u�ƽ�8KK(p�@�be�&�F��L:�}A�>�C��t��o�P��o(���޿#q{C`�������P�`��+�+�v�o�����/�0�Y�'E����w�(q�Ę{�%`9^<��3B������m�k.��[�#9"eG���i���q2ƫ��bTh�L����e��W��?Z��QCA�${9+2�-t�P�NuE��1���JKn��qh:�����B���'�>D|c֜���u�7W�f�#Kk�Х%�\��u��>�m>M�s�rC�k�\	� ҟ���Mp=���Dz���> � ϕb7W<�}Ѐv:��d�E��,46<@�"� �}�wr�N��6I��IT�3A�83w���x[M!C����,�n�!�g*H����2{�L��e�TbF�hg
�bzm�0|�?_IKY�k򶔔L�Sze���em>ꕽ�y��G����ޫuU<:oB�$��IO�^]zcמ.�������Z�o`��Tf�����V�i��0^BI����Pnaz�hm$�)0���iq�xݢ�7�L��<j��'E�r*��'eV,N8�Fo�I���]�w���,�IJ���� ,:�0�5b�X(�Æ״��z)D��[{)CBmM���ن�ɮc��O�j�kӶNw5_��.�� �\�j��_1�Z��k��qL��Q����h�t̍�Vr63%_��׳�%ۮ=�� ��=�)*%k	���Z��6���(q=�7�����h����Qv�w:�:_	:v�G� ��V�,̧4%~�4l�l��@����>�Q�z���& ߹��7�ŅM�º!˛�5��Oe�����oa�K��Ԍ�|Ky��V�g�D3_��j?��y�{Ih��|Չ��s���W�q3+�\�7���,�
�tA	�u�P��~�efh������ + D�ǽ�������Cww�8Ku���.��߆�I^��������?����> �r��{v�_�j�V��M�Su��a��aݫ��fM���(�2������
w]���	P��D>~ ��yE� %�^�\�	M���
_0V���*]J��{BN.AU���fL��j�J�O�6*+��6��@g�����	��T`�VO:&U��n���+%0����B��w.M��X|���A����ri��@�m�y���&]��hp̩�3�hF]�l��1��@1;7���.��������]Nq�N�Y��a`����z$zM{�����/!(U�7�F
�}|6�;���7��"i"��6��OR���)>�Օ��|2u�9k��7 �a��yL��
m�@�J�T��� �ݦxiI�9'w5�Q ~Ю6BN�������nZ_��ս@��POh��vC����_��%/3�(�*򣄊�?�A�[��vmY\e�@cbkߌ3{�?�NjG�i�6ב/���D��)C+�c ����������k�Nݕ��[�O8�Sh��/���䞔��4�חB��$- (�TO@;�)��ˇT��J�I�E��v=��A96�c��3�5������)�p�0+r��J���z���ʋ�g��4=\�&P�h��$�*Z��t��g���0wX�LO�O��I�߫�G�w:�ѳ����ň>�.Ȑ��"4�	�9�zE�ÁE�k7��3�~�\ݫkV[�~h�����iY�	jG��Iw����ͽ6��_�MC@ؕ顰R�q�Z�����"�B�#��z('��ۿC���Y���F_�y�_X�-�s�!DU�7Z.���Y艘lwg�9L���÷y����G�x��]�/H�օ���J8҉-HB�D����d����a���ѷ��2��/���!�}ŝh�����{|���d�Kc���n��Y�����v\]U��q�:/9����l��#� �1��)
�T����<���6��b�T�xIMj���1`a�e>�1��Nl1bA�7��	�~����%���5���'��m4v9��r$5���Bۂ�<�y/G6!l���|ϵ5�I<�p�_� ��Zwp#r�W� �3a�^�!���>e�ʨ��y�C�y��P���"!`YT9�'�\�|A��{�$�[�?��)�B�w���b��fj����:��	�(|Q�HC�t��|"Y�%�O/��g�ً���
��9w�aD��:���]�fBt�
�L��S7�w? tp<*�_�GD�8��{͟�=_I�մ�f�2qN���X����#��!E�ѓ0$�Kq��jī�K�7�S/�kn:I��ߚ�|�y���`��?a���J��O��$���⶟�Э|[����}��x�<�[h�P,h���ek
-�;��|�4NGq	;���.��W��w��ܜ�C��^yMa�����p�n�-aVyJ�Z肬�]�輽ޒ�$&�j���la�|K�6"�{��.�z7�_����7|����g�aO�S�$/4��6������V^��x��l�S�(� l�q�ۤ�m~s��dΣsg��m\��%JJ�u�;?�y"�8����(ACŒ+�dx;%�]ڣ&Ì{��E�22�,7g|���z������R!2�ƃ)R�`�bL����qcpB�Q�ם�Q�"3��E�"������M���O&�F)�\��P-x�tb�m�Ӿ$HcC9ҿ�	O�g5x�X��ֆ���4W�����8	��_LX?�!��l�i�1��?��|��0���enp��Ȫ�XF�G�А�\�����fԂ�:7V
c2�P�[7�E�WL6�g;jk�Yc�����n��Z0*�|�BR�*��O�Qm�Rrt6MGD���֞�]`����5��^��i����Q����/.w8�q�����z�Š�M&�����t�q6�6eӌ�8��|^yB}� ��{@2�=UmU��f�o�S�KU���җt�B��Cut؏2�cd��WـL��*(�*z-M)���U�����b2?O��縅ƫ����u�k�9{v��TsQ@��+�!]��1�Z�B^�*8�T��|;/��=��'���,��f<w`�?i�d^Gm(+�)S{¦ �^P��4�
�'�Y{N9ț�dkjJ�M�ĉ��Ө�n��]��_�X�����81Ep����n
��5�e��b{�O@��C�&�8�xH�0�,����[��y��ؑl�z.`����/��p�@�p���j��gHU�=�s?ȇ��MU��VM���gQ\��1WO�^_)ΓyDF��A��w��ͭ�~�n�����-hŷT�&&Έg��'i�-� '�yg=Z���▓�/��������s�^�b��ˎ�{�Z;GFf�-��R��o�(x���n��90:10�aC�-��6��5�:���9�la����&^ Z�E9���2M_�O��s����x�xa�X�p��)�(-:1j(Q��A��"�Cذ �z�A�T�,42��	��O��iit��H�xzB��(|��NZ!�U���&p������6�?�śK�b�Դ)�@nu�=M>�8sF-�-����,���Ow�la�D�X�Q�����Gj�5�����l�\���逅�d�h������MM(�2j�����ˑ"�f�%骷i�,Q|o#��;�ෑI{(�Wq=��1�2��*�a���NL��Y{c�4lZ���j�+F���g[Ƶ:u�&^&���Q0%x7ϖh�e��M!O}HIh�����A_�-y�qe�~~,���Z�Q� �E�E�	yԨ9� v��>Q���V��3,搸�'��nW���,(^$�>�Nat賂��8��U�$��� =U=-��Afg���u,b���|r�DB���{��¶���#�݇��o*4�����|���gx¹ع�yfZێ
�V�X��y2w+yUZ�@CF�2Ib���n¡��^F�q�4>VM�nɸ�+u���cf�뷬��t���E<�P�<��p�U��02�Ư;�8̧1q==�C�QRO�.�-�����ķ��Rz�bW�F�i��le\�ϵJ��ۼ�2�8�����]�(O���Z^�8=[��fO���n��ޅ�=R�	e3��A�G14|)_C�6T�$���MW� v�; �Aƃق)����zT�1��O*4��?t�7��)S�n��9�^$��ߡ!%@h�	I[��^�P�Ƃ(DR�������w��\vD��c[�s�>4,�@�M5}�|���
����=���/�L�2%��8ó�/&3Z�*����!#��Hg�4+��Se�O���i���/�?}n�l�1\8T���ۣ�N��������g''w�pLb�F+c+��3���Nȁ�B�,�(R)�tE�eGd��t�h5IxO�ț�}��~2�r��SG�{q������]�W)�9a�n�K	��L�Wi<�����
iz!�f�{���;�����4�~H��.<�|DN3	&�^���Xn�"��^�f��O_�\_E�&$6�Ӄ��k���dY��ԛ��z6m�½�6�:��5WǸ�� �(Mw<1Jo�<Ƶ��2�(HR���GSq�KU�}��hg�����,���Z&}Sjh n��df�cC������E��O�@�;0���3��*��A]��X��?�U� ������Bd�9�Q�\�7�<D��4����x�e�R��!�H|��Ⱥ8%���0���k��B̨d���`�ذ��h�/��REV��u�&ŃR�rAΩ���
J=�-�gc{;Js�D�KC�����br���|ƯH�En��mjn�ăC|�d���	 �w��NC�B��!m�3�JH*�����)~��7K���Xgߨpz���
zz(t���IV�H&����@"� ���Ŕ�$�-�pE}���+��Q�x�s��F�ǡ�D�v�蝢 z����	����Q�ɭ
ϩ�����K���Sg��!�,�T���}���q�<�A������;1��*��q��C=�E�~�L��՞ b9�5��v��т��]�$ϑ^�$����-�O3WjC���e9o�z��qvg2)�B�2� Մ�������ke��ZH���h��3x&��Ǿ<i��Ufy�g7���\(j�������o�r/�g:���i��gf�0���q�{ـ�����^	tmrKsf�����~GT���@�A[E�V�>84�x�6�\vM����M*���!;�D�d?�@t�}/2]��QnkR��[�q'�j*W��(��b��z�2��[ۻw_'���=�.�v����魯�2�96�~t�ȴQ�y�S��>��>���M=�K���n���\&8�5����=������k��'��ٲ@X�M�ܬ5L��@ �g�i�%��=���@�1��	h�ٯd��f-���B��w���L��E��z�j	29H2F�oŬQ*^g��̹> '��aW�9##�[\~���ʇe_E"�DF+���86Zp�����f�en7���D7�8f����t}����5RaC���hFB�����sj BI+M��E@���[�QS8?6�u��OΈI��>%��Փ�)�_�C�=�1>��^��b��b�a��{o�0�E�S9$̼�O�9�6M{�����J���[RI2�>�w��7���+�ḣ~#|]Nogu��G��C�[;���d��q�?!V�̄6�1%ydWq���E�Uq�����w�<8�L��<�!NG��Ɂ��,�ݧ�+9��(#��7��� ��}`�o�߇��e����+Zs����Y�MqO���3G[��&h���Qa��ܡ�%���1�����ٖ�?Y���C�8�\y�O�bbͥ�Gܓ�/��>�r&V+}�W~��E�י�r�m�35��tDg��>K�����xꓮ��b��~x�T��k|�p��(�Ǐ���3ٰ,ۿ8�Ɂ�����)�,�V�S����&y�sӨ�EzO� ��7%�O
8G���g�?&Q��^��a����o��Z�ں��2E7���|�~���Ie��fNQ�s�c�v�fF篱����"݉Q]�n��^+��[qzoϟ�,f��j�N��,�`������b�k�LT3ڎ�X��dr�W���
|�!<�Bm��159qu������?����b��HC?ӴV��#��7��$+����D5�Ԑ���1������� Y��SsqirK�	�iu�Z�0�'�j/�h�w0�}2��ć���c^7LȓC��xv0�.����n����%��b����cRJs��k%?��p�8��ݐ�Z0��d�C�&ز��C]���!?KA�q�P�<���WP���N9��NDc�.��<j0�<�p�|�������-'�T���~��RQ.WCa�te���!���l��q3>yL�Kw^9��~��;-S�=�i�[�#(�nڌv�r���|[�?T@̏�<��?%�-}�?Cm�lv�/�,%�r�5��"���� 2Ns< �8��sN�'i���7Kd+y���'�χf�����>4h���À�O+7�J^����E��3r���M$��k��<-�+���č�J���t� ��/ď�j����I_P�?��OD�����fb�6q1������?��\��T{�aN˺^��WW��1�'@kQ���ÎK����y��{'� 162��Z:yJs�f�_�\��RQE�߃נG���G�	8�C�e5��<3CE�-\��u��W�7Pi���� �(�Ќ��b��6�
� R ���r2m���z��U����'����g��+F?��˳��Û�0��(9�1�N,R�T��
�hi�.ΐ�ߊNV�x�Pc@J(�)kk9f�,����;s56�O��|���
.)x��h�� Ps��s-.��zBG�@�|��$_</�8sZ$d��7aC}�x�2�Dč��!�n���]���sK�C�ճ����^�<��%�/�w邜�`wn|�E�UH�Җ*��G��3�)�Z��i}���KD����3*�糕��bto�;MfT�h5�*M)������= �fǷ���Wd| =���E�3������`m.��'v Gq���Uc:&�W��骄X	�u�~�
=�M�"�ҧ�!B*�e���ٲ/��[� #RMS�if��dN��.��ڞD!p]J�k#s?��8�:�v�a��_��V�KGo
d<{H6����X��		�#��H�<r�L!\]��e*�nᓇ+}H�5�U��5;���x�����@��>^��4A���]X�?P�λ��n#lA��V�$[�e��N�����N���Z��L�J�w;��6��$�ᢹ�騝84��	7�6�"�f���>C}2�F>��V�X����+A8`Z���� �������	OS�����;F�#L+ 5`V$O7#�*l��(��t��@	u�ew�d|��t���1���?�M�U*x�ٔ�1��r8��&�g�6��4NPm�r}�Z{�=�w2��_�uf��҈�>�p�?����,�mI_m[���z%�Eۃ�ۿAp�����?a�}m���6#�%E�h����ը�J���]$�H&Do��2 f]�;�B����S��������B�.�V;�c��C&a|g��4]	��f��k�p>[��'�̄n:i=�[Lz<���U����Z�)�8@��I/���1mm�3��t���8�z�{�$\��n;����t�Ř��\u">s̵�����d{���vA,p	��M�j�9` ��UO����}�p"�a���T���}��Y���:��U��A��pF�%��#z��.��ja�?�-�9I�D�=n��;Ӵ��7WQן�<5W@�gy�ݖo�vF�Efe`d�aP�n�"bMD%Cf�G��:C�����
����r�=0\KdMʵX&�_N�s�i/˜���zE��"�
������~ӿ�ŝ�-��\m]�=�(�p��D.tw_������dox�d����p"B�N9H]�_2	+������H��� ����XC�P�Ss��r�1��LF��x%כ�g4�x���Ι� k��ט
#��߶�(�7"
�bS¤d��_��b{F�
8���`�)����<`�]���tH�q�w��6z�h�P$1�/�jA�h�47b��q�+~g*�3KA�h����Ķbr{��,Z&�W}@��cJ�{�'�y�Zq���B���_f���Wl(0��3`f;)�[�x�;�m ���_�H�ͧ\|��K�՞�
-P��-ۻ�%.�V��9��NR��r��"L�ڠa��(�N���=7`&�|ea�K�ŋ���K0�3D1-��=70�g"��$M[ĝF��9o4�GCH�>z����^�mؐ�Օ�ﵭ�/z6�K��]�3��xlɣ?ˈf���(A=z��5��=�R�$b�@@1(G��m)�z��Drd�dRSE�t���?������FIt✾�%�p	�]q�NH�֔�M��tY�_�d�Qdn��0*t�0�a{e��V��g��o_y�l`o�.Z���¢+ϝm��;W�"���{a���t
|L1+��Ž��$��ހ�,u�5�rOY׀opcV|��Aޒ8�M������1L�����g��&���eR�Q�n����8�P5H���<�F ť"(X�z��ܡ�# ������dC����&�{Z��t�I�&�	o<O6{S且^%���(	�~^�#�wwi�r�Z��	;���	�a��{�}w��=ѴiH0��x?(�3�d����/]�vnW�\(��M��,���{_!*�;&r���=Ȑ8����{�	z�Ҙ��դwS�5�vi6
��S�0T9�TUz2AMW��5�ݸ��<��X�d��u�����/�Јr� ���I�c+^96^���aqMzt ?2*xš��rFkȞl̌ө���`hr�� �5�`��C8.	у�!�G~�5w|m��Z�-�ˣc�[=M�]����*9��=N:�F���)Ph�Y��K��z�Ȃߦ5��i�q��8� ��Q��0,/�\�>q�(i�XJ@����"9$9����(đ>� �^�9�4�yQ:D�}�����RC
nC�sz���š�P:{v�o�Z2�KF��ߎ|f��7n���jsox*�fh�"8�:MF����f��y��	`��YNs�T�EI&�X�ս�~���ϒ��9��iG~�"K��'wp<F�Ժ��2﷜ ��"
v��q��i'x�F�Q
k����&6�j)g�� C���C".��Xk�����-��>�Ň�(�+!��릢5����)%j٘足scA�h}ᘃ���'��?�p�q"+K~	�8����¶�����VMk���o��}:�v�l���f#���$�WU�H��z^8d?�|G�+��h�㔴�C�<��k��n�qt���=n� ���4���SIrHթT�TZ>|����~��S�tt���Xj�³���M4�*"ucMs���W@/�P�B�I�31�s��dZ�P��X��@��Q[k03$� 55������zb������{�͵��0����|��ЮF�?�2��4���.������+CM0��-ٙ-
k���W��u���n���XB�?	��!!`7u4tj>p����+��7����%~�+�#VY��ea�٪Yø�7�:������H*t�jn�<�5K���]>d�v�f9$,�$�u�=#��]���X��s���
���Q���z!mX&v�	���;bkʨ\G��ǟ�n���Ѩ�)h<y��:�X�Px�'�p�җ�f�D���mceF�tR
�>x|F/�pd3T"jb&�x3cB$غ���\��9�:ٛ���Pw�����-S������,'fvV�Saw�H�HZ�2�x,/�Q1�%�ό�\]�x ���is���?�4���MXuQ�o�X�ԝ��:R(����?ƈ��(�_���ܜ���֨�Z��J���I�[N�믇�?Q�M�aC5U�K�?0�\���;��g��"�-��S��%0m�#� ��+ﵪ�����W�@���w��}��T��]z��/��x�����,tZ�e�/�K�O�y��S⃮���Bd�e��ڣ�E{~�L-T:<�e��b�&�jgd�!,�k�|�s�f�/�i��TW(��7y�P��\��Hmo8����ۢb6��yc�OR�#�Pg��}�^����̖akSq�w��r)���) ���mbf���ם�+�	A�l�"?o�k�%x������ж��@@�~�
��<Y�V�r������5�;��P���}�
�����=���}I���qXpM��xpu�9?R�,� ��?���vL��xC�p��1�o���i�IRRl��ʛ�� M�g�V�!V��1���W&�˪U\ٱF���tT/���\MF��={$BrI$:�M�s�}�ҭ+۩r��dF!�1��9�0r8�U<��]�X��H�.�n�� �
����_��C�����#x�#%Uu��V_ʷ��0T�׈�(''���P��ݛ���f��u75q�V�\��Uߨ�/�@ة�N#���D쎃�@}�{��� wc�� ��T�&!_�.�Ti��!��^�ѽ u'9�9=�z�o�g<O�'
F�2�r k������s]F��%�vj�*�+�_�	2��d�': �*��&ǽ��¬��4A�hВ[v	�'�Cun�⺛$���Px�۬xJ�-�V��a�^�XA��� �����^�.��J����%!,�����E�N{73��g�Y�w����V�y�,��v���V'�=�g���:E����CW��\_P�Íގ{�����D.�Z)I)��ؐE�H���8��]� e��4Ozvk͢q=��k>�Y�눩�9$�:j�Bbc(�ۡ+ .op���X�o{�&�*�ety.N��dF:h=��ky���}g\y��	+���d���O�y���x�1�������uC��ji+�T�k�S�K��+�����GE��:fBar�R��X����5��g� >����!>��t�Pu �EN�F�1ik���r\��0R��b1teL	*k�:�?s�2r�%2�'�,=_΀TjjM�ϣN�(�p��!��Ó��wъ�O��GC;���Ӕoz�zj3�$��Ȯ�w����9J�bA3�RG�T�o��U�4�-}ڍ�E�36�HӘp�x	1�������P�'o��s^*z�3P��Wṫ��_
'��<Z ?цy�ӑ�6�l6�t�Y�JC]�(�q&R��Z\v�T��ͨ�bjt�'
c`��g+
#����9�?�b�1�2>����/e���?�7tp�<���ț�Yn&
�_�,pN�eP)�dn�d�8�'S���!����7A�RkJ6e�4?L�g����5slk:O<�3v��ˑ�O��6�	H<���<���d4�����YA�	1�U�c��:r�M�߅zɉ�^ f������)����!�Z�9����l�7v.���x��OF��v�x���Tf$6�j�-Ā[�w�)X r.h?��rkq\θ׾_��ў��6���d2P��%�@j����=��I�+&���@*�Ŀ(������'���o!�&1�Sdm�$�S��23W�Y?����~��	^kn�2��,���#V�1ϲq�����jx>!bȪ�{�<��n��;�S� ��c�\�@�>�s��?�F+8,'���à���)����U�j�!�מ��b�:��w�C��::׉)�����P>r���`�mY>2�*
�_��&�u�ۼ"~���ׅ�@�Տ�(\<]"�)I�ۡ@��9�+�$�f$6���N0�5j�����Y�v"LP��CeIK���'T!lCe���'U��fo����r��������U�F�#�s=���l"Ϲd�!GbI�C�F��ܑ�-�IYA�·(>D�,��C����T�����a�c2�Kk����ۜ;�b*�F��q̣O��4�DM�!j�o/+ƕ���x�H).D&�=�U�H���BB[q?��I���ɓ�R毘q'�u<അ�o�ۜ��d����2�iT'�cM�����/���?�dsa
�t��M�Ɋ�`:�&yp�u�`B.�9ñ[�� [�zLz(�a����"򧐡��W���ٮ����<�U�ȍ��n���ۋ�{�to�S�l0ϣ�`�˿��"
VSV��Yeҗ��\6h�G��.�{�% ���{]B��C(�h���|MR:�J��~��� }����9tM�B��#�%��wD��B����X�ZTnYF$�=�3��S\{��Vz~��jV�C�FNj���9`,�|���?�b�/Mj��B�γc��"��lON��x�T����e5�����^}}E