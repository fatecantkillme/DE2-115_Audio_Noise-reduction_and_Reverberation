��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<�\5e�)��Vs�{_$��c�3?��?��".�N���Q$V�'�	���S�ؐ4E��{f��|����d�ա�b_p#<_@ⓤ�0`��O�z��WeP�1y�k<�t�`��~qnĝQ~�_�rm'�&{��ރ��տ׻'{�AS/*�6��?O5�#�p�Q��p��ɂS�F?�0������jJ|�΄��P����ɲA'J�b�k>#�6���2ڌ��Y
�P(R�p��`��4�h�dD#�e��Ֆ��-��C�S��++�]��>��_�q����a�=�%�L4�-��6��.q�rhZ�7sw�$C��p�˹�?�'�.Z��d;ľ9b��pCs�����Y	���l��X���5#��I��c��}�+>�ՠ<W�PG���q��3�o����z�0k�kQk�"�cn���\�ԓ���oZ��6ֲ�֏x��@ =�%��f��M.�7�S:�Omq��@����Xk����bߒ���Ré�xr˵�Qh�i��	�-@��5/���,�}G��_>*HJF\�C�D@��=�-T��[_��<��_$��͙�5L䦯pI���N�#��&����\(V�w�����)�ɓBš���B{j{)W��.K�D�b��$�{� ��5�����^���BÃM�[7��	�Mc%�$�/ONg��� qO�L=t��R�J��Ų��͉-潡��7�s�~IvŦ�s����n�tLN���k�5����!b:}U	f1P��P{ƥCB��|�:��� ڧ��ɡ�J�����"�izva�&�-�nR�d��@W$z��������x�0�?�J�����eŨ����!�V+�������Y4ʂ{yBG^Ǡ��T"_������]��u�V�|z�>l�>��8�������\���k�X4��P��ǎ<:�<C�3U�u5�ր�t�U����BpY]&qZk�@��s5�O|������2����6k>A�߯��r��p���|�k�aJ#QMu�D��C�{{P��D�R�8��.��a��'�)Q1�s}�9BIm� ����-O�2��b�w̙����G:3䜂�&���3��Y��D.)��V���{X�C���m�	�Fe2���s?ʲ_�����|1/At +���Y��%�$��y��Bՙ�%��o�w!Jw/���Y��V��b��>Y�Ҥ ���OS�0o/J�-Eթ�:��0�i�Fg$|v�~�>�q:�o�t+=B7���`v�V�����=��킕^��Vf�-`L��5��a �&c\�ܺ�y��H�^ĳ��&�I��X�_t�G
��l�o�,�Z0 J�:�]K��[���~���	��+N"��b���S�N/�Ś�_���)�Q�Ҟ�b����>䎊~n& #�c�3���/�t-W�����hF
��Jo��J�>rV'&���� ����lx �a�Py��v7E�_V6<	�E�ʿ�.�(�J���~�q1C�)�n(�
d��b���pu� ��M�OM���RqPx	 ���6��J�Pv��_ܧ+��j��Mg���m��'��o�0���c����s6�8���\f��E�۸N��50���?�M�$���w�W �ٞ�[���q��X#�좟y��t���:�����V���0]�D�.a���@S�p��`	t�溳�������դ��	�ro+6�˗�ۢ�<�Xf�E"n!t+mGr�m�])�Ek�Do�-L!�V��Ϻ&鋲��`/�����Wo��9���<G%7��2��U���#9��?��0tWJ{�`�挠A7��y�ʑb�i����x\f�6��`<3�+��sP�ZYwמNo>��w���;`(�Ҵ��YR��]�����t�:���b�����G�#������/XϨF�9���l�]�밎7� �+�����V�ܪ0���	vy(x͜��g�iQ�D3׼�y$�=�(�����f�>��~6RV�vfc 
gjyJ�oDZ�<�X��J�;�g���lgX>��F�Мxb���_z����
Uf�'N�˂?�#��S���u�dl�/��tTӁ y[��mQua��l߬����ٙ�-��F�Ŷ0P��[c��,Rߙ�<�IKt�&qF-��Փ��1���_��,�\���݉��0?���,�����Uj8x��XH�Y�.TDV���_*:���a�~��;�SD
N�	��;��{!3cm�����D��
~��릙v��������R�c���T1��c@ؐ5�c�X6�Qa�{�S]�Q�+�`xu�L�:��x/�ҷ�M��b��i8]N�L0��,du�aL���|u���ҽ��@��e���
9�Y�y@�S�d�?������o�H
�-���ʺ�Lu���?��-/^|l�MAU&	���H12̗ç���?,DC�N����2+���^����~���Ă��%(�Rp�t��on���ɾ*A�In׏r�pu �8�`"�h^x��06�_�P�FF����5�y|�,T�%p���D䞾��ⰸ���U���P��6h4��b��C'NFW�	��a�(~$չS������ȇ�G���<���L�R:�@:����z!e�u/��U�(hx�&�6!%���eȎƫ
$���A�!4���[?h��|������ ���h-.�Ek��EG����[]�r��Pxvµ��Уp����s�J���ԟ�4�(����j*�0�ߙ j��&��N0��˲��<�N��U����'E��ty3|��p�AW�����஦~��y74�'�l��P���_wį�E�ٓ:�!W�h��U/�9�D]�cm�4��Tdn����ܘХ)�� �EԠx"!�	����%v�w�RlOVɑ�%=|��53��D����� ��q�z	�䨆�f	�5�
�!�W+�'��)5�G�n�8�U�w�Zb�	�w%\�"1ē��붽?��j�� ���0�jӷ,լ���_)O�	p��4{�Tl𾏇~�-�{��=�b
���6��ڗ���P+&@߷L�X m1�f��m����F�6ʪ���(�k����3�iw�5�3\�o�t�"��ݝ��Xq��Eƣ�=���P.� ��h����7�m@��+6J"3P��y��^t)9���نl�;t,�'B�:���ԓ<�����9�d�������X�wb7*�um@�_��â���,{��M!ߋ:�8Ut�m7kvgtާҗ$�d�8�	�5�d)F�m���c�`�-B�ц�ڏQ	�x#��l�.�T]��A+΂�,�?�a�r��?�rtΤ�@P�ўt%���r=�_]z�{�O����'|ח􍓍�FYM���^�J��-`KX+����G�l4_���::q#7���@��������Y%П�0kD��Q���[�8N	w��=�߸��\9�+`�����!�Kâw�n��l��:�q ��l��pT�l,+U�@��[&����&C؆�ܒS�o��*�6&���ޕegs�տ�$P�G�T��JeT.�	�M�"y�,�=,!��7�º'J�4�����_OI G3�{��$�������(V&>�F
+�j#�#Q�|E�2?閾��������1�o&ph���ח��sOW�}I��Gj׈@�gVq��3��yX��6�lr�J�4����/��I��9��똄��B�)���1��`�9 �2L_a��=K�ؿxPτx�*����.'��J���a���J���$y��W ���J���/����n�X2U�mV�2��cJ �N�(?��z��򃃯��[1���,R�O`pKش4\/ :�?���F���Κ;�I
|>����b�[�͑mq�MW�p��\c�f��QS����̅%٫H��
.�O��mE�;}� BҰ���(�{Yyq<6�[hm|%��ǉ�վ���9&���B��@5+M��뤚��*��B�6*�^֭°���NT���;���in�YV�e��3��A��sLj�4��������̕z��6�����&�~�
K;�8}�."�$�za5.7�a�%�����Ô�b�������ۢ�ʖIa���ɋ��Dd���H�m���y�z�����l�+-sF�i ��Q4������h{�u�;렊Bs�V��n�^�,I�^Q_큪_�� %��=�?:+��F��jS z5�MRi��i��n��1�".i��q��{'�J��U�Tj]�B.8!��
v��F��}��g�o^э�Z�9��5��c���:���*�P��0���s�d�F�m��+���	�I�v��G`�x�d���Z���l�{��x�����n��2,(��]�gt�
vG�HU�(�y��G (E��+\(I�d�=����J,	|�x)r��c4��N���.� 89\��_���w_/H&�F>;��Jͨ�����$��)i��-ufk2��L�!D\�����x��ү���edR7��T}�m��~w�
HT.��5�#���YG�����;���P�aB0�S %���'uaݗ���S�Gop���J)�]��廥;^��̇)�J��,����G�����.NX��N���AqD�wh(�l��${�b��g��f�@�F��Y�ӫ�g4"|!�_ڴA��&�<9��xR`�>F�)n�s��U$a��Z�B� ����e�Hx��h'�t�GL�^A��	ܰ�����;�m�;{�Q5�}�_�5�3C�.R�6ڪ|_�7f���i���7��e���0�<���% .<88���jwC�+�̿
�hft�Q� Ψ'���}[� n�=@z���� -A\�5a^ ����� H���
�)A�%/c�u4r�i�t�j�&�g{m"�cG����wy�tt5�q'��	�����:��4N؏
k�&��	Zb���m��xۗ�*JWh��g�f!B����'���`���p@͉�_�ƀ�O_|%�����p<�Ў�J["�6�-U�������KN�Q��n�%��MW�K���O�e�O�JA��_��Z�x���{��I��z`ϯ��I�H��564���Yb�.#�%���P-��@so�T���/��E҂aL�I�Iا�N��.m��ۜ��E�Qؐ�������������(�D�U~�K��42i��ƨ[�2o�LɜL��:�(�����u���h矔�{ЪX�{�E>iD��P��Ԑ�-LO��l��9�T^�#����	H��pq~gW����|�C5|yAf�lm�4�m��������K����HU��)1��q��A6e�,�LY6+�Hk�`�LOK��[k��	�3�IT	��wnl�r���~�'=�d��8����~�z�HH8x��ݍ<��tW��Ϩ�=������7Q`$�eӺ",�?D��w�����:�.vBt	F�X��(r�T�j�u�}���ZL����X(3I=s��1����;d���}�:#�k)F�,�N�QOՀ�걾��sL�{���8��8t��?�0\��LeC�P�ˮ̢��BO.�n]�y�^݁���5];	n��﹑�7��ڝ�,�:$��;M�4a|��'y �gMYt�n�oJ�)�	Cu�q�+��* .CWn�O��1�M�F5e��3�ܰ��,Gb����'E�~`��1H��f���t�6?�_g`|��D� �~�ϑU��)�ȝ�2����{�sN��k�q
�!
3�#zx>�Y;^=��x��� <-�94�[������?��jA�A���*9~���x���=���ֳH�����ar�Gb��*�nؤ��F�8��hu
�t!����dBt��"�$�����?����O�e��:��]���=�A�.9���p�u w.���/���&�;�Gŵ!Y7R�ģ���<�Z��gy�K'e�@�ZpȽ�m��=����x�1��ՠ@h����˔���Ѭ8�8��_Y,0Jr�Q��`�%�*'0��zB�'8��������`#l��'�����9���y����z�M�w���>�B�z���_������
/��4_iJ�(j�ܾH(0T�+d�����lk�n�d��Cb�/-t�f�在ֽ�m�� ��&��$K�����Ru҂�W��yh��Oa�S緅*V��3��M���9d(�O���R��
�4�BAG��w0�h�LToS%�e�n������?������%�4�c�<���s_ĝ����[F7��o�� �3�h�I�| P�3</���V�&�P*��T��p�7,��$��F�X�#�BX�O��;��zQM�'�@Y�}z�����j(���m�5G�
x�5u�U�x���#��n��;�:�}�̭�?B'z�K[C���z���Au	J��V,��A���{���oVGWӴ��<�F�~Rr��c�8�"&
�'�1�X�#gMt��&F.�C��������k�&ȥ�G[�w�A��i��;�^*��_������I��~��#4g�*�nC'n����P�\ƈ�NUR���������а������0@�(U�l���D�G7��/bQ��'9�n�L�Z��Ct�w+��!Յ��Oi�KgO"�[j2��|�S�'vualR ��y1��5E8Bh�Ud���1��9#�Zd����>�{c&"T~���
�BZ�$�(M���ey��]�M0wa'T1���G�)�
�Ep�5�P��])H+'V*A������MH<\@���q�T�_a��:��e�p�8�ݔm�CB�'a�{e��'��M�����T����(\�¥��ŋ4��P�x��<��Y>b� %�a��� Fc��^�ŋ-ڪ9�OiCsm�(ջ�2��T�/f�]�6��0}���*�
��+1���S�z�E(�쁪�2��Y�va(��`慇Y!��,�L�_mV���5���e8��������C�H0FխS��u0��C�?�vv������-7L�����~*���!p���O��:I�Ҳ:��m\�p�Kl���"{���$3裫�[F�i�NI��ң��_����rq9�3����/E�rcM��#��"d-�z�\5��^�����Z,%�,Y�
�dm��he�H�Ré�.R��MTO5���9����w���!3F8���{��N���&���z���*��$r��F[�����:��l�o��0�|�D]�"��o���s��d�1W��+M��j06i����,Y�?Ӱ�'#f���@[@�Ct�$Ko�-U���kB��q!�-�{�=X̬f��6�]Sx�%��s��)k�~��Y�f��*8\�Y��K�rқ�j_v��)y��ky�O�BK~4�s^��מB�f��`��%�~�#L�,�Y�mz�*��8(�Z���Z�7D8ˠZ#�}���@R��0-4jXJBNM�%�=��EX��o����PC�׿�b��z��N���2�kd6d/
��F�i4u�I-x��7��I�h!"��	��i����Eo�@��}I)�냜p�o�=�)F+�fLc���R�Y�R���C����n�/��nk�+m�k�K�yn�k�BEa4/��Ut�tnT$�����(�E����&=l��.�GZ��A]C,��T��D�k�2׀��	C��O�����P���$9�_gh�0�ᅦ|L����d�Ž���U� ����J�`�j�U
9�"�I�GT�.�{��@����YR\A0�b��N�����H+S�w�z��� p ۫�T���M��vN$�s�1���~��	������1g|�3n�`F��f�p}�J^�G5G�\X�4�,&8��Ɛ��ʷ�K��|�����kE�P�d�&�ݘ�8����_�%U+��:�1l��d�O9b�A�m��e�i�wZ��n|�|�Y��F�(f0����M�m��!�<]X�1�=���X��i��o�%;6 Y�vo�}��F��ow�����F#��Q[�3.� ���Sq�����
�=�����k�O���$3)�;D79q�Zw�ί^��=��������;�/"��= �Ҵ�Bst�"�����<n���i��|�c�y�G�ʩ����pf6��$�R5�!K�p�L1��Yl]�R�zߞgV�U�M���V�tŬ�i
S	H�J����B��;���U�D���v��D?��j|��؝��M@<x���fW~�j��L3�r���7�4L �B&L��-}�Z�K�iȏ�ei��z��v��1�j�w���*��s�okr��)��app$�d1ջ�7���5�'
Sq�WE�a~��zɺ�A֬d���^��jE���w�8f�h����`ٞ��I�t�����Z���*y����m��˞=��c�Pˮ�1[������`�g,wG�3���?�d�'>�1���8�I�� ��ǁ2��؁osL��Z�xw`ԍܦ`N�z��<�n0O�[X� ��&^���@4��ԛ�?��y	�Ǫ�痶�v��yZ[�^���{J�2;=����U^��ҳ��>������	-�D|�h���Mܽ)���q�G��U1*5��2�T���|����s�+��S�\cʞ��a��/�s�	��G����Ϙ��,b�G�	��(��Lǒs+��2��kٽ+�T�7l0|PgK�)�� ��>l��U≓}�Kf��gQCI��z�*!�b�@e��˧a/�tݷ�l�m� �c��/ �k��ain��?����"4�����L�yC3C�V�?VDZ�0{��%���so.����E'���F!�����H�]���	��D�����Q%Ϭ�9��]��7��H��w��V�U�F�t��L��f����1�bF���es/$�T�`n��y���v�n��N��T��`m��ƀ>??w�Q.�W'���[f���s#j�E�^)�6�����u��Բ��%��Jj"�B�=�����9�&	�q��\��js�@�F���,�u{8�p��`6�09��X���k�GL�X��Y�u�n�{2����14�g]��h���i��n4N 	��x�12PH�|��pD;	�!P*�b�(�p�x��)~<����Qm�C���mu��?���YD����|�e�;���Oġ8�K���<�
9�#���XG
���$�<�I�:q��t�]��E��Zo�/�I�*�͕��b�ީ�x������3%.�<�Q�3�e羅f�����v���6~Qx�q͵���v"W�zhW�^~La�.����}�F�b.�Ć�Ha���y�w��t��0a�b;*"�L�e�"����[����$��c�lVK�t�,o4�Y��;��@33z 5�E(@2���m�����K�%n���.��U�11D��K��ˉ���A�M�꼛/L�B��x�i�^�z�xl�g����E�� �rn�F|��38�_0�[�Y�_�������cj��>��ڙ�E��[�C���e{Y�0�<��d����u�n�����O�e��q�R��M#KP��f��:���W�+ZU��n��Ӕ=�|�@VҊ ��*.f��USu�r�OnW���fK>�ʮd�^/�7v��
����LW�ah��- ���
!! ͪ�*ni�z����`�E�<'nl���:�`�ڍu� �*�W�3�1q�*+`��'ty+���A����p�nLb]��!1du��R�cW��YFM�7v-b԰C?P"�f��|��rV��y]�&<{P� ��q�=���x����n���+r�>�Sǰ�`u'�25��DD�&�'����l,Xu^ ���%�����/v�$Snj���;��!@��BD3��!�uoR`W�O.Ȍڦ��$����"��+ɑ�*��ߎ�Y�3�ŮZ��G�~4���_[BL�@�P��M�4#�ֹzo�_M�ȉ�2n~������u�s�F�M��>y9w咡5�y�p:L�E�.�V981e#�v��9E#7��}�+p�Y�rˎ(�����4��PT�WE��n^���w���!����U��:�{)	[Cn%��<r`kb�@w2����T����O��؂�B�uI��.q�4i�Oo�4	R�C����엣0v���*2�^��3�@���EV�q������X��&�BBe�yb
6@Y/�)F�ڃ�#�z}���>2� ��3n�l$SA�R�!=�W@��EA�2��_�K� ���1d��/�|}���ȑ�O�׶�o��HIʪ�f�#mT;R�50�J�ff��m���ڲ�0�RP�F�M�2�Ak±���Q���ܖɮp�0?4�Գ�V��9��/�H�)���l�Ń<C'ڢ}��qK� �ݎ-53*r�����`iv."�A8z�R��H
��:���r�Ҿ=$r�0�W���y�აodH�!xVx���#>쇞ٳp�ۡ;O�IW�zc�� �r�&�Ɇܬ:��m���,f����u�o"�qS�|���9�p�� ���,�9PnZ����h�;f;iUؖuSЪd1諨�;�%G��z��`n�@��W�����O�* ;�jH�������)Kή�� _-R��S���o�f�`W%-'�A&��+�h�|�×��DH:B�v���~�JjfH����j����(m��E�0!�z��Rk��*�pK�`1�ݿմ�а��.:/�~�9[^n�1xOq/�Q���@��4�y-�_�Y��+����-,H>8G��RQ �̹�i��T��8h3g1q�	uI��[��)|r�\ɘ_P��fK6��O>U�li��ͼFB�u�q��d��r��rd���x�z�� $������M���)���¯\�J1�'���V#њ�Ne�m�<�6�#����,f�ml���'���r�ㇺ
�v��h���J����$�B�\�~ N.->Y	\� �T���-�E�Cv���A�0C%m�G��S���'�C��1�[G���}f�%�8�ٲk�&;� �/���P(E�f�����u=!Ṡ5��"1��w��+���Ϋ�6�qмXW�4b�;������ʵ�n:jE���B��d�2-6Uʳ)�ℐ�`���S�^��9��/�����bB�"Wo<wKJ�b\s&��ɍ�������[���q�l|�]N�:����vU0ۇ�H�b7�<gIဢ3�Gn���S��L����$�>�1�% Q��w�!��Z<xf	HT�GE%o/r����T �������2�C>�� ��7��t}����%�"P�`g���_��}^���ڢ��������
e���{y�O���wm�l%(�Pn9dl� k��LXb����S��RkO�yQ%j(���J�2��I��>4�q��?�Ȑ���l竑�3p�o<���8�(��Ó����L�7U�j2�N4��dZ�0L��\8��c!r�B�6���88��ǎ:Ӷ<�T���.�b�"��E�0RFު*�����v)�E�x��h�{�lxOJ�^�ff�.H`8e�c?�c�K2G�5��ߡ�u�P.��ª��pĊȯ�K��d6/�:���su���\H�lUy?t&�TD�(�2H+0ҟؙ�&Yo���>�6/�iP%���z�ܵmFh���#��ů�d��)�6vuuj$�`����0����<�Ҥ08"BҔ�vN��Ӧ�8��JAB����p#��gU�%j¨
b�����~h%��+�Y��*yFՄՈNy˄����E~�1��&�����drY��i�Ó�"��r�S@����n��h���E/rpp�o�_�q�e��*0l���NzZ�g���Xȗb"޲:��.�d#ߴ���ːzmO_X>�������5u�Q�"�G��$����O� }�4oJ��7z/`	[��u/H���/C��Q�=�\�U.�	W�P 23$W�������6�&FL�FK��U9��5����dd��)�(UvjA�0b�X��5�{�z*�aܿ����c*��o�6l-�o��D5xo!Y�P.5:���H��*G�EV�7}�<2�)�4#�����Y�ob���w�[v~Ũ�^�r|�,��=cJ%�/a�
:�^(3�V'�/�f�̕jÞ�AF�TT���q�x�o���X�p�n-����[�-ק�CL�s(ǘ��f�%��D�>�6�Ox��cw]���k��Y�B�Q���h�*��/�I� ��L�*8)�i�I���Ge���Z�㜜>.�H���Y�G�o%��и��<���9QN�7�2��TI��O駾����R%eed�����f��G�Q��ܟ��e�\>�I�k��\WB�dk�;��L<iJ>~6�qr��f0R3��>w嶋���F���Eѵ״���0���	��6�ˊ��q�M^\��}�Nzn��\Q\&A�BJ
_Sp�0|�.��G�Y��O�c��{��0�Iܸ�Fp��_�p-|�T��Q�m��FH���L�����_�ie��Ϝ��+�s[��d�"�"ώ��ئ�fw�$�s1�>w���cz{nu��у�t-��խ�o=�8#��d�����11����C�s��Źz@vD6A)	\:�%���]������N�t��6y陉��T����� d[��I~7#�C�+�<&�?�O�����s�8�����d��a��d��~�i��`���J�ea�~8�	xiF�I�>����2(q�+k��=%����'�J�n'����1#a����{���t9�CR������Q�`%�+n���-�T+�r}g�[��x��E�j c�k�z��YZ`چ�l�&\�`�G����RI��Òⅴ�x�{�5_MDN��P(W�t��G�1��-v�%�P��P�آ4�b�|;�^�"��*<+y�e�\{Kl��ɾ�msW�R��)~�f�)Ol��+�����>YnP�<��v��_����z��cF5����!�x�mw���=1?g�6��x��P(��6�k�C�]RKN�e�18����p��,:�x��R�2ڪ؎��ţ��=���#GE;2{(g��d����;����d�Ev�y����%3�^L�_���m�1"�쑩@`ﲾ6-@�f��^em�:��/����?�@�;U���^*�;)劤ߓ^U���6ֽr�^^������ٵ����HJ�#�;����C�$����qE�������H�X�ψ;��q�ψp��ӗ(a�HƜ3�~��'#����i�bX�C��\���@l�����E�Ȯ�\ik�I�j{��s6�Գ��a��!����nRL�J����C��t~iZ��HO� XM�:糜�>�4L08,�+��m9�tҏ{!��yz7T�Y)u��[���!Y@�"��)@XX��'� ����E�O�Rپ��l/�,��[��6��OB+|vYJ��A�+�R�lx)[��k�7���S9��QM��*� �$��N���R�՟y;-�,X_��,Q��5��~A��҉XCR�_ ���c	�+I|�Xl��3/���=��<�� t���bЬ�0<cP	�n�v0��΄�GzS��9"��W�^yѾ�OV���oɂ��aȌ�ժ�hp���`>�?�R�S#th��h?��3�/�Qz�o|�<_�Ƌ�9�� ����j���䧑P$�x�Ll� �S��x�{l:>z�/1%��ȱ�Z���Y+}a;C����ۓƉ���\������L	q%�!3ٳ����8�y��T�������M����C�R#y_`r]rq!xB'��A�$}	�U�G�k��M.׏�5�鬰-E�&�G���T1�$�ۈ��ݥ`���R���Q�2p @���,�>c���_�.uQ���jNr��k4��ޞ&�t-{������rZ%��XoNA�a$g��[�N �aϷ�i<�e#���Ob�a��������$II=�x�����q��Ge�_���+K�Cjc�S���ں$V��X��@G��H��t���1��՝�;�v�óO=X^C����5�"x؏�����l׉�=��	y�W�zc�P٠��mZ����q�p�}w��J*�X&%@w]�sӔ�`�O)F���a�g��8�\�6�(�(bo�x"σ	���&M�r)W��*:|�:F����Ze�s!���y|���^)SZ�VhweQFZD��)�'wR�J����H�J^=b>x�����Is��=�J�v�
�A��I�m��!�Vڻ�|�#w�[���WR�bx�|����Vt���f��p�����ƫ"��hLue�Qjn�����*�S�m�27i<{i�:�)��񶁩��4��M �d��J�}�G݀�A�C`aV,���ya����J�=!�d>;�fF�ו����Z2�{���#.x��y0� �UD�r�1[6�з�%�<��|٧���J�Z#L<�8T\o��\ �qL[���"�n=�5n��&C,�� o��Po�4�5)�5ȏ�B��#!�Z�H;�LN��-lG�C���ހ�����'���gE�}�,�� -!J�݈��3��}���4	� ��9Q.�Ō��	2Z��.���R6��(�)�k{1m�r�jI�BmRtlր�v9���!�,˰n\����.�H��5^b���R%Km3��*lO$��s��]��eb&�#�E����#��=�w�e߰�亭:+Y�Q]���� ��Ī��D'1FA�K�dV%����[�.w�E��sO��|�-���0Aw��
 _��׮*5m����=�]x������SY|񎮆���X��:��0O��)#�(Q���g�2@)hH���1�6s+�ce�,D��21[MIc�[_�7�踟��臶��P��2uW�7�s���'���}�ra,6�#OO����m�F�,u�|y7���nL�<�A��տ�����w0���2D���>&zĘI�S��@�𛃾A(ġA�(���p��� OeWve��h�FP�U�Î�Q��)���k�~K8n�Rw�=q�=��w4��T���%��;	�J8��u�&�����%�`�O�#�T����J5f6oi��jr���3T0���g��Qy,�b�/,W���Rr�� ���,k�E�α6�r���˫�n���O�6�~���2<�	� �#C�hU82L�������l��b�����˘԰pR�½О�	��ĝ��b�)&��@�$����3A
�$��P�mj5& a�-�{��e���?ӹݐ�i>TH�כx��]��{-��a�й�A�!�z�KVy>�؄��)�w/0CN�˘"9������,�Ĉ8�7a�C�0(�-ۏj���P�9��=)7?K�b&L�+e�,�!�j�!��קּI����onad?qP�TͰv���`�@��5��Wso �t0C�rw�����}��s�"��Q.1�B�ޱr@Bp�L�<迓$���)I��o��d�=��#3�����ָ�F?�3��ο-ln��/	����q�٩L�lp�����uH�a��)��98�<��Ls�E�kGdcG!��̋��p��eN��<���X*���3��ouJA	�f���Qb�B�Z��L�y�����]��V�"]�����*$��KD�j��P�����0a��
�Ь���X���9���H�]�2.���[�h5���]���֟N±L��>�;K��*��Ѳ�B���w��`�Q�l�n;��k W0B����!ix^"��w�o�����	*��AX��v�|	A��qU*���H|��h�78ħPE�NT�u�"���1�J�I��G@�S���)/9��v��+=8?��=v@��C.0�U�.f�^�� 7!����e����v֍So��`����B`z�#;�W__G���2�J�2�Mٍ��b&b��e��u�ۚ��]�Q�t���b:�Șm��;)��{V:��:hrf�:$"���ks9ň,��x�$�"�o��8�C���hT�d[j�8��O����	_�4�
�I�<���w�ڸ-��`,�/K��w#�wT'��H%ő͉In�GV��ϒ{��Zt!��+��mUO���1B���T���|Uv�_�����/�af�������<ef?�\P8uF�S�_Xk��|:�-�DCWU[��O�K��w�H��E�hϤ��GrEH H��]S��Й�4Sw�&�=>b�K�ˋ�V�g��E�ME{`.���h �4׊�}��� ]���[ �����7�%'�/�9P4XMͬo�t�<jaIeA٠���A�Y:NA�g7O]R`��A��L�~��#Z"fnzMU.���v`W���.�ߚ�꙯�e�-+634�1#D�eK�Z6-�,Lӏ��%a���[�S�s�#�\L��7���L��ڢ����E����a��r���BN�V�)���� aç^��^�B��1����%����)p�[a�Pg��x�]����C� 6�F��Xp�$ʥ).������w�R�����zT\'ur��Lԏߗ�ـ��D
���դ����d�co�`��"߻�n�aβF8v�R}���0
�;y{����ཛྷ�Ž1L�������Cn������q(A8,Wp���W�r����^�[�c�W5	��P~q湛�d���L�	G`�<$8zb^5��E�U�
��KQ�fJ���l͵/��E��(��Z�EpKt�+9t Ⱦj�jM��Ʀ�}�]��|�\�D��w�����N�gA�F u<��Λ�p������wy��ٺ�͚�`�i\�����ʌ����Mt���*���<ҳѕ��tm�Ќ����:r��Z��r��޶<��i�;Y9����]��M����py�
�=��iuo@SM�2�j���$�dH�Zc�U|G��AFG��zm�4�pP �r1-����=$
��G�'������;~2i?�.T��.�H�����1���9�����sU�v�bL�Bd�i�\�+��7�C7{��{��"x�3��U���=�&VX�z�r��|k���~�)��yY��cNy��2~����V��>�-�;i�T�:[��,�cء�,d�����ߑ@֓`憖}'_�?�2(��nPp�q��TW+]˨��~���\4���\&H��ECN�a�:���x-������=R[�S�0���ʎ,� �)���r���;R*n����v��FDt�~�1�ˠ����D�8�=ɐ�W2�$/ru�vK���N��pz���`'�.�0(��Y��A����R��ጛR��?�-ڹ�������g\xkL��5�v�p�}&� @CEq����c�n�6� 6s�'��(2jP��9j9�"[@���0�qd
���?�O�"����Еr��(����Y��֘XNűe�b����/���V:�%�ƍV� O�9�D��sb~��}b<BI�������%
��/��'�Nu�\;�Z	�PG�r��: S(�'��ՓB�xTA�:I�S��0���}���S�.9��!+�i>���e�e�?����˅
#�,7��_}�H�l/��'�q	�
vՆjU9
ݖ}�)F;5�m����SJ'��KD!9Y��ҾҠ4�g&_�7�So��v�hX	�{��4~>K6?��n��^K`��!��N�{��J2v�l����T��eh���kҰ��!0�A�1���9��.r1�\zX������K�r��ܽļ�oڮ�s�JIJ���ZA��߸�gYs$5;J�o����G<�ɣD�����+h�p��OiW�P�ޱ<j�*I-�X��~/�	:����n��@LJW���8e�'i��DZٰ�L���&�ܿ��ym�}�S�%�14AF�YV�G�
2r��4�گ)!,�M�H��@ϱۧ����;gm��,�3:�ew����i�Ǻ��ɽ9�X��i��׫^SZD�<fڄ;�m�g��0�n��Í&O�T�Y�`��-S4]L5�ī�u��K�A���d�^m�m��t��}o�QS��-O��+�`kO�EV�P�?����@ѵr77���K�YY#Y�uu�8xc﷥��&�Za�P������̕O@+���Wۼ;1Ǒ�	c��E�r�̂�N��ݮ<;R)K�H������I\ �`�а離��m��G���@�
 *؄n�[Y�mk��/S��.=�������x�9����C����ѣ��E3�0���|�e'�����v%����d��y��� ��m�dmQ���F�j��{�
�����������l@���J��݇d`��E:C�]}�#����n��*|��@Q��#joEq�,�NH�I)����R����¸г���I��:���jsb��XӔ��ʶ����fv�<#�&fա��n��<�ʞ�yNy*�������əJ�ſI�����|�Qĕ�$u/!=bk���L%,.�њ��R/����cw�W�
��*Z�k{S|��6���� ��6�L*����?BD֢Lw��oh#˅�z�r�_�( �\ţ���
��#�qE�ia;��v[���m�*�l��!�I@t_$��JqJĴj�80�o�PP��f(zy뼧���8]�?��ؚ���F(y�ӝ*�ηٛT�m F�*���)������,~�����g��2���}j)�/�t	�?�)��@!FQL����3��<�A��H���H���=��}�&c�8[�l�e~{�J�c֠�7_+/�4�Q�DV1}���_�q�#x
���5g�J�QrMn[��U�J]C�0���+D���6yk���r=ȶ{K����[�I2Qu'V���nB�r�**]��D��*a�6Q#Gc�F�i�6CP�"Rs<(OE�-��q��)�/��W���#<�P�E%k�w��W���%����Y��wp����=�)a��bK�pHQ"�_���묍�̕�k� �To����*��(
��,��Hѻ��Ѝ^���w�oFE2��X��v��+�p��P��9�rW�M�q�\��G�8��^5��p�3�h���y�*�� w���j�Z%˖e~��5�B�9ׯ8+XHu���k�ސ���$w9� � ���=�@���Z
��ؖ+����`j�4l
��c����$K��/'iE�["��=F�b+��XEV�s2 �ۉT<4����yǐ8�p��/���%L����e
Zp]����0cTL�c^@�r7 �֐��QF��8��0���V���7=+&8�L%��>�`�t�������т8���TotE��U[�J�-���  �����U�m`��Хyf�#���5�޵R���V��{6�(Vu8J�pv��b;��|^@[�I�[�Ȧ�k���J��ӑ�ty���L գ�6q��p�|���̯Z V<�w�̫:���|��`�A��Oh��=�~OoM8X�op%aa��J=�>�����8�*�H�	�1[z�t�R0��A����QT�L����3�0��
��ze��sx�Kxןë�E�?����C��y�^-�~=�B'��9��\}՗��ل�M�|_SA_�|��Ѝ]T�f�<����F*��s�s���\�U���R:��3S^������!���Z��n-��z���ؙ��1�E�-�Z�A��0�Y�B�g����oP��@n�{O)���IPk�pNocQ��)�q��<�i��#�G$����"�D���1��Y���o�.���y��k��A���lh��= ��MD�.�t����
�[��l���'c���C�	/��>y�����n^]���[,��v2�m`�p�,+r���S`'���uf̞�3�o���~*�@Fܸ��R�=�l�|�����INI��z@X4�q��o�h��AY0L�*��7�!��Я��$ ��gߕ�
X_ֿ�fA�B����"�8��&�N�b�h��/PDW�tϫ1�!p�(Q�]���^�lIՙY�������d��k����5�$�ᩎ5�sz"CŪ;-Cьa)@d cܭ{�'�}�������2�Z/}0����(���ъ�Dt�ц�� 	�����s�� E]$܈�A���"Qz0�j*!͘��d���"s��>�T�U��/�ꦥ�M����1��4�U��k/u��*qD�f��>�Y����0?w�Qc�]kм�{�M<���6�>����9�[�&:��_dQe0n�H��\p�ؓ����1��v�\1E�,����T�gK`h-N�V���l���U�LTRgs>N6#��N��VXLx@��{�OxM��BL%�:�P}ݞlb������V�hN�=��`��S"m�$�	Y���F�̷]�m��.;�t�K"���H�Y�����X���]I������2�&����AU�^q�&�Ql�Ojr��-��4�l�ȡt�t��J/J�2�G%S|�ha 6K�%k��Ê�uk(��d�L&�G�	0���7n|.�vu���$c��~�T7TQ,�_�x���y`J� �wC��E�!C�e)7Ҵ������mi%m��n�e�F������;we�ó�zyKH=��N�j��W�>@1(�iAك�ɷ|�!�:ƴW�gI� �����!;�U��N!:]��3�D���v� ���o�onܥ2��IY���F�%s�@�{��qzť��x�n� �q�8��P�hā�=(@��42,R���������Orv �X��?�"n4�]���1�ЭO�6����x��'r��1��+�e}�֮b���,δY#Ṟ�˔���b��S�0��nl&���u�����������M��Pڪ�{N.B�$���˫?��v:�+}E�۸(�*��=�3B�L�fL�h2����gٝm_�֪F�A;��5?=>h(�]�N��_=��U��a8M"�Q;�����w��#I)�r1�p/�N�w�s��3�=��鶆��Pq(���C�U4(z�(�mȕ(���.d�k:�>u�W[��E��'�+�<9Iw�I$���҅�kE�s��sC���Vz���$��5�׌��dD��W���u0�O�HE�yM�d�63Jh����tx4\�����),�|MX�q4�۱�l �) Kc�� ۵g56��4t5�w>�4���r*�iY������LM/�n�������*h��c�1� "��%����$�-�O$LFH��j��u8���20�9�@�^�`�.��S �e0U䇗)���Nu�^@���X��r����
j,7=�~"[�M¬�N����O���=�
Cs��35��u9�HE5�t�N�<��/�i��!9��H�5�!�@P ���v��&��9���e1f
����O�1F��7Qd ��)���aH�� ���D��~j� �KG���pv'IО��^��yKU.���
z4����B'*X
q��V7�c�RW\vin�ZVQ�D�R����i�G�3�؍=9Չ!��G�[���`�p}�Ĭ���x�k�=`����~xw-<lS�cR�Hrgp<e�A6׋��I*�H0�f�s�;�:���a	��"T��״��bʭ �;�b��l���"�L'����\lG;�{�6H����!�����{33_o�sZ�Z������Z�ĆU�_����i���%FP[�uS��`K����o��L�e1~�� 	�A�	�g��|�<����|��gp�u�f���^� ������Q�ɩ�ć}�r_��^V2������� -F�!��v�)e�xU�rTs�s9��#�|�Ct�'�m0r��1�!��y監͵j~�U�� �EQi�C{�d�,�V���&&�2�g�驻��Y$VE�A��HKq�2�(�����+�{9�1��m�s:�0@7����!i�Y�)�[j$�ְ�>؄���	*W�7�!�<qr��1�Ci:�"1`^�>�FWX�i�)ߡ�jKɀ�h�&s��غ�1���E,�TgLX�g����ou�j�e��~���7�;����zar;��wn�X�J2���ޑ����;��]�p=��MaJ��7��U9�=V���A�.Z�����.ĸ�ˢ�|Z�@�x�0��y:UъƦ���"��fo��s����j�v�v�k�����2��
&�����-c?��
X9D<��4/`l
9��ܒ�b\}�vVK�}���\�+e�YC��֊� ��]���NX����Fߢ��L�<\&,�y�ƭ��L�8a?�|����ψ�X����ȃ��p��-��X�؅��|;\�� �8�|��{��]���C7s�O�C�5�ćK�?���uT�-�5��i�9gY\T���E�%���b�������K�d�?9���%�x(���k<��N�s8C�U.RC#��R��=wM%�٩rM��0Ċ��|��so��%�F-��6�O��N6�;K����c�bX��$#H�NF��������ҳ�s&J�˴^����/h�f�_����BYB	�\�!pe\.��R�*����۾�������A\N�h���tn�.��tcU
 M��jھ�>�pt���oȝ@��؉?���E��)?{.� �(p􍅂�� PS���A��-�%�_��h{-G�Ւ7[*��*�VY&雮ٳ�$Q�`I>�|�j�C�\p��O�'e,v�-*iSXeMe������?�y}puj:,'^Z�4�%)~�a?���>��Hu��1�"e�`a���X���m�3������r��"D��2�	�������Am�\N����2QN����vJ
�#&]|f~��������lF��G5i�F��h��،��wr�_jR���]����6���y`��1���������(So����U������]���.ģ�{gM�׸�o�Kc��LL�=��9rtT��ڔ
_�@�����7�7^���m�)����q���ީ��"d�1�9�$�2+�q-|�d�Øm-5�R,��0$cO�՞��*�Gl5r}\��!S
 4�j�T-��	���E�Yl�+����,@�;�$�%e���W�s�S��<�o��[��]�{p�@��K�t���W(�pwh����laq�a��},K�9s��0���6�S��zvBrD`�9:	�Gѫ�ACƙ���H_)FJ;��u��;���x��e�;�k~���	�Y�� %YnJV?l���/K���fw������]B�lE-m8��Ȕ���G��v��xW7�c7ڙ�Gܰ*<Q�&C�#���vC,��!"U -FT7���܄�&�)��%׍���Ӏ:��$�P�� �@E�Y��Q���My�d�i�]��~���5�iy8q�-<��m�ߏI���)�Sړ"�����死O1�����{c+�� �FC�w���q�	��Qه� /*Ўo{9<B>���n�;}�Z]�ӷre����!� �{�6������1}U�N��ƎA���d\���x�_Ѯw�ה�l ���H�=����ZX�$,�Nés��N(��k!,?2��{�zEH<��<UM�����~ދ�ȫ �RyTߠ^:���hM	[�}p���J��z0����m�B`p=�n�z�����1�G0�uś&�\g.����3FN�A���S�d�iəp�l�;�x�q�Ԡ%����ʱhS&)�"P9�q-��� Ϲ�(�Y&P]C9.{(g���o�a��tsD�|��DC���;�9�c	Ãa�!�'�Z@�U�W;�@���pʱi(��e?dC�UG��z�&B���R�~A�UoT�O��X�kd.W�|��-��H�Jj���9��@����%b�Aj�;k��Y
�ր��0H���ekW�^��{�W���Kw����������υ�w��p�t��	�(T�N�y�ٯqU�[������p�2Kն�����Y�J�>M�]�T��U�Sd㌳P�y��r��ZI&a`x=-N������{5<^c�c6��h�����D��7m�uT�RK�&m�L)x�^_Y�!4):9m4TPqf�vJ>�<G)������+b⇑�����Q��juC�s4-��h��+#SՈ�9F��j����la��%�[P��, �t�-7�kZ��EF�t����Bi�r�}R�?R��y��"��j�4e�����Ȫ'	�RA�$w�ء��-H��qd�Ya%���ؕ�`Ҍr�q(�Xb�{�S���M�e���Gϩ�"*$�r|{V�y{��mZI���U�>�|���Q�4O`�_�uZ9ٮ
 9f�S��y�IiG���x�J��Ps�w���6[�4)8�<�>�Y�����Ǻ翫n/n�o�~�u'�p�^�넍Yx���"��������V����y_ʣj����7Z9���$=���R���+��t�L��̻���W�;j����n�c��aGȼ��ma���|���
1`��:*X��	���Q\>b�)�}IsPR�!�Ee�̠��(�v�b��[�Ɋ��ߔ,	6�J���Z��V����W������Ou]�p��
Q[�Q<��A�D����1]�xih�c��f	��A�~�P�� �}`U��lj69�R�&|$�D�TCE�8�:g-=�.��YB��J+����z=�?�j��QC�)N��墈��+�1X�����\٪�Q����.�YN�/,O���s�ѱ�]�pp5-�;���dD�x
|:�a��$�mrn�u[=0O��k��N�iL<���b��Ϣg������ �#˫�Ĕ�I&�q]O}y2�We�F�\W��1K��b�I�)���ux��ނa�K�t(3�������P�R�U_���#����aI.pv���:0�'�a~ �]�am��� ���O��l1[N)��JSe��n�ٔ́�y����ė1��������&������1b�5�����g��	c��U������1^���=���2��k�ŻŐ�k�z�+\U��z]El��F	o��8�䲶P-��	⮭"t��j��9���'�8@�j'��k�X����e�,�S�M��o���:}��;�fҭ/�m͇T|HC��1l5^_�$�f��u�a��1�*��	����v������+��$�:5L��U(p�=�X�1�$/��]O����)����݌"�0�:�h*^:^ ��׺�wt?��6���U��/q�B^:�͚�9{�";}�����g����C��"�`Z�������;mu���X6nĄ�6�D.F���U��S�w�&h��h+'�0��HD�Jח���8��������rL�5{�T���I���Mk�faޔ+�}åC�7W�O�ug
�&�b���+?2E�_�,!�{j�����s�Iݬ׋���io�����t�Dm�ksM�܍:��b�f�o�e��كCk��M�	�C�-���n9�
���H.;ۓ��Û������*b�(	���z���v�R�yv�E���,B�t+DM)xۡE}�'}Y�e#��2����>�������z��� Z���càS;r �|�e-,�9�1��Z���
�C��:F��֩�%��=4&�\ ��/L���E�Ԅ( �e��.��P��lG���g׍��I�Z:ѻ�Hv\T�A�T����ri�HC�Ň��_�j�h�I��S�bd<Ñ�ǡh6Xj��B���p�=<�����#��MB�	҉�}x$��'}j���%z�ܰQa�/T�N��'�2C�l&�ڙ ��^�s#W�|zZɩ{s	��R�(�����g}��X�����'Ū�� !�v��0��n�E�*l���f�%�?�/��w�cz��*�t�����J�כ1��u��kr�ɜk4���$h6� Ωd��6�U(��.Y��%9��̶�
�E#wI���H:C�%+<�գ��>G�-��`�j|��E����ͤl�S��+��D/�w%)�u�z��S�WeՅmq��}�zm9� g�MQA� ���'�B�����ͽ�h��YA��9�y��'o�%����������z"a��G0��lQ���n�#�������(Bϸ�Q�@ػ-��7�"_/"5���(�ܩ�Kx��O哺��2%c#6k����:֍r�>O��iw�4G9x��\H��#8*��#��S��l����侪2���Li�
�V�4k:
^����� �@X�΅!����C1��D{C���g[��� v�U\�Y�Û�28ҭ`S<��V"��~��˸�B���)5w��9iS�[	4_���a�e�m�1bEU#����d	_S:|�V��\0,�J�4�ȿ�w��<zr������'����y��H���̢�q�ß��x/	��8��m��A-p@�)�Ph ��"u=��F��P��S�����[�D���l�;Dbqhvo�P������!&�����L3��ݜ��ϥҕ����W��1��ͯY]�WM;���4/.���3�>��9xB� �qW0��>��>S�Eb���9F"���'����Be�yi�Z�	2E�Z�p�C�����n����*�I�$P��ݲ
�RD���<j��
����;�u5�G���J���J������ڟ�"8$�����ts���K���ˠ[��VQ�W��5������F�I�̈���q�B��ɒGAX�-u�h^�.�Y#~廮.�jW�?�� �{��D����Q��x����L�8%�˩�5��-��ñ�͐�9�9�$��KD5~s�ѣ�;�W�Fc�%J�p�h���wUn�����j�o��IRg#e���J�Q>� �˟A�9>���db���}�ՁL!����5�<��Ɉ)-\�z8�Э�5��Ŏ�����U�%�viY����m��D6�9B�����EhP�A�$粖����w �^�A��ʰ��� SnjyV�iP%�@���k��U��'�?%�A�����UUQe�05q��^��v@~DR!qؚ��.�Sz�m2��Xp\�L�!��1X�dJz�����v��s�h�,���iL�
��lj�6we�X���<�1}��в�)���s���߿v"���u�k1���/;�\�����o0\�DL`A�u��W��]se�0�"�D���^j �3]R4@��yg��)����_�\YL��CMx�i����|��X�*yy6�l��x{57!����W����h�	(�_l�(-JEA^���N�m%�h�o�P��*��ܵ�;��ЅS�b��i����'�in+s^�"�`��0��,���-6�$�.��r�w�k<���=�ʵ<yL�C�=ɦt%Q?E�� �����4�|d�-F����;��"Q���@��0S��b�K�H��؏]%;寢�m��o^��@*ZX c&��f���0�e���+�{����j�챵X�Ѧ�j$j߉�4c�I�f���o�bFo��J�GGu�&NZ��L�z�1���>��!.�9R�?FI�[r�b=N�!j% ����/��3��ŏ|�1��`S�T6���t�b�*�2hIi��!�&VX��-j�S�8|�x��s�^nFf��c{�r泉6 �a�t	��R�V1i��	J��p�P,S�&�'�j��7��^