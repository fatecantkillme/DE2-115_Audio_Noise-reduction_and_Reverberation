��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<E��D1�a��Y��0�q�9,���;2		�<)��`k��84�`Yr���o���*�֊:"�ل��/�Ps�tߛ;@�'2d��z!+t,]cL�TH_>�3ۙv��i��LgUz �22�⯸:�]�-��%6���͛��9¾\J��)�')����Z���>'§�����Zt��K`��e+#�ʏ�ܑ#�@�Ia�ք�Fm�QK�̆�FB����㉞���]!3����kMrZđ��E[��(�BK�}{�b�-��D$ܾJ>�����4]4�<�R����45����}c\������^�iUK��ϧ%��2�ֳ��n�+ⴿ9�}�_�O ����}��|j��#U�wX��ⳳn���GXU��+86+�M8�	0��T�#SD���k-D�i��
d̏vX9���E��c«ۥ�+{�3�#L��`;��t.8�[8nK�<�Q��ܕ+cZ3�)��H5�tY;1����5�\J����~4�Hx��bn�9�f��2�n#�l��-F˘�E�i�:r������n7h)��@���`�Qx��n �&�=z[����"Cԓ.o`�$1����{�=p[(���k�#��C�aC��;O-�����h�Ԧ�wDs�HQ�)m�;W�),x��iѣ'�
�ҹ�
�b%�W��C
B�:�]���_�-E�-�|��:�ߵ���<�]� ���K��)��a�s+a���Hc�Pw��M����GO�����j����d րԖVH��$���}��Y��E����YAN��7�^@�`�9�.��S ̊���i��醺!X0h�vf���y1�j4'{�֞��aa����k�o=�Ȍ�n�ٕV��M��*���K�����m�T�N̘FP�����	�W����v3O/8�z��fij ���t�`�iny��-�3z�z`C�p!q�n�:�^�-<1m�h��a6,Y�	.�V�lļ_l�y���q���:�*@� ��?���W8Z�@��;%���pQ݂{�Qih:�d |-j�@�B"��Q�ݚ���-iM4���p�a Ɉ8 0�]`a���^ʠ�"`�}x^���\�䆭ȏ(Ӄ�.�֮v����Y�P�����cU����O���8:�^�E8U�_������'�'W�/Z̢����؍�@�e���D>D_&��*�g�{l!�B�BU�[iv�ut������ƃSմ�#4덐��XMW;�j��;G�T�˝l�qβ�!d`8Qy�%Q^iL��6t����l��yҜ���g�x|�ۄ`*@ˉ�������<��
��S��f�A�3Y1�Oi�2k"2 װ��*��kW��lk��
�D7��	Աt8��濶���g���	L�@r�Rl�R$�&�c������0�	�y�����LXq5l�P�K^�	Ĭ�`i�x�=M��y�s�����h�.V'N���>[_Bci$��Gs.�%�-n��#��� c6�5��.v�e�9R�
X�S�=q[!���ݑ7ZV:�bu7y��0�=� ��C��
d@��7e5���~Ȯ�u�����H�'x'5��{��4=?�W���=�!��9pƕ�VP{�>Qƚ�u�D��*��d�5g� ��H��~�޲;�Dj]��66Z�qh��mR|ݮz#{i��w��D� �S0�,?4��1��YX+h�QC5=*���4Zy��Sb����Oc��ҍ(H����|\�N��_��.��.�>z���vJ��|��C�d��S��2���xC�б�`#�>��]��gr0��q+�Ě=?b�(wm�_��%h���Ag&�&p���+Er$�'�j.mJ��bw�΀�z_�����}�J5�>?��,��$f�x[�Qp�6�Ȋ,�Z�Bfm[/[�˧ B<ii��3���a��l��v���̴ՙCz�^`��Ak��w6E���Y�u�`��q�E}%��GI�10s�}����ȋkk�M!��^
lV��G���rSxݗ�RI��$	���w��G��R�u+�l��X/�yjpM1S4n��	0D�a��0'%��,���� 0�o��{�0�^�?<A����-W�Xr�%�w�<7Mݯq.����B
���z���L�G�sj7u��;R��}�W��W�D�y���yև
������$4�k�9`�ȇ	T���2�������=T�-�#�3����õ2@#��aaʂ��}���@�����z�LlL��X,k=|N������VQ�x�D>�V�BMnt̀�6��r����T�S�%���')I�#�t�����7��m��*4�V4�/`�ca����JL��j��\^%ǟH�G���&IG��A��#3��J���6>� �5�p�s�q�3��{>�i�	���O�.��r�_�-��i���V��.+�hSh[�Sv\�v����]�j�Y�۫��V ��C"�7/�{o��}��@릤����a
y���S�O�����ԍ4f���_S���~�D�8<��S�!t��<n�T���}G.�C�����2��f���A;%/Ԙ�KYd�R_���[�4�fU�d����B��� 2f{�Qߊ���1��X2�n���=_sz�1�^�!S+bST^�L�]�3Ǒ����V��H2�헐9_̙���q�uX�^դi�w��z��޾�#Ar��c�,��6�V呖��P�'��Zw�c<�O�	��5���SXr��?=���w���ы6�m������dB~&n�\B`�E ��{�Ǵ�����تլ`�u��Ќ@'�O�Χ�d��QW�47N����ݺ�W�ahα=�2T�M��Gǡ[�����'?��𾯃{����-#XIC�9�����,���i\�@�&�5�%	
-B�`�Yn��;U{zo ?���1t��3@#tUb�+�:le�տP��_s5�|.�/h7)aMI��#��K?���^#w{g9,��Z��p�H鳧dHh^u��71z�&]�ηB�M���M<ޯ�D���P�����������y���@�Q<ax�<�o=�(tީ�����r<��$=
�h7�hI����E��0�~KaT�}��f~�鼵�0�}@�����Q�~ʊ@���4x�gCY�R=0�:�ad�+p��k�Q�몚�9)��ɨ�<Xn��<騹��#Q�m	�؉(��{�G����5h�>�|\H3�G�A�-%�ID1�9�rD�h"I�(ĥ#~JR�H�Bka�A��/���ˑ8�Y�ȖN\��U`���?52#�3�}`�s�ܫcb�w�NsZ��Q��T�;�є`j-�U��̊�����	hbtی�LVn��� ��{Pm�7�!�6�o�i3p4���ai�},a=��)J.���Y|Ð��{3��\��̃°�U��&M���e6n�sQ��<(d�{g;٪}��bc�n� ,���}:�����\XX,@�b�0�*v�_I �R��v�-�	?%3F��3^G�;��i�_h%����4H��������9� M�:��G��*�FN@��裼�'���g�B����w�L��ҍL"6��iL�vP�J{r"*k{23��`U,
��u�e�u�I�#�Epx�ϘV��� x5׊���ø�|��ۆ�;��B,�|�K��oyQ������F
����'Ɲ�҇�mD�2��CE��D�߿��*"rЪ��=!SV>z��zSHP���&�[X΂x�5�3�k�u�2;��ۛ�#^��)��<�6�Ei���c8�OZa�c���~�B����bG�]�v"oij����2�BX>��Nrs�WS��r�C���|��v*b}8��1ZpUHW����N��u坹��'gz{(R���}:~�����J��������D�g)]�'���a�s��I��)�)U۔����,-��<��oढ��
h�P}V"ćN4i����R�s��-}�����^�XLI
��?�^���\����`�/�ڵ뚿X�7��#�89��:jCdg��k�%�ga��w�>Av�&K@V�;h����?���pITU1Gh*�
X@vS����h5 ?)���Ѻ�7����Օ�h�X9��O�N;�a�x�5`$ Nl��dqD��ީ�u�8���-�f�ўh�ǻ$ (�V	YcW���;�Z�s���k�BJfa���͇h�@W\�����wE%���*��du����(`�>_td�L?�_k�=�6?�E��K8ȵ8鯸7��V�_���)}�-�0l�"`1c��K^�q�����gvn�56������`�����N0\Dj_7;	c��|f�w���3)�E�|gz;	8?	tO��!�#�h[�a��W�M�-	�L���g��f=�q)M7����vʽ.��T!놝)�1�?��!e��li��gv��8o��]z�T2_H��G=ډ���O?s��dj ����A��~V�1Q�C'4��׽]��ׄ]Q��ˉ�+��_߮��[m��Y9�=p�p���9u+>۳7���ͷ��El�ȸ��x�]7��W�5������,^+��0%�n�&e
�ո7W�m�z�C�Ɪ�7�,�MN��B��}��N�yaI�"w�wX�����4�V35��,��8���f"�uS7�]/� �'�ǂsA��S��5�����X�目����U�s��o���
:��:u�P��>���T�0�8�`�7"H�dǍ��p���>A��Ѧ�S���&}���V�ɔ�C���]�����?����]����K��Ɔ��c��q9a-`�>��$ѻ���]	Yr�1�VJ�X������43���29�$��`fckc�)��u����`�5j�2o�B���g�+�v:�Ȭ�p�jU
y@ t>�Sǹs��D��:���l�bwrJ7õC��t�1p5u!��͵͖+�����ӟ�	�`�8�`�P����{���m�0�v�q*o�gil� -� �[̷�b���a�r���.�tBZڞ���I�1�~oZ� n_(պm��O�I^^5��c8�%Jv^���,X/����+��
�9?}{���eJ;(�n��S�ʲ0A�TqY�����D��yc�R2IiB���_ I$NE䳭3x��#��s����P��Ks�MX"�7Jո���NY7i�y��4�#�4gMny�����5�CxG%-��s�"U�_�d<@́�"�[�����deR�����2�o���)��$ș-[��^m	c4��CVv��Um����b�aD�����赻�7jH�2���ޭ]�����Ŀ�E%}<�!���`A]���D�f���#D	ň�E�=��\	 �C�J�R��V�8�Q��7�D	yxw��aAÕ^���6F�hM��QX�zm�d�g�ua��2<�e���o>3��%�0��ejI/:Wehi ��?����{��%�q�t��c���? >�bNÄP�Bv����}ԓ��P��_A�| ٙl�a/i~��A��U=��9�T�r����3D��Dm�$w��ˑd��#4��"N�
XNX���Gb(�O�a��z�U��:s}"�}����j�=%e?�/ũ4IP3��	���wi�{�&�EP��p�4<�����KI0�n���-_���u�(6��gD%h���?se��h[��q�Kl�d�\}�C[��!�_�8w3�?3����5z��8�[Wd��xR�
�'�uj�'���]����3�@�f����A���3 +0��mt�]F��q�{�B����e��:���h]N����6x״���(�&RC�_�
?W��N�w������*J�j;���Y�ޥ�� ��M�c,���s$�p��<���N�=F�j��}1�ʿ,S�fO
��B�z�8�g���|�+IƸx<'[g��i�@�-�&$��MTW���3`.�W�c���?�x�,l�`k����`����-���� u�� d��x^ЖMߺNJ�R/	<��w���5���?Z��PTk�U-��0�4LM(��:��S�%I4��m�-'��W���%����IC���%�0g���k$$?�P� *�B�|%�5\�>%�BdD&=*m��0v��^{����0SM+Kg.�T��fw∖`r�M��6����E�"a��Q8P	L�k֙<<������Ʋ�8�E!+EԷ4����OM����e�i����*n+��m����,���a7�y"��r|W͹�oD�0_��=�nr`'M��t�.�E����بCJ�u��ʆm�m0���]ϚVT��F��j����>��C!��ryǳEw�h�|B��7Nޒ	�����*63^&^��7��U�].7��
���+͙ٚ�"S�������,ue��4��Z |'�U��3���r;�cѯ��Qz=Z� 9���$M�+~W0��c+����7q���!G5 '^�%CM@�q���E�7M��<�5ni�O����?��W���0�/B��oQ�}�_��,ڻ�e�J�Le	�Ex�P��r��7�¶���-�dФ�@N�߬3q'h����h�x�"V��q��i���Ԣ���AN��t�B��Λ(���wʆԃ�
n|գ�l��.?��_a+��;�[&����6��<�����]&��jlma!�g?G���ՠK2$M o��/���)R�4o+�A��種%V=����q�c��\y>���#l�Y���$WZ�,
m�B��[pl~���xl�|�D�����&s�s:1���w�h&<��p��7��\lбv�'�b
�I�e�mH���F[N��������SA��^C�2��G�Ch>A]Q_l��bt��<=���f�|��7���^
+2�n��g��}c���]�W�{�t�����5pz�@�W�_��������S��J4��n�ԱGOD��7!�eG0,"�o���D}!5����U�Δ���Vr���DRg�[x�eE�|<���w�u��o��JɋQ��4�v0�<2�05ȷ��7�$E��,��^9����6^��N�A3'�>��cBE��Й�n����f���C_5���#�i��h�������tu��4��F������Tɖ��
υ�����^Q��~MS��[�³|@�z�%iDe��U���;�c�F��5�ԡ�CJ>w!��^�2u/���NYx��j�v������k|Y�z"0��1�Uz�*�$����@\�kU�Y+1�9��6�f?��c�����f�|�j @J��{���lZ����������Ƀ�q�L[�Uf��9���۲	�iƴ[Ӽ�uLlC=t��Jx���FL��~Б��z`��J�x�w x2�2��d�UUY�ܪ܇<٪�`���Cڃ�G����������^A�'LBe�Pn��&7D֯"WkWP��XK�C)����<���E�|����*�͙�:�����ɏ	.X�r7��뎳N����a�cТ �i�E��g�����Z;�xTQ�
]��2��oǉ������b�?�����B��XrA�)}�t4Ӑ��x�wp_ъ!�>+�Q�խ�s�=Ϲk�x,g�	D�ۭ�Gᒚ��RH��R���+x�k$�؍>N�JBX�?��`=�rk�1��ܢ���E�{�z,������	fE���*�
n럫��5)�J�^~WZrG��1 CcŶ�A�,����혔�<���&�]��8��o@+N4��(��A��/:���@��S�@���2���ji+��y��u��#�F�)By �cd���w����mV��;sa��zJ]5�����9w��=<���Ԉv���M�2��ܨ9����*��bٕ�
�ڈ
P/����e�r�Wv�j�~��[ Y���9��)T�I�È��pR�Ih>4����YS�qgj�msb��%�ʀ/�?A;�`�[YX<Ҹ���>���A��ܪNq-[V���{��_�����*�nF�� L�7@M�W���XfWDs:�!7�i.�b��	���Ơ��>��8���c��ujKuz ½�G�\����ʻ*cW���x\8��#3���m�]X��� ��L{���{;k������!�B���%�Q���9Ao�����΢U�
<�!���.���e&R��x�S�iF(oW��
���*{�֣�o]�6�d�}iEЗ/znfǔ!�oq����Y���v��(G�mn�����ǂ9�[Ae�s�F �ӣŐB�X�-~��6*���-��c$Ce�=d&ܿj����o�y�z^�L�n�/K��(�k��+ß�<��:��uoQbMg�l�/̷T�Q5R��w����x�C&ǣ�M}3Z�od�}b�KʯȞ-a����U���^���E����%\yR^�x�t��"MC��a��m{�iHE��\TO���c�ժi����dg��"�b2|�BP*���N�6�䬺K��w/��J�%��Q��l�AOry֑�6��=�� ��#������ira�f䷁8��?\��w{Y�)�uq����~q�,G�"��[9Za��b�U�0�=z�ppl��)7R�J��G��yq���ߓA'�L��d�$�F,�q!��O�G�9�/��� �۳,!XԐ�,�W �L���7�4f����l�-^~?")e�o�tҚ�޼�(��	�� C�⎫!7{��3}�y�=��ɘ��ac��cB�1X2��o�����������Φ
NC�,&d�e�e�Z {��{5���	 �G#;n.ZPإS/��	`L��L�`�o].V��"������M�<�y6V�X��l[=��. 	���S7�3�Rh?��t<����k���_4-���đ��d;�rM��R��EX���O���^`68G%����@X����}
Gh*�D�gT�����4��ũz�}���"�>B����o�p�*:���)�'2�D�r��� dH2����@�/��f����r�Z�c��j�CUP��H6)������Z�%�D��43��O����Y�ǸZ4�Q��V�GK��У�����1q�S�N����A!v@R����2&š�h
��89O������-����hVP3�,gT�	R�K8���L�� �L+2���U��{���ǅ���V�S{��H��	.�/wg���damC�:�.�~a��B��������=��\�y9qiA��e��>!�aN�N�.�[v���yT	�f�eZԥu�㴤�b�!nG�]��`�+��K�dP�c%�>8�Ԡ�M"=�Z���K�+X{���j�oLE�d���x=��7wO��<��G����Kw�����e_��ލ
N��X{1b��}�Ov]���4�雸la��Hsn-�P���5�&���m#�f����s(,���^�&7�������,�A9��S�RVq��̃�7����Ѹ��a��7[
�I�l��*$j
T
s��O���C��x�>ă$c��q�R���6�%�8�@m�Yo����iB�xZ#�dY�E��7���[��o�顛�'4P����nk�1���3|�1�G/�}��b��)��G��M%x��P������+qh��� �#��ù�z;�l���).�C��݃\*KK�d���4��fR�y<��W���]��Wj81iO[w��3�<�i=
��%nX%��լ��"oO�X7(|�2���9����2�74���,ax��L������$�]�$�c�b+t�0�����չ���Jt��[2�v�1y��]Z߇²9��O�v�cQ��ɥU�OE�
��n>�,񣸲^��z#r�{��X�t'�D����<�\(���l��f$���E7D�g����O)&�~S�׹�6�- 4CJs���r�eJ/��
�����r�o(��Sϛd*�5fDT��{���j z������W46����a:�J`�#�~-�
-d��ZO�0}ҝOGF���o���n&��Iz�!�V5�WK�������:�����%�d�"%���/��Y	�s�q� ����X]mO0��cam)?��(�|Z��
�Ur�����;)������g��U_F/�l�n2�C�*�߇K�-�3�+��{P���8��'g�	@��m�@����
�r�,k�/'P�
�9SCWx�d��b�hS(3胇jD�~F�c�GR�gZ�%!b����	(�ю@��-�Ϯ�:�Z��sIە�PJ�ɾ�/�ro�:�?�&�骕���B�s��W�+u]���҃�3`+�@[>�޵���?��A���)�bS����^K����I�������/�R�N;\A��h��&���S4�(G�g�e�)�CT�J?2+�M�}&��g��j)a�A￼�g�^�>d�0�@���U������!��Qj��X�����t�2!�$cq6<"z�p��vk+��ԥ����{u�-$I1��h���p��2Q7��'�z;��uw~cK�*E��i�`���