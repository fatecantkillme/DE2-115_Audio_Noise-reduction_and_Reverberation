��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<sv'-e��4���-i��Z=���?O��q~���rt�u��25^eW�g� ,x P���������ƀ�^_��i��⋞^� �e|����;n4w��xl�/�ղCZ��q=t�@��?���NkGs�P�^�m��-�5��U�d�6=a ��F-=ʦl`��6 ���4�^kB=��Is�fæ�_R�Q�#���g5![����A�'i+	B�a��,��D�n`o�\&\G& ��ϯyB� B$q�P��Ra�Ȗ���j!D���~.����":��i�b�'01���1��N�a7�ȅ4��T4T�艵�ү��Kb���\�䰮F&(`��V~_3[f��t 'j���Ծ�;�7�C�s�"w.���	md"���ߠ���Rղ�V�^L�|�XNZ�e��ߧ{�@���D�.�g87ۿ��*���C�"(�RNQo�g�=q':ҳ�������0�4� ɑ��8<%��~�����*�}�>��_[�L�	4�@}Ne"VL�cIͩS�=��ޫU��%\�Z��A�ރ�Ȣ���lZx��I�*�͟�����O~�u]C�nǄ
p���V����d�rgܢ�z�H��2�I:w2oe�"�w�:�λ�k'iUg9{b��L��VP��%�ͱ��?�L �f�T��-ueq3Ϡ��J#�;�|B6�[��'�.���7�����^۫�0�J�- ��X��p��{���n�{d�C�S,g��q��P��+�Ym���ҿaruǟ+2 9UK��Ӓ��(�!!�v�N���G�~�k���<5�Ȳ�j3	�;\��S%�������Sڠ��/1��,���Ub���H�^e]RS؂��%I�+�5(~8aO
۞�p ������/�gI���O�<��ȁUU��qp��-a�H&QˇQ�k�n��y��3�r]�vrZc�]��-��H���BkJ�6������>٭_�!����+^��s'?��0�[<M�f�橅Q�(f�'�� �L8��U3c�Pg��X�]�� X�l����ۃΑ�ݡ�j�Y4�4�� �An�ؕ|�9�w�siοz	"��![��,ʾ��x��j�}�s@��N`ȫ�-����_��˚���]�ǒ/�zO���T�}�0�̈́�j9'�5OG�c�&�7�2.%"v����	h�v�Z%����{�7�% 2�<ReB�B��j�����D�oBd��e���))�)Q���|+��JS3����Tx�=����8۪|�p1n�e:� �AҸ�	H�g��3��QW��Cec�=����x�B!|FE��W=���.�Q����W��kN��l��z���;����Z�������C�=B�Vy�bG���«���r���~��7��X�:�	�);��Yym�7�Y;D-�-}:�(���)uS91��ncX�Ax�y�c�<�ْ�����R��?��r�� �[��{ʨ`��q�I:|�����5�*�_%@#c8�rI��d\�Z��9�Ą�>�>�m�X�I9�LR�`��2�&���1�U4�g�INv�-q��l��y���y�`�}-�w�6�&f���J�/���s���h~��V65�|J�{G���3�~g
�;�.<w�`-8��a�S$�J|Xw���2V� TX�x�[,f��Pot
���X� �Ű*-L�Mfe����c���(��
%��&ҔA��n�V��T���1��BOǀ��" �Eq�������8�S��)�ɫ�K$��$��<���n��9gM$�f�"@j�/����uVԺ��I���!�-�GI#l�w��{�@�V��."���+Tp��!ZP����["R���,��ܲc�8=&�z�,�M>�A�ϫ�j ]mc ٺ	��ix�g���b��IY}P�Q�I�X���TK���mP��Ԋ&�!���!zI{���/���ז���atZ�h9U[~�kW �f����q��� �[�zXz��r"���(,�K�r7�@��_䄖�W����g���}gU�t �V�Y(��H���r#כc{����������~7
���857�
�>�xf	�o���	��?��y-[5���t)M? oaO�x�r4]`���:����C�O�r�"RΌ�te�:r/��g4< �͆U'�)2�mRٲ������kA��p=BLY�24؏E��i�&?&9���}m�E����R2�d�)¦M�u�����Q�
�g��5
ɪ�v�`�F<\�:5�|�_��`����s����+�vfE�L����x�"�ƨ�ӟ4q�r\7R�r��{&H�N��x����"�C8���۪(۹0T�u��[˯��˞��
I e˵�lO��8h�h^���UA;�������ù�9�*e��>�i�� �r����&,�F�v+��Ř�v��a�W<�L������a��-��O	3�T�������~!��/�ͮ�����6TާEp��6��	Y$�c�c��r�B����̙�g�AQ7ڔ*���&�)��(K���!�Y��^��<~8�Kڤ��!G���-�&Q&H�nN��_"�W����\ߓ��:�L3z˫�|Z����_+�l'a�RV0S3���v��-�]�9�I0�W ��P�0���*
��ȅ�=��x@�zO|���p��I4`j��7���l}Y�
E-UެDw�%� :���X�(`��g��iB7��`��ꅾZ�\-|9�;b�ʹVG�H�.NJ����	C����,W�����{��-����	aRE�1�ͽTd@H��;�s]��li���ɴ�c8(�
�Kp��h�b�:۹_0�����"����h�;�)<5�����5]N��w�Ōfw�,aݶ��9��Tڡo�sa���N&�ĵ�Y�"<X�1NH���Ml_NU/m���}���OĖEgk����v  ��~C����">�f����):߼��
Z-�v\ஷ<O�ڊHo�c!�M���3&�tMW������U�f��K�>�>�|T�b���e"����ѰeH��A�Kլ��Ug[mRU��)uӱ�T�)�e�2fr3־w���_�H��/�U�?N+
�Ś�g�ا���W�`���
������㭮�Gь{�t�F�C퐕
��,��x_C!�b��tm~gm!:��m�iV��yht����4��8���}n�L�9#�`&I���!V� �]-(D ��~Ȯ����]�O.?rI��VF^37�Jʌ7�*���o �N�{���9��UN&���u��ޯ$?��C�k�lF	�!WX$�����"]B�g��a[.x�o��Ʊl	H�D@�[B��"���e5�������ykd�:��S�^4f�,�@OT}�~oԽ|�l�N��BVysj� ��w�o��ǌ���"'���`�)a���cdr-I�_+]I�Jd`6��!,���~�[����&�!,F� Cb�\�ݤ3�	��g�G[�&��5*)���:�{+7Z�Xr��!^�b�rs朇�� ����� E���Pcd^�ɞOZ%��m�r��䯘���C\1�%���q�?:��e���'�$m�-?3�m:���H��.���3���.�WMk+��9ĠLl�aP
���_��ܕ��p��L�s�&!4�tf��W�2�	b>\�޾c�'،MWQ����%����S����+�p�����Ȓ�C�/�%W�d]���t�M1��k�v������|s���2�U7c���5R+џ;R�Gm1{7С?�pu����L(��������U<F���h�z�ؙ[0��%��I�9��7��me��}���^!6��0�w���;X���L�)�D��͡���V��ޠ������x�����^a.�ߔ<��P��e�h ��{s�
��T$�vq�g�	����#=W4��]f���mϑNo�+v�!ޛ4a���MB�Y��$tZ{lc-_!�*��_͍�>����d�����/�k�.�#a#�Li�V�	B
x	���V��.�.�Gƭo �*� �ǜ�n�2�k��������l;�[�3�F�������$<L�3� hQI��|q5p0�6Ջ���Ն���1H�a�/�Y��������v3�M����[_R>�A��>��v�S-g����]�r�꺪� �1�ٜ�<���O{!��w�񵓷AE���pq������,cl�x�8����Dk�缱݃�ա����6]�y��y���