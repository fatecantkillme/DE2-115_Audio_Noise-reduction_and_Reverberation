��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv {d��ށW�\���k�(8Ȍ_"D� ��x��k!��E�$��Ho5h.ԋ�Tt�"z�	�˃ ����2a�)������C���V$��#�`�R�V��"y͆����;�3��e߫�3���Oz�|3i(��=��l�H�5��5�YbB��f�1=#��h�	�8<C9<��	�~Y?q8=�Lw�0�$N"'������g�%��*rKۧr�8'G��_���V2�8��4�~	���+��K/�x���ңM�]���c�Ku2!nѻ��"�y�}4�}���n��*�V/X�G?�Ѽ��/L�d���4���/`�>#0��T61��f�<���R��Z��,4�dOORF̕�������%��n�nR�P%,�~c+8�QL7EV�@\�h������S����j����Uo�b�8�f�GJ]�z)��:��#� �����? \��S6��5�+%�(ʫ~���$5򬓭|� �$E�{�����>���'3h���f��o�M^�j�rub��I�X�6���t��@�{V��[D�<�����\=X���&���k�l�� ˴���Ms�nL�%5��J���Ƀ�S(�;΄�'�ۭd�PS$C���Y_ŵ�G���{��"�%D�8�	�#�������0�D������=ی�#������yy�>�- 0��h���Kȱn�a�o�Џk�k���ݧh� &i���@5� ��f���6����w�	��S�^݇C���4�C1r�E�`�"\���ȳX�RՎ�v�~]��Sj���{IW��	��VǑg����iut��5��xv���DF�Gϋ�ɛ��$�1��~�lԑ��+ �f�j8ԭ�=rDF���s�>^)/-v?zob}9������F!&���\��v#�����,���P��y�z�%�8�l�8��i���-���܈.k]dr��uַ�X򠛮)iP�bF�*��[zs���%���Onc`������ˋK8�Ԅ*��N5����_4����̅��U�Jb1}�+hSs��v?�����RCT4�\�vI��A�����sXt�&k�L�ҟiz<1����1�
�`+K����;�/ZMٝ�7٭��rAΏ��	��d��{Gd7�)�� o����'�C�t������])c�5q�cZ zq�Й��,	�m4l/��x�t�׽������?��c��E?��{R�a"|�R��S #��l� �Ԅ�s�b^>E	4�As����`#��M�Y�)5��qj���L4��k���cH
��2�?mѱ3Q��#@lE?�\��f�Oe��ۘ�VG�b�:)�ܭTGꞀ�د)����&T�'c��=l�H��2~�� T�w�Z��S�U�{)�������������>�2ls�{M��#y@��L�t-:�v�uJu62���T-�}:o]{ʣ��̩���D2��[��D�^����1�sVáΔ$s�l�7?[yqF��ǥWvU�S~�1��k�I���C�|��[� dl����7ƹH���p���q�D+<n���h�D�KT<e�v��QL�R6 I$����Y�f�ې���.ΐK��1���a/�������a���U=�`vO����t�z�:�P��2��7��"cţ:i�-|� ����NH����<$E��u�t>W��v�-�.��K2xEq��s�Ud�f[���vd�1�e0����	t����C���u���**J����'��ع���1���'h~�s$-,#��cE©��0�v8�ҩt���sT�:�,���OwDK,�FБ�p��MHl��`:�F��5�z��5h?�"�@n����q��7��/�2���(�p�w���C2��cGf��F c��ds9%�j�JE��f��Y+l��`�:�u���q���]�*�4^��[0h�|a^��O˅�~�S�M�����E	QYTbaj���}aeğ��d���a��� xb�������q�C�b��f�V�f)dF_��v�]nO-��:�Ќ{�(A�~��J*�*4�H˝����5U;�WΨ	E�bP�_��?��v}p ՙ4���c 6�%��U;���LF�[ t��uDgRZ�%P��쳂{�𽆿�bXJ�%ǌ_1�D�̱��VIW�
9�S}��^��]#L{��˨��ѻ�#B&:� X*�����j�Ϝ��S�}����IG���s·Y�Mnj�I�I��(~�öb�%���
Q� �8�v�����d[V��iy��0v���Iq$���"�_���1�����bq����N���+\:"N��=�})�m�<�g�	+��jp�s_n����..Ar�s������*�Ҕ�A��_!`N��Jϟ��nCb$�����AE9�㨾GR�m-:��[���b����[T�)�!P>ɣC�K�Na�*;_#��\��n"��Z� nn�c���c=���ᶖDO�n!��U!��	c[uH���!'��`�昸ke�ĺ/��[����?��DވY��D`/�H,��.�*�G�jd%Xmi� c,1����
/�%Z��]���c!��8�~�� ��i���ma�2~m�����&�&��G�6� �6b]�gfm���4$(?Q�^-�I�������C��ak�ouƽ�J��s��jCaPք)�o:)��.�5�wXV+ۢT�
�y��G���F��qǮ
2;��Wah�0C]���]�M-e����ݪ�m����I�V���ĉA�Q���Cihe���Z�K�_s��JOlJ�1���OVD���QC�K�ZZ����`��G�4S�w���$O�Ҝ��!̓r�Rl��q�2��չ���Qvr�^D
V�V��ryS���戻>Q������0>)��-4��	�`�O�m�-�N����M��t����t�t$~��Ɖ��zuۃ<q�u���'%��#�c»�Rd��K(�����_oE�ޛ8�%�����1��i������Q��3��[h�0e}{�Z��rC�;n)i����?#��>���B"��8�<�"�9���[�Kʤ6M9T�"�Tk"EK{q���"�L8�k߇&�DW@W�!<�'!��
�ꠋ��>����9�������A<�[���A��u�|�m��c��V�+�����+�?a��kw�#��6 �� X/(mU�׷X�T�T��&PXx�&3�W�g�8ZЌ5d���*^<Jb����Œ"�ݖD�����c�ގ�uV�vE�K���FO/x���i�3�t�Z�t�̺��`�� �J��>�# ������K��Ir/mT�y�2��\R!DAY6���҇�9����i��@��h���J��:1�nm5���c�,(^?��AJ��TyN0��Zl�TY�Q���rb�;p�5�����rK����[��d#k���Ht
�ڊ�Ôz�����n�ҍ���5"��!X��y;:)FE)�%d1?$"�~y����g��ل�{$^p���-��4��HOrQ���j�����XL8�~���ms�jA�TO&�� ���#⤑�&�����rb|�Np���A�bqOBM�⠊>~�j�i��d��2���l�Y���*uG�vŘp<�MX1�,���;�:�zQi�AT�k���e����<I$�c]���Vko���	���5� 
	�x͵/u��e%_�G����2�=/�ߴ��<-ƶsN�ZT� ���sS%|��hɶ0:}�Z���m>E �r~7��I!�"t *����� ���lr#�܂��W'�������<D�ð��"��P�@��ң�Z~�j�.U���q@◛�0]����WO��7I�XBo>��*Mr�^�\G�ps�P�rr���	&��h� G\~��N�[ <WC�t�eZP �͑j�+�b�g���Q��[!ů�G�8�შD̘��|^��QbFe&�8�Ź>�4��W.vB��z��I�v������������(�t(��z썹��,�7��o�(^6�J*��Z\��ӯ�_�5U�O\K�а׼�X�_�9���o7x7���evv4�|���
�)��a�mF3�<���d�Ӣ���j��s��+*R �c��Y�e��s=S%3��ОN9_c77��6#L�9��*̇{ܳN��Ҙ����`���ҭ�:�ڲUz�N�~N檈cc�.th�~��@��$��	Ёۇ��;2�3�G��+XG�\G��kN�O��B��I�n9��>�e���m��
���A)+&i������C���u	������q�RF�0 ~!�,S ����߁���55;ڐ�5�Ɗ׭��ӪMM�kBZuNG�҄��J�0�Ƣ0�6=6�}�FG�����i�iS�=qL0WY��0J�pӵ���S�ż�+TrR�ۆҐ\6���,��_Ʈ_�Nȗ���y�y��8�uCCW&o��z�*,��ykZ��m���8�7�_�o��.�R�G��.�F�zlQ�}^��YKNrN����4 |k�b��jNO��Z0b�,�L��P���1�?=���\%S�i������n}_�..��҉�>�	���$]�,��t�	�Ƀ;�L%�Ʊ�r6E#E�x�/�P�.�b�S��m�Y`~��N���U�S#p�gd��>${�
����9	GΣ�z�,��шn6X�wkMI��8��Y���-��x0XcĢ�lV����uU���KP�&+������������v��+7rPJ�|���n�udv��2 ����K~N�@3���� u�Vo)\��j"�9Xf��?����}��Ĩ��SIw��R��m5?̋��o?����L2}Řf��U����t��m�6�@�A����佪%�,"��� m��<۰+��LS >Ɨ�P��k��(yY4�lD��9�ս����DK�A���=P d���Z�K1��5H�PRW1f�z�7ұQq<W�L;�@
����WŇs'xLh����#BF홌愈�h�*R�|Nc����2'h��`A��1��|za�0�ʇ�>�􂞑��T���b�/��ٿ�_G���^͂A���i�^�(af9:��yIߦ����n<���[_��S@rs�6!�_$@4�4�3Q4������wOb��a����r�0i�=����T.(�]r� +X^����(T�aJ��B��UʒE<G9'�	����~<�������;y��nL}��p����y���D�#���ĔZ[�ҞF���Umѻz���6��[�Vbz�8&���6#ypԄ��XK�xͦ�æ�o�Y67��i��;�����+��P�:ԀҒe�T1G�>�Ϝ��[TTp��_�gd�;���Oo��ܰ�[�[��>卥��E���-��R7��Сd����+��G=��� �T��,���D����@3���Xr. a��yPqU�6ɓ7{
�>�0���v��WV�Ga�����U�P�&v�4%�����T/�%��E|�"i�}UZ��#�qxp�?���ï�>���m�D��2I��l�H?�7i��`��D�x�Ļ��v��%���]�����`������?�,S<Ȱ9�c�U���/��k�l|�z�ޏ���俺B����1H)P��b���wg,�tB�=K�RSć��k{��BU\���2ٿ?��"�?�)M˄����u����VbnNr�[���Y�ɽjZT�S�UB�z��s�#�BM��m��$hֳ@1T+��}��
���_G<�C2y�ո����)����
�����^�/E���w'���b���"YM�!���${1T��NN�>�8n&��;�'���y,��A��gc���Kd�e���D�>��9sgױ��{��ӭ$}`ej˄��-~`+:�o]S��AM�ᮮH:��9���m'~\G�}sn�������JP��N%Ԟ�"r����:�� �˅�O��h����чb�FƋ�~1W�_M�	���λ�[�؛�(��&]`������gsE~�:�w5�vL����G�$my;J���$��M��x:q&ݨ�/,�g��xM=;$��ޥ�~��UU��ҎH�S�6ݺ�H�c���B�4������޷�H�`!߀$�>S��:� �MېScė�~��{� �w�����%dq��D3���9A	��D���bc����o�j�K뚽<�Ѿ��R ����p:Z1�D��(��npĸwț(5� ?�-���ᾩ�:�5s/�-2'�s���٣xm����*ݠ`]��ހ� 5U@�g16T��"2��hڥxۄ$�`ĝH��W��A�|
�Ju%��f�Qݔ����0X�h��v|Ұ��n�9P6ʃ@�"}�nbv��t@���o��j��e���+8a����'3����v��98�d�*.Z��4��B��O0��Z��晖G	�^bQJ�F�wI"PC�m��e�l%Xn����X)�5�]��EVF��
|&�!QK��ҡ�d����zƥ{<m��N��B� �3�꾕�z3�b��%"�dL��-��A]֥K�c��v�#jY�W|����B����Kֽ�o^���hK��~���R5�(��O��7��!�4�S�T�$��>_�V�����u���Ԋ�;���vH�����H$~mSE��H����-�թ?�4��soO,�S��z0�[¤�#�?_�P�(��zg�J?Tx@GQA]�WC���+VKW-���d�)�Oo!s�7%��\[�ɾ��t�t���M~��&a� -@ X}b�v���{���O���ڸ��6$vv���|4�f�1���iN��WԳ( lԖ�J�w�@ҸH��wK�D�&#F�����~sw����;�!�ء)�;�@��k2�s]!��5�v�k�e��Ȟ�9����MG�שG*0����H�;w����r K����zO�4�%��>e{�j�HwB��"��ȳ���z5�6�����o���S)v�y1F|�Y�	%$ҫ�6NUN*��-�\�h�2sctR+�V�Z{UD�D]��Ui�7a��Z���D7���8��j��6��j�hC�m���䳏G�c
����E0��/9Uւ��ʽ�O�S��|^h��1��ɤ�|m����K!��\�bH�=�����n��j:��h����w..����x��F��s�m�w�*7�Pi�ùYq�E��Ü��Z��f�z��fo�Y�#��@=�b�y��]L'0���P_�z�q��Z���,K�8A]L�6�����B��uƖ36��`�gm}�E~���Ʋ���8����ˆ���I�ҷ!ǽ���w�BkY��w�)�5׍&-���iDoU<����wS�K���J��Sk�����o����H�'�6��{H۴��#Ky����#5SGUg�Kށ��.�1�).�3���Vg�����h�P[�*����@1I�S�AMU��!W��$C��w,�����쭷f*�LDg�#���x�9^6~�O5�@jC�^3��w��;��FֆdDϔ�1c�d�C������t��C:�H���˟�Rr�������0k��(��)R��Ό]�����i.6�-J�N�r�3����Ԩ��J�O"l
�?�����e>�I�]�!�k�u�-�!�_������`9�Oy��B��ֽ=4���͔lY�(U�B�mE�k����.����RU����?���bɂ��^�v���������E��q��E@oCm�|$b��2RH�[P�8���$�R#"a�IhM�A��	�g-�-�l��������%��C�HP*��e����x�)&uNJ�U������R��7�=a�A�B֝��Ꭰ�pu�_�U�� ���<,�`�����+����Z���A�i<H����ʉ0�i0ڀ�-���������J4�ȫ#'�����2������%~��m�28+L���q��"Fԗ��G��a[&N�Vx9�ӱ8�?E�#��um�����b�%|�G���5ò�Z��j����U+{��z������(��GP��ú�U�0T(��xaw�wd&�|�)R����#���5Dq�U<��EV%y�C����#ũ�?�G���p~򢟝�~�	�����.��Kl�S�ȕ��q,zN�5BiT�iX0�P_�v���B	�z+���f��#��o�8xK U�<zO�L0̠ܕ�c]x���W�.XDC9R�ǄPH�Io�<"�� �ƑkFWw\R^�-���Ƥ�����p�߃��Qt�d�NJ�����l���\��ȳ��]௛5�����K"����b�����!m�dܦA�����~�p��q��p�p5aԁ
�,�Bi)�X�4盗K��X�i��kլ+����W�~�K�K�l(�Z2�])��Rk���=�^�s���P�?�צ��y��8���D����&�8j���=H��Q�h`o7���+F|���@�ը2�n�.���1�/����NM�b���������hq��i�_��yl�5�
̸C�ݥ�朼p)����FR��dX�%}<r�7�Fe2*�]un5�:8�4�g>ڋ9�w�&,xt����F��[@�e�h5�~�ؔ�68����Ǜ���t*�3+q� ގ=F�+-�"��hO�1|�w��.�<e���;P�Ի�S~!��d�c�P�����+%�dUAT��尓#����{G�q
��/XN0��o��0�c��ѸrY����c��~����Ɇ�mR0'��)�l9GF|�B�5��j��y3@�#��B�>��	B��t�HyKؘ
��V�Il�����}�L�ؘs+�`�Q��QL�㵨�t�Hⶃٶ�˅��������F��B\���=O\����N%���'�O+4J�G��F,m�XBU�y�RH�L����Ƃ̍W������U�/��]T�?�/�,~���Y`�EW�f��]�h~}N�Tz�+<�,_t���Ʒ��	o��cP�S�,����?G怐Z��#>Q�j�:;�p)�$n)����?�;]���p�����8���֧>�rı��`�Ҏ���ৡ/ݾsߚ�a�E�ZXb�ʵ~��Uu	��pDپ�M��;�0_#���I�}���ݢL���kҊX��H�O�
O!Y�"�׊w��-T���mGO}��[�.Dc�yB�9G�[B���G����nWE_o��X~3�i�����[m�ʀ���S�!x�9�i�I��$|3k��K}����!�$jZ�����سL�0ڲC (Dd��XE ��#�@bW^cP���{�F��<�x�+��3��@tP�+���tnp���)7A��P{��М�r�2+�W�3jmǈ�\�l���ş �q�4#���X�.GXA�%	��dW�3����.|�l�xu�+�>�\nI��_ڌ������XS�`��x��$�E�'ٝ�m�����;�o e>1���ɪ��^8b���n��ǝ���3���(l)�^��)s:�7�5Fx"�l�{G��]nͫ �:�
�{�8�������+�o��F!$i��, ��������f�NZ�<�^�i��E>9�����KM���uL��$V:sR�^��wi4���'tq�w�k�����A5����?�IH��l�c|l�1VT�8��dMV��^���ҕ�,���ӟ�>y�Z1�@5	L�ӳ��A8����7N��~�ѻ:��|
��]F�_[W[ek ���CTى�/ܘ�LK�%�Ac �H_;�e�`1]��jny�T��WG�%�
�3�c�I��b�d��{Idi��2�\����h�� �_w@�E�rsno�ui9���JJ�/�Ae"'��X*x�a?�(����:��hH�z�X��e��?��"^����=0� N:�N,ĺ�r%x��>�x���J�~�L�p&�>�+���'�����3��%�%�I���h�OO�L� b��dPS�!�f�'|��&���%�9Ms�G"% 8g�����o���@�n���E"�t����-�-���N Rjы:�_��7��ʞ�_?�D/�}ܦ�s����A�t^�kz��z�AM���] ��ː="�#k�Q�J���-��y��L|U�e�)���VO2)�ש�N*F�#3eo���w��Y�}��@��0Ӭ;����Q�B��I�!)����:��鮨��D����e3ic��h'�����֗a�VR�ru\�&}��q��&�]]Mj0oJ8ܟSX��\����ȡ��f�UT��ѣ-E��uD�d!�?xX-����A�v	=r'!�1׫@E��Y�!�/���	`�Lk�~�*!�|�E�.QY!=u��NZ�wS����V�NM�ќӓ�
樹x)e(�T5��5hJ��o��r�Ksk�S�`�%�a�h�*U[�F�G�h��dC�M�/]?b7;O��Ȝ>������g����+*V8l�u�TC�nӀw*�T�$77`\�>���<Yۢ�'�yj��,��Y�ϡ�շCg�^��F���r���b�1����>��nBY��c��=H`d؏	�n8�� |�_>aeY�N(}qٻA]S4�b"�M�Ϛ]��gA�IK?�F�X}��Ă�:Kj�;#d��Z:���ۗ:���Z��	�����/���;�j����O_'	�w|՟��6j�93Hl�e�w �D4$�exh�İJn7�˼bs���-1��-�9�{�jl���B đ�k�W��*X3AW\�$����d�'��-���'Wh�7����B��j\�E����PQ�%^|	�H�W��WT�!J�j�>�8�w�?=F�iR�ho�[iR�
2�y�k_�,��ݫ]Q�Z
\�/z�ZЁ&������i=@=kP�Y;��+^z�ih�y����Sg�C����m�G�Ƀ83�%�`|�z�A78S�:�(��4�PE�3c�B�"�O�b[�(U�6�v���^+2��|a�I��a��:�}��R2�p���ܓ��4q5���?c�Bg`��!C�	�x����d�\ѸQ��?�OY�v��깖�H-�-�e�^��˰6��RM߻���98�N�(�\�ï+Z�P��Dd���(t,j�W�������"Zr|�+�Y�������4u���i�]9eV�H�����姽M��WQa���j�hTZ]���so��暴�|�� �JTK���)�`YF���?R�9߀��4���?$,A8-p_�Eg~��+���M�`$�u��o{ʄ�h�M����`Fǋ�#�Šk({�����͍T��K�s���ZN~b����_;
�g*���A%/�e=�방��~*�!Z��uu*Z����洱ʍ�iW�/R��q�r5�»�!S$��Y�\��p����@�g��9��h[£KRV��2����M(��Su�w6�'���v�KGB���g�9)��>�v0�K�N��^MТEQ\�tcm��昒�����S��窟����9���}l&O>m�F>��A�1����+�",���-b�.�� Ԋ��.�(ZK0+����1���$��������tj��!a8v�Î�;PFY'�9�Ǧ6K�����x���r�t��TV+c����H`�������ǰ%�'��j���lr0��&�T
0+G��.�E���D	�P~�"� Gǻ�b]���E�v ���yҀ'��j�=	9�q�u��!/Ӓʁ��^�66�)PH�4*:*�ѧ����{~� XK��1�gk3�@k�+���E��	j�#y0�6+u�T��H�~M��=��ѕ��a~�=Qy!�GZ���t��pF����E��i��nD�ؓ�-Um�ŧr`'���6��D!�&}�.목:NI!U�1h1�BY�&��KX��0�P���;\�g�SdG�nL����7u~�m$,b�^���f\�q���<�������C���_y�y��W�
8��a7�'�����ʂ�/�Cx�D��'�\�T�Bw���+��̈�X��;ģ��(c��w���J�S�}Ṕ��͸,�{���PY�yY4ϟ��KK�}�M
�A\r�KZ���9��e_��ȵ�T&�����,�s�T�-K�w2�4�!Jף�#��2!7E��x��8h�Z�*:���6��X=.+�2</U:>����h8�(���^H�X�BѠ�`!�l�,�Ē�	O�ot�*�R�|P}�'�2���-S�䕀���y(O�Y���i�iz�ı�#IA{C��f05���� /�0a�Y�C��K =����^��E��*��w�k�h���ps�q��������P�6�J�O���6�xF+H:N]�8�36X#/�F^A�"���6@Y���� ����j�yBb��P��C.�xfn_��$��e�1A����AIBU��B)?�[zl=d���	+{�.��N��Ws6���W���/q�Qh�����#���N�Q���zQ��Cu����bz�����JC���`L��}y����F]	�@XEϴ΢��ͽȰT��UE��S�VL�d��\�����?���v���;^�z���{T�q�S5cN��/k*Soy�Lޅ�џ�1����j�E�S�v���.|�i��+�DĠ�@���Pt���h������e �����rD�9ŗ����X�%A�,i6ͳ8y�a���n��������c�W�Q�/C�l�K��J���ۏ08�<�c����z����zG��`�V2B��RT�m�[��(����u҇JX�Bk�,�7�8��*@ICە�и1%3�e��!E�3�=��錝#��"�SZH�㉴�2����UǞ�pP�)G�ԕ�/��5����Y0���q��5��ҕͅ��S-������w��O�:{���,��8�����p�8_�iAҮ��w���ڙ�3ƣy��J��Q�Qx�C<+rP��!>�w]�-9��I�V���Eg�C��0ʝg&�E�E�&�⎺톌/�1[p���.&����9�A?�&��~�ie8�6�1ݼĻ���;U�Iv^P���Yd�$�5����&��(X!Ddp��Y��H�p�&�/� �B-���lc�/S�v��F��C�33|N���a��>w�Ṷ|���_�Ћ���Yj���p��Х����7k%��
��Ю��S��dp�j�_�E/����utg�x�N,xF���zuGI�q�eݛ%��,�r��i3=�N�]�,@�DX�{G3CuW�?�	�M\�����-����Dz�"o��O��a���Isr�V7��Js�Gx�	.�f_U�F*�{kQ�f!��}"|<qe5Y��W�Nx��-kVЬ���`7+���<����u%�L՟�Bˬ��e]��~�
cD����d�:�Fi�,u`"�z/	$��k�y�r�������j|�.-Pf~�4|I�8EZ���z���-=�O��X?����3:QJP�5<|�[rу��7U��>;���z9�WD��Ų����JtR�:�F$���痞@O�8Z5��r�OP^f-	$SE��2��t���8���{,�c�N�oS��{��v�*�3;�#,��Ȏw�Ů�X|�mA\f�����9���a��EX 3��)WD0ڗ$o��~�#��p���{�o�����/$���Ttț2�Nډ;�K�K�����6fk���6¢�	|q�2�K��
C�] �է�E"��=�~@�X9�E%��g]0p�}�և�B�C�d��R���S�?[Kq��O��7J�,���S��-tR����M�[�W�L�i3qiwoM�rD=�b?������:Qvbu/|S��bEY��������-�r}T�Q� ���?�/��N�W$[��*�㬗Ѕ-��dG����jTCs�1혷�,9�[��`6�5�~��1d*��PuZhP������X��$,uy������A��Ւ��y�����+���뾙t"~D��NTS��B���M7�7:���ĳöwJ`��}wB� g���*��$��4�r�a��<uϖr2)�����»��c0���X��c��@B���%�ؽ?5_�5q(����_d7�`f"y�L`b��R'��&�׏l�o6k��������79S�AA<M~δ6w�߉����A��s�t���^����B��mu�a�2x[��7il�"�3�����oaV��!�"�)�l���*�xT��d��1�����x��*��5��fwr��u+�k(��Ц|�bmE�{j\w�U8��5��!>k��j~X�nAwV�.�G�23y�=�gV��i�z.>����S�Qw�U��y�'ڱ͍?9o�ۚ��SI��B���H�WNꕨ�"����Y"y��|�߁#"�:2�t��L���/��0D��^ą��5��, 'a�'\����{�����χ�o����תau_�F	6e������z�,�酎��?Ӛ����>���A��Y]�uS�9�Km��!~���U7��M���o{(Ÿ�u�;�]҈{0W�:�d�;�&ڼ���(�<��ar�K�{���o.��\�����b���kG�oG��.�&�P��s��}hw�o#0w^W��.��a{���{� ����U���9�}H�������M&U�8���R~�)��tR�wz��^�8���W�`5y�\��F��9&�7��Q�|bGZ���L��	�'{��z�-�P�����Js�(�tm,B��J�!U�}����bxO�ځG��إ̰�ϵ�6��{�E������e$�ۇ��sm���f�J`�5��!5<�򝠢��A���k":�}3��7D�O4�:�����6�3���k/�A"����0?��eNA�"��IeD9??���_gv$Ac]|��K�r�+��;���V~�F�3�.V[�ZҠ�zR���vŞ�B�p�9>x=�������G"��(��.��a 熬 �!���c>��^A�	��7��\
�a
��F�t�������9�có��q'6�|D���!�5��Rh���<Z|t���a��F�e�j� ��D�$���'������%�%�
u�S�(U��>#��&'~Nяf����2�Tƚ��:m��C
�q�x���g�i��u#������6#��̽�e�������R�~���j��D5+�%r����y��[^߫jD�W~����̺�r�5[�`�զ��U}+d`�I�(��!A mL,�FtMk�c �����gx�=��
_�:�X���׹AM�^�����/��Rď��%�7a�C��X�P���)_�Q!o�x�8cJW:�gi;�o�ek�0�허=e��a��A>X^�Zqk�:����L�Q�,R\�1G�񘔐���)�2ّ�(S=B����6�.��"�9���JlC%�f��{8 ����X�v�)�ܿ����n�:���]�"^/��l~����Kŕ��u�x�<�T�����Y�F�s�@�|?�������%Q�v���Q4~��Yz͙�Gք���Jﶍ��������W���{�����2��7E�~@�ǰ<��3%˘�1��o~#��ld�v�W�qA�Afҳ��!7��_�P�H�]���	�C�厗�o��f���uZ|���|�́p����Hh�����O}���	_�ѩ	��J�����"Y�����"�E����	��(�M�^�U_
� �n��ف�ӈk�j����`��;q�|�z�)#�CMuP���jD��x�� �ǢH�zF�� ��k<�h,��e����o��4yG����vrH��卤��:��7���<k1�{V�*�8�2u�� uH��7��w���ʶgF#���ёgq5�x��7$Z[3-H��K�]:4�FX�^u�s�#�ϖY=�&fN9���*�-H}�eJ�d��Aqa>��
�*�c�����ĞY/?�m�@5��G-�-�{�[�4ŋSH�96K�����?�f
f��P�!(���,8U�t�ǢQ�֟�y�r���;Y�9��R�5{�؎ω5���Eh�ߞ6�1��R���q���}������ �m�x[��{}����{���m�oC�I� �F0�����L������GǛ.��R �s�eYe����W��Y���4��{E�F����(V}4l�� �clRd�5<g��}U߯�\�(߿�įFTӎ{��h1o�"Y�"B���M�̤����+:��4U�|�,:�ߑ�dXh�f�{��A�Z�멒w�N�����ڜm!�̓�\i�j���Q��+�'�g	�6W�D�նz�o��d�*EZ��dc�5w��HX}��\���S�/l�$�{����]�m�����3Z��~(��:����O&a��Yܗu�8�΀��K�3Փ�Z��?h�:*�.�KE�8�n��nM(�ޕ`��4Q:b��9�嵑`�6�*@Q՜g�bFM����9t �Y`i=rf����Z�"�7�?�~h�9/D�9��Ei�:CcW��h0���f0�����ϵZ��m#z��"ƘV��Ҹ셡N�K��Jy9�k�R�0�����������A �m��X���p�ɱ#[�� ��5��ȃ�1̚K:�XK��H��qr��f�72�zP
Y���vS�\�-L���>��2�h`ej���HVΨ8h+�4zƢ?�-'��cA�)`�<�'_���T����	 X���Hp�/�R�R�s0ù@��κ]ώ�h�&/��nK㲻���D��wU��u�����5�d_�XZ�+�ɄZM�GlO
���Pgpo\[1ԯ��<�4[{e�h=�n.�͠���jN��Ig]��l�$����.'��<�$���6�7�}�pk� 8�.G�x����!�D��QQ����j����c�/]� 1-<S���J�^��"M�\�|u�8�i��h�1fXEgX�a���+���q�ɟ3K<��?�����Af^�3��ԥ=�j\~34P���˻�`i��Sw�s�J-��2"�
�@�=E�!��x�.�0-x��T��^ٽ���������8�vx�%.&%Z|�k��D��hE�Pl�\��i�<�J\-F��|���	v9JۄHW�7�b6kN����rA��3 ɉl����T�4���!�2ݖ8C����a���y��i0�I�������m(�y��M�A���kMr*I�s��������|Ɠ��|�y���9ց���p�����PA�2�-�����	�d�J2�����ǒM�df�%w@�2FS�<���%�=TI���`��8Ձ�="�!�E��7j�O}~��07o��ۉ���_���=��<�l�Z)�>���JX��T|;
j��Tr�;n/E��w�~�z��o��;�f�X���\��2�����KW���L�"d���g$%���2|�#T��G�����ln��jW��+���Ƨ=�d���������)�^�$-�;
���4�����2cO+OܝC�m,D��*��B���X� �:�yס�W�FX�wOt�A*}�%ٿ��
X����b���L���q�_�������(�ÂC�%�蔟_'!YqR���@�~Dh����Ov���ke�,�)ThC�R���1>q�9EBI�!ٶk0�I��P���XtdJ�~EI^jp� I���9a��\���]���B]��*/�
y��a�=��{¹�'�d���mp�(�ʺg��My��`�
��,�p���[E�Ƣ�hk�G�U�u��;O�oƖ�>��.�P2�`_IYU|��5�!��}�����,��A=��j�HW�1w�U�lh�=:�c����J���_�x�l����g(\ڹ�T�Us�d����B������6���8��;eJM�H�6��'��J����]B�+�XBb.�\��)w�d�V�+3��D{z���X3��u�=D��h�9@���P�� �}�R�'R�nZP0Y�����Q���6ԋL��{p� �䯬D���ּ;�5{I���hx��`�'cV�qz*F��\9B�!Z��В#��5��@vќ>׉$"�5�=&\c�:"���h��6.��)Z���ݙg�L_-� �6�����B6�Z3������`�ub�'�V����|�%����;�e]%O/���j(,��l�����>�˩%+�zw yr���/5�R��Sr�p�%44�4��W��9���9؆���@�'����EJ�{��(�5Q�{��KN�nJ��eq�L��ݓ��_�����ۣ��)#�iq���eO��#��j�O�\�����pFF|�*�	�gs�^@)I�7��w1�psπ{=-���S	�6�C�/�w��x$�Q������
�n�J������[��D-��.F�z�`7kJ�d�U��8���Yg��:3�b��E�5h�l[Y�e�,�[ޠ���q�Dq_.l�Z��㳳57D��r�䖜�k�yna�\�-/���e�$���x*�I��lC�VO�,�Rbw��@��Kqn��Z9vH��^Ԅ�x�����y1�� ���u*Ć�m����%��@c�fgx�
�LM�˭�S�F�
{5ĶΗ
Al�<����[���|�Ç�,��5��o�G(�'�D��뿶ًg�������V�p�3+���@.���O���#l �D��\y�:c$Ǘ��O����\��������%��$(����í�ϒ#v�g���S@���ˁ7?3�q�  gѸ\1�a$mv#'K��n՘')�~�Kd�亠+�T|�$
a�Sz�V�f][�2�s�$�bi?����
+	�x��$����Y2zA2!Bi�Nܗ�%K@M�#3#o%a)׍c�ђ��\)7[�Bf�����Ҿ����UWϬU^��$l�3�hQMA�M{{�F��%<��䦞cX�cC���K�h[b¶�Vӊ�NVC�<q��~�/���%WX�a �ğ�w�Z�oU��*��O������{���X��Wr��1M�Hc(��� ���L���i}��� �b%+�H�hU�	�pA��`Z
Ր�s�������ɽ0a����U�T��g�HV�Ґ}j@F�}����Ԛ��:[>kDE��E�Fe�`-훓��Y���m�g!��N�.�"�~DX���ԝF6V�;�eǲD�����殶�1w*/hs�#�M��M�� �r~�0-���{N���"j�3{ɮo��³�91��R�����3�3��$������F�BO�0	�Ap�'�`n)w��LU��1V����A�k W[Tc�]_ރm����_����Ͱ�0Pb?�_�@��9Un���Tr��L��	th��{9�g���B������.k˽�	�^�pwSd��,4�F��ˡ=C��y	��N4��͚ӛm��"���
-{���G>�8dA��ܙ�# 17�TY��C�GBh!7M"�'�<й�M�������m���������^�Fa-�7�O"22������US�r�;5�
�R��)�{�P~���m�J����GP����{~����1��q�ܥ#����]�t��7)�j6C
<�����_�v!��>������s	*e%�B�w�wӉP������3� ���S�ܥ��;2v �Ϻ��T��]��U�\�th�W}k�8�ޏf�;���_0d���l��?<����yGXm�UT����:��U�'�?6,���OH�V�U�e����.ʪj���' ^BBG����rS0�.S��}���F����nEN}�ˆ�������%�O�Q��	�s3���p�r�9����� P�✧�ѵ���]�V�W^b�O�f�5�k9HuB��)�(MB��G��d_1��ч^n�4D�l��Sg�Y�{i��RB����(@5{j����P�Jk����xr�bte&O�"�@�gr�g�QK(�������oZ��(����yy��#`��W\�.�l����o�u>��-|?��A�h�M�b�F��p�#�aw��,s�E��uG��L륟���}{Hv,4Aqp��i~iO�	E�V�O���B�Y7ͲD��̷�v�7Ơ�3�<��P�*2��a$i��t�DK��}�ɨ�v�__dl�� �ȥ3ڦ1�t�	"|��y��1��&ᘞ�;T������aT�o�][z�q�y�4�B��4�d8*�ڂ'W,�G�+�"�.8�~���B�8���.L�c�S��j@Gy�f��0�����WU�/�#l	5���Z!��:����ǈ$�N��O��ƶ���&���S)7�ǒε46��h�h}Z��H�!Ov5f�o����7�ǁ�<��h%�amP&���p$��JX���Z~�ui���zf1��7�ϐ���J�(��
��b�qB�T�����9�A�5��� a�&<��s��=�+ޑ�r�(�}e�A���3��@��K I�^+y�F�De���ŝ�6t���:��!P�X�h��q��B�J��#|�e-|��Pv��Nt5=43���2vfl{�l�e�FO���k�A��ە1Dk� ����J�B��C�@<P��`�+J «�r��sq�� ǡw�#�d|�Ɓ�u����[-�j%��_�7�g?��~*���Z [q��߀�~-�J''JH)�9�뤫���[,�C{��!���]���Bv��.w��UK�_����ޞ���Ӭݻ�u�њ��.�q.\�.?gw�J�$/�%;�]˿f,���S�JMh^�\��ϽT~��]L�g{qߧ��Lx+��������I��F��]�j.r�W ��=:�1���nX�3R	:#J�R7Wd�c�a�G�pJ�e�dehpۚ`��&Z�jC�H�/?�+��>S\�ߠ�c���5�)D9~Q���8J��O<�����D��݊����W�2���M�t��ўZS���U���D�\@��b��ج��(����V&�o[2��M��}�c8�B9UO%kL��%_��
\-	}7.��QU�:0v&��1���T�iɸ���� �Z�q_R۝���YE#�|$&��̇���P��Ɗ�<�>{�3�H��`�e����h�PK&�Ҷ1R�~�Q��-��!�h&��6��S��ؿ��#��oj*_UC}��d!V#@��,�`>/�=$X�?aqUf@�1����}�"��~���1{�׌�'��4D~��beG~ie�~�<<^��c�ݑ^N�`�f"v�>G��?�����Y��',Q��������0���f�`������2����i�R:� Y�Eڠ�
 ��ݧ��@+�\���3kߏ˲a�%v0�ƛ���h#Hf�e��4؍��<�Ij�i0;�!�D�:�F�ۑT���r�O[�V��±�:F��К�\u�2�ۦ"Bǭܘ%̩N�QC�yYEۛn^A�k��ԓ^n{ڽ���л��g��+}^d��*��Z ]"�Q��4�W5�h�H�V�Z��$��!Ap�1��{�m���av��Ӡ^��Y�R�8!D��Ur_X�~�k�q�*'���16�!���5�O&��(���Ԧ����nz���F�{$������$��S���J�H��P��*�n����p,�l��e,���u��6f�r	E���sK'S���T>:"��f��n�o�Y�2�����K��%a�d��㉤�J�7��Ժ� \\~(E�Gt�1��u_zG~��xݚ'�JĴ0�3��"�it�rL�o� [�������@p��\��H�+=��Z<�yd���(�(�[�E���+%'�^�M��/nl�^��
�K� �U�UG��]p�退0�	vA]���cLw?`��}!�S�1$zH��WC����\���G9gU�n`�W��^�X G�0.����K`C�n1�i�,�H{
�R�ag�T���yZ�1��V�bSXxt���`/��`�g�a�^m{�� �`����Dwy�{F�Չͧ��S[V昙~��Q�1U�O��A��F��D��ά�m҄m�}?��c�#�d��7�ډ�$�5T�{�&���ca����v��p����^�^��>��?��b;��.G�����#��2������/�G�1���a� �w9!S��T��o���hy�F ����9dJ����1j)�>uC�xf�w�i�j`\��U���L�uyL/9
�վ�4��dͱ�}�˾�\����gy�mc���}O~;]܋=|95/�wE�bFHR���e���ɢ�J�r�Y���-���E
%�߈�����-h�����z��˂z,�,�M�����KrLۏ��QY2�r����;1JYa���3��Ɯ޴(� �y(�2�ZL�:��m%�	�yz'�4��5>���X�6X�䆪��`��Yz2��?�)���ȥ��̔�y6i5�	�A�J�>f�}�[�Q[���y:+����po�