��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�8k�)9�k���J�f ۘEN�R��>�Ug:�&�1H��������yAc����T�ƿ<���7��
�ַy�x������cCA�,؉N/�R�����I���YNv��X�q�>�!���O^�O��j@�c̭�i�k�U�.�/���H<��C����c ֽ�rR��H��0K�k��pȰ8cB[��5x�^{�XA������쌌Vb.
+ҴΞ,c �����)���)�L�.!n_/�etj�����;��y2�%�69ͳ(-�-�����g�碌~�FX�u �z�n�J�:�.�����,,�(�m�������4��Et���9�۠��\������C1�@����p�2��s�xr�4�6��8��~���vܻ��&X�p6��rz��E��/!c��ȅ~+�����Ɗ9|!/�Ĝ�U�������B��������OҴ k��^����77�(���Л��e;6Q�2g���yS����b'6T�2_]�.�u.�N˧�!B�\��q�VX~��*c�G�R8�΢&"_���đçnpOK����1Q�#�l�$'Ih�ߟ�6�`Ȭ�_������m|�n�b�ogg�O4�������h��r7�q�vU�����x!+��9��omK�E0�����%�3��<QΎL�PuȲ]�*�X�����!d�v��З/���;�ly}�#j���|��1�y-�;�t%l��E>���9����?)v����yd��\n4@�7�.�b����T�=��_"�;+�	�U�A�:~_�EI�C�����gN1�F""��<�T���)�؜}����z���'6n#V���U �;�lH��l՝��L�Ã��(IK�!D�{
;��4���qK�	琷�u��
��A�dD�!�{&��e<c�xWn;67��/,B=U��L�c]�O/�V�L��c�R����Qv��ш�ϳ�HsW(ۀE�^+��5�+�A����.]�!��|��,K֦\g!ت|4�$�Mpm�b��(�5{��$'6�E���m��=� B�b�詻d���t�hB���\?�z���f���or|6�ױ 61����Z��cI�@���O�|w�=M?��/)� ��I���9��|����u���_L��A�F�?�B��WݜF�
O��Q��	-����l�d�񕕲Y��6�/����[@f.�CZD��	(�Қ������o�=�\�s�ƻi��-��3ܫ
��C��-�Y�͛*P�U�q����nL����u��&�Iwﭤ�m�]I����'`W��<����Va��4'EV�$�k�L����>J���mF�]�@�
a��eAH������M�P�"��U�i�����8��2Y�&����F�uݰk�O�J���'��L�1s��մڰR*#\��h���e�xW�1����M'��V��3ؕ��Iu�RAw
S�~�J�� �*�tlԖ�>*���Ls�esD���}b�%�(NF��5���;G/>l0���n��~�t/�x�.��^U�����X�����YX��$(њ�  �TJ���rQ">n�%x�m��@�3�ŉ=�R�0\65���u��Ej�LǙ�]�Y�8ߦ�11�<��3AT ��s������M�j��f�C:���������l2f���ƍ͂����N�}���2jP�1!:!��k���l6f*�{��1��+4�ՠn ɞ���r��B1x�ڡ��}@:��]Zq����T��_E9D�e����P�� =k�4�r%B����m�8q�;�-�0����:��Zw�ѯ�����{�!P|=��ymH�%~;�E�6�S2��%��������M���Ω���Fy+nM-$ᬼ�K��ݶ98=B�8��[��Z�9i8�#�j��6r���%�x,��4�Oѣ_1�>��oFC�z���\�$7��hn/$~;��"b|����j�A�5��ׅ�t��:{�^�KI�P)�@�L>�K,��#���W���۸������M�c�hϣ`b�<�.QX8Ĵ�4%��K͕UJ�r_~���w�NH_�BY��xi0J	,��d2s����g�A�1;��f�3�ʶ�$��O��$�t�L�����)��O� 9#:����}�J�t�����H��[�D�wd��t��csC��M�'�cSZ��|������� �h4���bV�P�J
u"w��a�he�
�����A�.�B���6�Kϻ�Uu��]|-��� �@S���8��T����)D�*���>�����E���)�{��zK��Jꭝ��j&C��V_O�g��>�S��h��t3x�L;;U_+d�s�������"���Dx��V��*4ͯ"G�T7���*ָݲ9��-�������d�_��㩀������8�},���'�MBe	����}7�9�Ͼ��芌���8���2w��q����16��=De��bo�}�=Y��&QvZ
E��k!�LA/XE�jo��{��4)���=���/ݮq��mF�4��X�;_L�v��;!�Qի��o%�b��z��.��vn��̨�J�ɓ�Kӷ��X7LG��Ś�%��3��T.:��TRyI��m���zh>���Dwָ��m-�]��7��!�d�m�؛fpD�R�/8J^�@y�x)�(M�Y�tL+z݆�5��
8T֔�8U���~t?�9��\�QN�М��IW�{�ߴ�az��m�s�����Zo"����#���vY�U	�_�1����;��H��g{���
��<��Z=Z�;����z����R(͈:Ȼe���aXH3P�u��]�J���E�0��@�a
�����I6p�����.��PT�ٞٓ$�D�!��t}Iva��@���p1}^>�Pi�uWx/��⵱����`�kqBT(6J�8(���[�(�?蠒�h�J�.O�f_���{D���:�� c�>E�+�_�eK�C�wǄ�Ybd���a��?���2k�[��ެ�Az���~<*?)<�F���w�����jCPa���S�*�\�������B��� ���ϟ�Qήw�4�q��"W}�0b6Q#��#5�*�
B��z# I��bņ6�t�0�� ���p��*c|�{bU�X�_���I��訳�_Ôܕ����t�ܹ�t]z �|j�>��z�����$��L -쀥XX֓���bq 6��ɚ<�b��:W\WM�<^zH,���"��+���x�=�H������w��1ȼ�4F4)?sg��a���[��>#*�x�H�R�h���	�W8���`�֨ܛ��s����>1���̭i�i�,����~9l���h
0�aQ�G�l���|��8�N��Ӝ���*`���n$ڶ+���u柠a����-��b�Ћ��(�h�ltw5��1����	��"�fF��F!B���?��]'�a�r\�����\�8ou�n�;�3GH�����;�l�;8"U� P��F=q��a��:��/����>D9���ĝcނM�g�?#~�&,��j� :�>�=��Z��/�f�E�,���~����� K���k��W'e��Ѣ�y@��#�A�L����:57|�dBa����d#���6��O4qb��;�bDj�	�=��'PW�����jv�:��͉C�:��lX�"�������5��/���Wf��_T���_�h;
vZG>��N�"*�(qa.��1���i��~����� �W�UX�t�D1��#��e���:Z��K5�lo�]1�	Rm����/
�x�r7�Ln�58����5�Av�=׼L{�R|�R��-�o�9�HKj�x�$Bĳ�F&,2���2C�v����2p���<6+��!!xN�k�����z}�r�W��w}��dC]'��Z��F*r��ޒ�6 �q�G�7�D���;���v�r�LT�\�]�����ߜ{�_U�;9F$&;q�&�Z�A5*.�I��qQ��,GWb7܀H������j;��mr��cM�JT��n^P�K�\%��2C#Hli/f�n�Zxg�a���lK�9)Qd�eHK>�S5m��`w�����N`�N�����&��sA9ě�Z链e��hI5�:�����N#VD�&Ay���×M�&�r�|e�x�3]?p������l���a�;!w��s7�u<�<��RJJ!TR�`��K󒜃�ΰe���S�9�7��F��!��'l"��\�"�Jlo�MF/��Si_=wS��ϭv�~�܃�S�2j�����>ߺ�2�������ʀP�1A%W�׃����6�㞏D�,�Pt`�)2yq�*��E�wP[K'e�h]|j�rC���_Kߒ�m�u�0�����.{E�؅��y���%��o�@�8	Fa��J4��.x�ZKkD���D��6�I���Ɏ7�j�p���Ţ��؃F*������c,�d簤+��biU�u!��v崃?��z�bi1o4>��2r�ʭ^��=T�H�Ꭿ���8�843y}��A���->��� �L�<��on�YCUV��d.(��0�QBe_>rL�wM��� �� _�Z�?x�Z��:&�����[T"ʅp`ce��[Zj8�0�Bzs��AnS�H�R���q��J,3.��z�������IjXDoG.�nW���k}�y�z�!�O�N�z#Sl�
��1��7l����bII �"�&7#��^E{�|��˚d��eq�f�"�T�|��3,��݆�5B�n,�R��oQ�]3`����bykzg����<e�%�%��1�Y���_���]��(��rJ��Q�7&q/�|��娑#�egvF=P�ۛ�E叽�V���ޯ�}�	dP֢��i�X&[��a;�o���t.���ܩ�g�V��2�C\}/��2��n�n�60��Ԫ���MQ�)u��]�H�t�*u[4n�K)ǅ�����R��qd����/� ��z��9�)x�����)!=#�~�Ro���/o��s���g}5�w��WI=�l��"���<ީ���C��D%(}�W����7\����E��S�U6���%)�V�՚��oy(N[i��V�$�<(=�*�5
%a��'�7��"'{I�P�3�9� ?�Hg,�*ƛ��-.�� A�#��(�'&�g���A�B�����ϝ��ῐ+/n)塊'�Р(�6�V��-�K�˃006��Rj��V5�l\��r[�}F����tk��!k�a�C��jj��+�n_��L�a~Iz�������J�eV-M�b8?�sd�,kvgol���n�p�mquټ
�	v��ᱯTydſ��{��y��eߑTH�{���{d��"��p�2��xK�s��Q#�㌙mH�YB.��~��u�^���B��2�wks��>�;���=ؼD���㡸�3$�A�^J�.EK�m�U�A��t5-8��=�墧�n.�eݣ�_�p,U�IE^��o�ָ��0�5�뤴É�=r�'V�z۶����4���(���2!�{�ig�b��x���ǘ _kÂ��`��F�ͼ�C�\�Z�� �m�������1g��
ɲ��Kh]��&7�W3�I�~ԧ�6?��R?����I�#��C��0�
a�(���R�MA`u=D#я��q&�2]�����/��li�W����y�C�p��1�)P,6��7�1T�Jr�o&�@�_�����
�=<�LZ�o�@sԔ�ǡ~e�*�Ϯ;s)��D�ږ�+u&�ۑa �
:＆W J<�&1<�Z���U�Jee3v�f���eBo�)��w2I�+	�ٝ���v��L�eH�
��B$��8��ig�ącJ�eɆE ă�[4ϑ2��S��`�{�y+�A��6�Qd6T,S۬��pR��QƆ�/���Ȇj�"g���H�mx
��t�gæ��7�xя�ԧ6�LNB��*��7��ib�,����c��1F%@��=�TӉv�s�xri$�CVh��e}�{���_������IsD��~Z=ŷ�������������bד?�F�x�j�0�%�B�▵��M�����/�A��Wi`���&%�4lx;�v*�2�Ҳ��HC	ؤ����q�����