��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<�d�k��R�u����[V�J��C�X�t��W�'��nL��&ޤ�q��xr�nY�8V-�p}����)�ƚ��0�gL(E5���饋�:DZ���!
�J��IE�$b�A��}ĨR]chp��]Ar��,�$��	� (��/�&�ȽxzN$ΤP����2D6~3��*	���jӔ�1��l{jj,��[��UG�	�7/d��y}.�u��`W���յ}�	�ʍ�`l� �4��L��2����d�q+^�� �'g%HؑJ�p��7R�wa�b��xq�Г�^xqV�[���p@Iic��@V�p�����$�~ﳻ�L�����;R|2#��4/���p���)��Ɉ�؟�mۢ��6�F=o�/��	�k��P� �C�N�z��+����M^ؠ��u�1��I,X��hb,��'�}�aZ~�<�m9.㶬,�"�@�rYb'0�<m�5�����u�Y���P��)b�^��ڲB��a���=�bЊ�5��ip �(�X�*�ȗY����ǆ�Ѳ@�'v��0�(�x�[�P����:ɭ���fNrx�|H�˪B�w�a�`T�f����������Bj�ZЖHt�m��e��fO��<���E0,����k%�a�#�e��^��}����9��̽�0<�wr�y���Z����5�>[�aA���#�����a�{.�O�N4a̜�a����İ��=!Ǿ`�-���ny��ķh�~v�5	RK�k�ԕ�@�&5�w��i�x�i�?��ޝ���5VU���a�*sQY6�ܿf9V�9���������pjР%��	�� ��>�%����'�?�6��1�#%����W������?�%x��qSu4��@#|ю�I;���^�8Y���H>,8�q���6m��QU�w�����H�7�B�L�*(�V��s���X�/1Zz��?��Fw&@���S��s��� 6W$��`�� #o¨��08c��G^��G�U��|���ڣ�}e�k�sk/��N����m\J7�k�9	�%Z�x��75��������W�
��5�:1`��\���LlG�{�g�_�
�0�*�����㠡�A�Bg�3�*��e�9V�{���F*_��E��|mRO��7S��`��:y�W�"n���y�է�rF�������yi2�LG�;����H"~ScC�,l��c�O��aޜC��ݮ?��-����һ����]#��T�o\��>���O�q'�7��=T�L!�V�����.�s��,�%��CXn][�.�v�4�B�`M�2�zT�� ���Y�^NN��qwo��F��P�����y�	}\����e*6;�\>��dNZ�!~$i���?n�'�ғ/q��Fɡ�)d�糛��~��P�����6�n/>=e�����T���q&�Q~0�[k���#�N�͐j+�hV�����N��[�)"�E��T��-1��ʁ�jM�]{�24�a �M�#�C0)Cv4�]s�f&�k��v6]��̃Ux>8]*jKk�}����^��h�R�a�_��;�����hi7��u��-���~���x�����u^��2Iv�ֆ��<��x<�j�Z:XHz@��߃\%��2�B(F#R|r���S� k/�1���OL$s�*���ϩOF� 4����WXI�{
��z#���� ��MH.t�;(�2�=4�ڢr>�čI@u�������cC��E�A���T<=�h����E����Z�՗�w-[<�.�si�����-��`���&9�5����7����[�c�今ug��C�c�ntX�.��e#r�����A�[��� ݦ�B��aT��-S�r��u�ּ.'<������_,�}��T)�*A?,��L/ft*|���:!� ���d�a��	ɿ�y�����Wt�E�Ш� W�� ���p3�
ngRqvFie�k8�jg0�[���'<�Ws�_�|�����p��By���圣)r|s�f�����D^�"$�{#�֚L��ˊ2�����������^�?Jp�p唛�f5d��`���yB�.�T��X]�$����C�b�A�2ت�h�g�����C8����;���ا6dF�`lg:ɓę˯��]u���gbf=S��k1� ��7���2 ��!�ĂY���A��g?N�pU�ȩW*�����W'7����J���өXrg��F��&�h+���k="M��t�O$�^So����>>�Ȳ7js�!��g�ǲ;��[օF?�)����a��F]*=*��X�ӎ}�q�";���վ�x�v�\%�ˉ��[@N�^�TtˮD��!u�6V�"�$x�jY�iɅ:�j����`�{h�^< pj�ޫ���D��A|�=ǣ�*h���7@c�,6�gA�`�O�.=�G�G�����6��1��J�`���6�������w�G�w`��'��x�2��j�5C���a���������Y�J���1@W��t�uQ�]D��ɐ�u'�u�@�[�[iʢ�x�˻�G�Se�r�9�D+�&TR7����1��/k��[�c�O|4L�\2xT�%W���O�����6l1�~M%�v�YU��Yw��;D��<EqG�~%4��4����|�d�/�(�W�ZҷS(�E���I>4��ޒ���3���V̍{j�6�	V�8z�{��!���GF/��$���Ov�T��7Óz�����v�8��8I�@�L�ԯ+0p?P�j���y����#������T���	и��W�E��
'�l&���i��>����C�5�&:��!:[�%��]�=�4��p��,���햟�m`�8R�GDq?���`��x	�٧���\M?{XU�;t'w ��Hw��.� ��o���6�
��'���p��f��5]r��Z���8ǔ���{ș�=0*����q8��aOY�/81��q�Л�d��!H�u�ƻ@n*U��"�Xj�.l�ia��yga�k�M�o#��0�n����_k��B5�=\:�8 T!�ހ�Y�c�\P� a��ytR��?�<3o*{zh�A3��Hh��Q�G��%��!��Sh�Y
�[F� ��F�p;����f8���3ã��v�Qt�dEy.��Q���F��WF�
r�e	��G��w�S�����蟇�r.�EQo�N�fzE�m)
���Fbv���F��4!��A�oQ#�JdjT�@��POy;�!N+�н{DH�oĕ&��L���Gm~E������Su���1b��Ta��G�~�W;i/��W�'�N�<%��+���Y��nSDd�3�+nuwp�<q����Z��[��\���	� �~��V���[�>�ϥbpᘦ���64hg	�^�0$����r��&�+�q�ȴ�0���S������Vn�Ew�������"x��F>[1 �5G��-�ԨJK\��)��X�ø�-ZL�qZN!\S �أ��lQ|)�W��,������,?Z����6�U1#x�`�i̪�H�|�=��mG�l�S�a-�9����/������,](fx|�ī&n��9IZ?�b�P���j5@��Q�4Ԏ<hm��)H�!$B�'q=6�{�b�3SF�ml��g5�D��
���(����Ϯ��A���ѐV[4eU�ݷ�p_����g�{�Ҝ Z�Ag�������n-��P8��"����F��@P�.Q�e�ځ_���Y<d�៍��/o����
��D=60u	oP�������=6Pg�o)�����E1rRjg�52p�9S��5Sa��p�
�_K�,�	h��x�J���x��y�� �J����O� 3��@q�<5*�.�]����3pW)�O��T4 M[DvZ�C>�7������}�&����CF����A��&��l��w�uD1�_b^HV({�]М��w7p�iQ����R[ՀR�R<�����q\Z6��������<�-�E4���㭒uBͽ�M���C凷�Eb̫@�WɸL�|~�4�܁E�M+z6�U��t�)K+W��C5�V�w8cҰu�b[��hTk3֐�Y���U��;u��һ���6�QqL�X����M����������L[�kp��{#�����Il*��j��2���hU����'L��w�������ƴ�-���nh�Uo�1dCm.#&Nȥ�/��0���<����js�Tͅ�F��pH�h35�^���s����C��ڬ��Xk�����ɬ/��
�#\]őt`�,:��yd�7/ˈ<�g�F���>�V�cȑ�%�:�u�3W��Zm�A�yKv�F�3��,ŏ����uҷ��,�k�Y��;�$�T�F��� ����x�o��vG=�([� 6�GJi�F�'�Yl��u��*9���`�`��2�'O��6?vn��\8�I��t碭%�ɯO
��F��,�<�}�듌���!ǩ���

���%�-Y����[0�-i|�uLF9)��d�5m���ىi-�x�(L�����/]�]�������AC$Y���S��/�+yp[C�֋� ";(�rk��"���K��^�Fs�'
w�;;�PY��0���42B�b�Wp���[��p�V��.J�Fa��0n�N��?\����&��6*�����؆��뤌�g��
�M�UW��cc�����@�@����[��˪���'���o�6<F)�W��N.E�!0e{m����:m0�m�o�qVR�4�=M�h��ʨ��7��J˩bh���嗄z �����@���OU.,3��}�*BD{���R{��JN��a���w�q����9�%z,�X�Ac�?�Lh���.]���S���6��T�F��J^d�N�s�q
�O���ᆑ��@q��):��&Ǥ�5z��9�r�(��Cϲ+q� D��Tк����N5c���&�#yBD�Vr��}�,����1��,םR(Bt�%aK%��]�A�JU�>�X�}A�':=���?��Ztbr���v_�!���Q�󅣰�%��V�4�DM��R������d��<�SJ���\��i���g) |��4�x��ķV�d��;�wVF7���{N�0K��6e�W)��\����):�"��s��9[�Q���h3w�ц�THNn3T�\>��Y���%�P�n�3�<>��RSfgh���U��Jی�G?G!,�tg��Z��ahŉ48|^�����nF���(����O�[�	���\�4)��i2��晊�~P���@k;��A�nSOB�����X����#�!�b����8G.���h�a��Mh���0Ņ��f k�O �����{��4qW"#�����z�c��}`GHl����䊷?�73��b{�.z��H�r}7=��MXm d��f�b��˞�۪@Ƚ5�<���U~#�z2 .��x ��u�Q���&��Z��~��iN~�tq�;��a%�CK6;�� Yco;.R3��*���'��+*��vL�8h�K��CgH��8�`�4�@cv��nh?nΐl�8��bY�㹙j��2�y���X��o��eD�xk�z�6I��� Z����\z��Pn}�u��n!�A�� CW�J�H�Evn�ۉᴞ�wf����q��c�u&�Ň}<��<flc�����TO���������9D�*�b)�F1/|�F�ʢ������!C���F�jy[���C$�}�xs�-Ӈ��f�aH�)��y�Q�a�|��=U�^��R:$��/��LH��8�߽Gug�Mv'�N apyIW�I�A���R�u��[,:�iڴ��1����D��Zt@��6���^#iR_Pz	��-�?���?���ڏpL�&�ῑ�t� ���4���#{�=e�/���`(�����*��/5��W���