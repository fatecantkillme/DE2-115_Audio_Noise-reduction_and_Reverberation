��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|ۧ[���v=k��J.�b�ԓ���y���Y �g栦O^e��8�����W��}C�͞u�!ēB���sy�,��7�ޡ�nѽ3��.��HI
�8���b
�S ^��y���"E����ڜ��g��V��)Q���T��W�*���*��c�5!�B�ЋC����
/.ZN[6߳�oSV�Yt�ۉ�|+w����f��3���#&�O�pN���s]rtw��ҾF��R��"Tq�nP5F-A�{�y�a���\�d����b�5;�Q|9V~�&��{�V �f"Q�7{��z�u�J��"tH�!}�,X*���+�욠fB�+aA[߶9�>15���@������ǡ0 �G�*N� %�M�k��@�
����i�D%�yX�š���xo��<#oe�2�̼����4��5��!3��\�R9��ʳ��G�f��7zۆ�]9����/�<W�����|>x@��&BG-^��-�i����y��|+��9o���i��b��'6�Z�t�Ԏ�^`�$��IM�
t�<���ň��u�/H��8�%`3yp�҈�o�&�1��`�c ttw����Jյ:܁���:(^�*��o)uJe4�9ؚ-��9�`�G[z���H���!h+i8R&��P�\�,i���պ?���9xMk��))�9��f�;�
��rX�]?�_Ƴ��N�SG-�N���b�D�����p�B�ťgo82'Iɽϛ]j�� �u�l�:a�P����w,�/�@2����I.�����IV��N? �YN�*�ʀ�Y(�\50�Cҥ���k
~^q��$�O(�2�UG�Q�M�ϳh��BB��
$n~V5�d��9I ��pV�}�f.x�)W��ZO�\���-0�����?!�mu���ەMB�lβ�ǰ��bK~hN���zn�\���Z��<O��ٿZ�����������$��}�M>�#~��Vb���ѫN8��c�����|J�c*�"N�.�K�jVg���d:	G�����S�{���H%]b��[R�l�@��'|�>�U�$�[B�ҏ@�TV�x�O��d9�יC���[�x��]-�i�M�������noZ�|Hq�
�
5��L��BMMI�l�U޲�ԓ�粑�gMg���G\��-;�zTwk��pDc��"��M�p�GoV�R�f0�ܨ��O��G-��hW����`߮��G
Q�	w�9g���}��D�x�O���蒹ܐDL�{���`�NR!eC�)�D��Eua-�jH��e�sҖ�u� �ZY�F�oL%�N[o����_����p�ҹ}*�J��&���
ї�f0���,��c� �JҖ�gTc�ѺՑ�!\TlAE%V��1^C�!-s�4��@��}rb4Ў@����gbSX� �F��l��.��a�9�O�n�]��{-8	���س
m��ꐭ��[�5?�j�i@=\�̫s�4�qK|�%(o�'NƋ:�x�.u�ޔ;��i � ��Tu�Īx>-���x�(�̿�~�(�L L y��2d�"f����H/偽�.{��yɵg<�+��ސ�߈��$l��T���#���ع9뺰����z{
�`Mo=��	'	R�;���c��H���E��	g;�C@�ہՈr&�p���.�n������%�g�������+�����1>�Z� �U�n�(m�R"l��=�-x���y9���b:���r w�ؠ?�13댤��kҤu� Q��ֲrg�Z���p��S�J'�r�0�f��m��T��$�8ʺT�O=a�V���TK#�i�z�	��90X�x����h�8s%耚�@0��Q�D5�1d�
1�5 z��ڶ�y�Ʉ��I��M�|�뭄�YW.��EUڔ܄��p�DW3�uf*TI�F�����������/����V���_����2%�[o&ґ[���BB�l5,E!�-���/nˇ��g�b]���=�wqa��Y�^��� G��.�kk�-<�	�<&����x�c�2.���M����0��Z��I�Gr!�$_O`eGL���(T3ӹEW��2�K�OX��!2>�/p��t�O]��~�X����O������l�� �r�TCg�^�N��vڕ���Zv����\n<�K%�9���ˉ�n�ś{uog�L���I���M������!�cK�������Б��[C�w�-	T.�������?1��ѩ�]����WC����+L�x <��zD�.֚�p�;�g�E�R�0*B8������N�-��K_z�尓*��,"`,u����+Z�Ҵ�POLU�i��b��-�a��L �D
�t��Q��_�m�8���9���gk�$ב���~C�^I��ɋ�#��P��!{��X��x	(�Ի:ؠ���2�qL��k�����ѝ�c`AA�H�E����%|un[T��L�:��o���e�&�;��Cv�^��,��e�i�vo���8�B�9�0�yE{�����s��7�����\L=!������.���,��y~���5.�߻8�������J<F? ·��"�m��L� `��3��T�@����7�� )`8L�q��.���Ɖ2����yA�d�c��K )CF���f׃E.���p�1�\���]$ljiF�}w�0�Q�#��v�> s�*��gs�j�:b�	��@*��Z��u	�@��cy�	�0S��'����y���%��p>������4���LP9�	!gJ��n�u�y�vl�k�V��f���������*T���^�0��H��2�j�ǧ���omv�O:;��](Ol�R1�w�j��i��"�b��L�B�M��G��0J�A�J��[�m�e���	]jV�"Cy��zN�pNT�w�"U�{�������zx� �Eox��Wm������"�,o��Xw�k�8��ej��3F����Y���Aī���TԚ5,(�/�e�� �OT����mL7����B���E��\�
~�N�G'�(��k�V	��2�k$�U�g�x�_�8���~ 
gU�)T���l�?�o����5�C����#Y�ey!�G/����D(zK�ͬ��Hx���f�qC.�JD�;�$f�)2�[؊м����;��7�7�?3��I�i���=C��*����
����c�UhpLJmc=f�S�.'�I.��|�c�2���o�=^6o\j?b���0��	�N>}!̸�0��m�Q�u��u���*ȵ�8?o�o|����Z�]�Q����m���Nz���_x��ECTs��淄;�� _��qͲ�y�|=xj���0(�)�U�������AD&�[��;�h<��n�ȉ�X��(y������K^�ky��Ex@]�u|a<�XX�������g���WYU���߻O�D�k��SM�wx���V���/���=M����P�|I��Z����� �=m5MW��Șͼ��,�Sd�I��<&k��$|�W]Ӱc���m����o�7����4�j��v��)�yϷ:���o�+1�i'�ܘ��������#�u��e��R�?kY�-���]�T�xL� <]Y��Ħ�Z{}�Ů7Z�Z��YQ<J�a.'2y���jJ&Z#�%~2�p@ek���n�H��#�l�Se��f, ��`�1S%y��NE!�(��-�k����%G�ʔ������C`0Z]�����[���P|D����`�0*q5.S�Fe`��8m��7�����Ơ	����K^i{|fcq;���.���w�7�?�B��I�13˵*!z��S9��<�R����̹J�u�)� ���Ȩe�.�+�}�mU,J��"�U��Ьa�X:nW���N���,�i��k�Ea�D�{����D�K��#��"C�Q�xA���qҡ�cYx'���5� bQ������]�b�����֘�>p}̔ј`��[<�yb�tG�H�?/���	6~��~����b�����sJ5ܻ�p�Wt���}h�˦�~� �B󬕌��@��'�"�����3�<�!���]`����@�j%l�B�zЂ��<a�Ө�X+eR3���O���F���%�II�J%��F�r7]������bv�	��!?��Q��9��*�m#��z��zQ��m|��FHՖMZ�6��K��FĪ�\+F���c�G���}=[d�-9��n�nR����"D1���kΔ�Sw̷���6������Yz����N�V��` 8�|��q��;�/�t/"��0Z����&��B���<�>�ɴ�ε���8�*������@!'�jk�Q��@��
[8q�lk���P]���p"K� �- e�g\�*�&��X;A�w���AT�?df����=h������(z!���Ԧ����*��Ş�?@�A�7O����Z&Q�{	���w����v���j��O��sN�~^~Z��j����D��� �z���-Ù�I�26p�t�>Ft��a�g�+rx�!��ԉ6�eg3�!�Dހz��Y�^�K�"Fy��@� ����8�"���r_%~/�{
�t�U�I]�L�n���C$��p�2���F�GY���2��n�����L����#��C��%�g�����bGFd��zȲ�bs�����SU�����i#@��e8�3
���`�KC��Ҙ̘�y~��i����|�O�[d_]����ۡ�t�9sf#M�8]�h^��O�.��&5iD�F&*���}3����4Φ4���3yH����u�vG*�5��
�T�}���g�G� �����v|'�GK�A5�?��:cf�{[��H�%W]ʳ>��� �4˂�U��#\cG�q��
-3�Ź��H��EL�s�o�1�`Qnj���:���O��H�+%
�c��C�{yp-*R����� �r��$6O���ǘ˥�J�%��9�/�m����'
2vTh�����	�#G�x��2=r�RK��`�	�ڒ��I�9��T(��3H�N�C�	��:���/�*i
$��=���ZH^	�V�ûƣPJ��9��C�;Tn���2�^���#�!{�k�<D��K@��Re����{�N�-��d{�.��Iqi$B�Ķ[��&�+&��>ϟ��)���BL�4�q�z��Wswԗ��\PY���`���B����-;��J�{�甴^�?��V�"�[b��������[,���j�i��_$r�/�̝�/V����� hF/� G^_H�/g0�\����}��� 5�yMY�@�j9� �U�tZ���{�|�.n&��v�4�M����I�Y�
M) 9Qu=�o�z�θ�/��"h�r�.��G���0��ry��Iz�T�e����%�*�����-�MjhE/�h�$��B���搜j����9�\��+.#x��4�4(|S�NƦ��������ӎ��}TV��%�	�m�up�ߙS�U�:Y,;e��<�/W����psv26E�N�$�C5�7_х��5*��E���nW�d'Z�*��!�W�G=�H��Aò�	;����(�;�����&��X���!��8���H6.�=�큤P��Q[(~���	����qWz�[�
���p�Xn�M�o���F*6kFd+��PL'�k`o��;[��Б_��[��cޢ�eR�C�w�A�1m�I �h#�8����P�0�6����[�y�����Xv7���7�� ��'�ĸ��-N�:C)�}<��#���A/a��Q�7�2��V�������{ܧq5�¡��kC��4�@��MDE�^��#�19���\�����0��bw���VV�f=��4����㼾�O�.�r>��t(Ն����<�2'�k6�YȽ�NVq��gR�@-�?R�n�X��F��'��&L	����*�8�6W�0\O��aO��"��4��N����Z���u�0EaF��\��W�J����p8�T~S��p��� �O�V`��+�~w������9�S�ѓv&�W\��TX���5�<\�L�+wd�ќh��ڸ��~�%L���A� ��1Ҙ���N0[���g��0=?��va`���"���p���ik�������+����9[Y4U)/�%���f]�|�f�t;�X�4�
�>��}개���nY"�<ڸ!��됕��l<@,~H�4*o�^��Ry�����*�Q�Y���g��]�׎C�VN��P��[mhq.��q������k�t�%F��U�G p{�NT<υ5V"f\�Q�$�m����*C� =����?��tY��}��ޏ���,�����dI|;ޔ�İC�]�h���RA'.���u��t2�c"�R�"Ep�f��/=���/�G�l"l=�S��r����?��<��Pd�5]n6�)��U$�Tv���7��Փ�\0]iN�vX�v�]�.��_��âO_�8g�����*�j�e>#��K�*|���<��y0Fʶ��V�o���Z��Y��=4�>�u��� �^���,��a�s,����[NI(����{���7a����U"K�L�~�y�A.��]ފ�n�2�S�KJ��e���E�%�S���_��o�"�[A[����عގѺ�#}����#r
=��,���rAkth3��{�	!�t��ñ�q�Z�F˿6��Y���?��c�^%}� ̠7��**�8h6��^V�eHJPc�/����o%���`��"�]˴��^5�Qh���,l���4sOx����v���ź
^*r����!	`F�l}}��9f�Kx�k�E��B�K~���|:���il��{yOC�nq�f�67̴gX�"?�Ğ�1��0إͲnVE:W�;�.���Պ� J)��̒��o51��T;��h���5Ash�_��AX O�(^����
�_��C�\�	9Hֹ�~���@�����ww2���o:�m�5D�2W��߰��:�B�z%�r�}vJ��\����O1�����7���y�A=J�ב0���xɐa�tѴ~w�r��f��R���{t���J�h�?T�$<5G��3>�q�0���'m ��p�6��[9u��3b��s{B� ��~<@�ʀǃ��W9o�+[�<�Ε��"�􎥕ay�¹�=)&���/��"/E��ب+y�aB$�8�ba�O�C4��>���b�gAQB��A�%(�0��F*��k��A��ll؞3��T����q?�w���)�±׿[?"6z8eK}��
����d����
-��ACD�u�6>��yJ�L�t�S����)��������uU�	�dm��,��P���/���GO���O�+��cA�R����싾�X�KJ�p�6�6��*��N�"�g+��B�h�LZ�{�+�j�	�{�:��j�}���a\ ���I�5�ҳDʱYTz������&��>9�6W���	�2����O�r[��8v�9 _J,٩"��Bə��_����T��9n����m��%3g�Ar��t�ͭ��.��v�;��sB��#��4ۆd�DUw�h�)M�=�-�-�L4�@}1 ������Zp碔Xţ����1(u��8��>lc�^ӼT��I?8i���$�Z�M�=/	��t�i��o̵"ڛ�#�IO]=υ�A'���8�Y�Q�Q��q3���LY��u1���(T8��,T̉��8�_�쩅}�?g�h��1wE�ZE��!%��%wb���M���?F3xN;s)9{2	����}����E@�<�҉^0iD�9t��a������p?�-B�����y0c�jV��j�)��E~(c߆�!��Bq@ W�i4}vE�\���j\kxN~�p�S[���9�YC�`b��֦�@�	E�B�!4^\J+E�������1�l$ؔ%�ZH.���C�Nh4>�d\�&��z9��XW� y[+T�H=BS�5T�$��\"��8�o�<�����fϙ����G��$0�������R��+\7*Ԫ<��D�ҥ�����d�o�4�����nᳺ~��I �5�Bt����Lv2Á�s^`ur5�z�8���{��yp��8@�D��7l�fK���{{�)C�ů�D��+��`S!)+��w�L{���}@�C��-�.܃L���#�C�4g�Đ5\��d��5N����T�\��AX��|ی�"�#q7[���.�ה����<C��:{�&�z�%쨪J����S'��uD©R]|���$�M��-0�&�`�D'st��V̃�̯��i���u%q��O���E�@�f#�>��S�U�(��K���2_?Hc:�^���B������M��lng0n�I9\|����^#��<�b$�Q͈ �"f ������)�����=�	��d�JEu5|�д�g��=��h��L&m>ϋW��X?�vAAխDC���}��0�6D�lѠ�͈Q��6)�cS���EZhØx
X��UC(�[��+[�D_7u��=�;o �8�P#5�i���P����-,�L1�d��d�A!|r��7����Ϝ�qڒxCo��anoza��KB��~��dk��SR�c�i��R9;}� )�-�񎬰i�*��!�J�ɳS#OG���u��ldXʟ=_�q0y�-_�k1:U�{ܝ�zjGx����e�G{��ߞ�#D�n�GU+��=�Ǧ�|ʋ�L��[fY�� �ĵ][�V��3��3��߂���»��/%7��Zչ���L��\�o��H�qN:��_=;��]���E�)��l��鲽��
8��Ѹ1�(�"�<S
�bC�ހIvk�Y��x��,�m��<S���z ��m0T�?%�����.���X����"	���(�Я����^!����݇����yH�H�ް�z$K?Q�m�x�+�Yd��R���x,���q����J�Y.OtGc�E���v���[����H @���E��i����R�3{��/�Ӯ�wk��6b�������D'e�����Y�ǿ`~��e-�9iUuv[��ZlvF��<Hs���)�s��{�'�'�"�E����?��F�x-�T��m��Ve1�,X��!w�$tma��3��`Z�����(Õc��&��"�Y�i]mF���=k�(�ۮ)1��Is��Ri�Cy������:�����u���5�g9N�q�4�E��u_6V�x
�x�R��1D$�i� �V&�U��Lr��m�t)�p�����F���ƀ���2���e�.'K��Sk��lR�:�й�ѵ��.�]E|PlܸDk���l����Be�-�`*��(�!Dq�%%j��
7�q��]���Rw�i�F�b+���z/�╝��C?/~ۋ(���[��M+�����x���2��^�E9!��ϡrcB�l�A��y,�wN^Ia��W;t�.�{�\������k����]��\�s�sV�)�:�y����F�Hzg�[aQ�|�������o���a6�~��OgQ���5�N�򣖄��Wt��K��M�]�������2�^#��X�=����M,|�>x'5d�[�����\���P���m�,#83��4��Q����=1)5��R���+���U�-��% �\�s(�X�r�pm�%��f�e�F���J�����Arg�9��iZ�	@!��Y��a�:���O懙o/[�"��l�d�D\�]��7���k��2b�a	�Z���b�����6�n�"���3b�Ҷ��������H�G�����C�W�)���\�4_p��M i.>z��SE��کQ��M��5����Nʸ��%��F�Z���#PݑՉ!8pF ����C��C�y�ыs�?�S�s,l�������{ �#����5�����"� �-﬐p��c�i$/�˷b�+�d1���)�D=����1ĝ��r8O�NI�sjN��~T�3n�!\OF�2Ã� ��Sb�r+g[~w6v"p)AQ0����5�c.�WȹR;^����?�0'�Ɇe�f�`8I���Z�d��&��7i���e��������J��S �[8���J����G/N�O�|o��))��3^� ��b+�:�|��^�;{�r����rpP�7.7���7h��';��~���H!�=Aq�'2�1�u9�h�SU"ݔ�����>Bm3�ǔO�)I���Cn���O�*X\LҐ�b#8���d.%��w�^��"6�q翷E�-'�]��-�s�/^��� Տ,�`޼��T#u�Q��S�b�Zv���ݘ3<e�v��������N��'���iel��C�:l�_��*(��S>]0�S�,�Ǵ
��0T�P�Y.^f�BӞ��5��7�E��Y�C����Dӻ$.�,�}��:W� K��r7~�	���1)�6>1������}8�����y���W~2������ԋknq��`�8O� �pz&��g�2�B>[M�8���| {3k�Q��PDfn�� !k�a�O�$`H��q�e����0���m���iE����#%G���+݅8H_� �%������N�5q�*Y��i*����1�P�i�KD�͉B�<ԓ�'93��v���W��Բ ���ZޤS&;���Bh�ES��δ'M��2�Ź��D撨 n	��C����~4�o���'&�p��C���PJ���Xճ�L��f��X�d��4�Wu[�uAA[>�́������[�����f��3��iv(/�j2��ÍV'0?�i��IwT�@`��9kiFX8γ-�K� F6a(�*�e� ���"�����~5,IL�N��5Iy˳���F3��9Y�3z�G�r>$8�k(ў_���i��]$�ǻ��t�Ḱ�D>��al0��Wr���gY�uar��������F��mt�&#��p�!��\����Ã�c�4(���P�8o�;��WʇO��VG
<cFZ�ej��t�I6��^⅟�[�����F�/��1�~t)������]���E�/m�ܮ�~U���z>�-D��/��m��^A����eU����[�B_�X�7����Ԑ'@�W�8 {���v\J��͉��ӣ�9�p�k}��S�0E�b�7�/�Y�ʏ�<���<�u�[7�?��^@�m�?��A����FZ��~�����UA/�ݑ/ݫ͚�ޏ�ᳶܴc~���s~ߖL�UJ���',���ΉC�v�6t���T>�9��CV��NO�=������0����KB#���r�m�gM�x�ˏ�y�ѳC�f�	���Z@�bn"Zc۸$UY?�>Y�V���b��cA��'�����
�X^�{u0+�?-ҿei�#�gx�1��
B3{���q$��{S?D�=�/� )��+�����z��tUɧ�x�Y��S�;a.m[7��:"�S�b���η��EI~
�Z)����J�_
��ZK�D?�?��+�P�'n���n?x����=���L�]%����͐�S�%J������6�-J��| {��i={�N�Ѳ$0i�����-���א,�O<� { [���^�����GՊ냰)�'�;涉�����4Lk�\����$����a��*���e����G�4[�GiZo�q�n�'
췁C��M,��<���!3qq����k�XJȎ^����#��*�uGC�M\��ǘ+����R�d4{��H�z���t��tչ(�X	8�>Hb�����C�&�Xs��?�XY�E�����J�Ϣٟ��Z�i�L�S�=�9D::�'�3:hQW���^�V���0ȉuը�R�C;S�|(��R���-�<0��[�?{؜���sS]z�����_�y�ҿC�O ��̜���ʱpx�˄S�A��s9�;��sե��`�.�C|�A��R��?�;M?��P������{?d�TyvAm"М���R�X���EY�W��n��;; �~�+v�����V�F��'Ac���"�W���Gn��� k�Ÿ�G}%�R�+�=��&����H��|��gmɂ?&��i�J���=�̕A���`�FgͶ����0��Ex���ݏ���]���Y�����~҇� ���ʣ;.j�5�S�]1���IFD�>��uBT������:�$�	@��8��&���Q}W�@u�	=�=@+軘h�w�7�ޮ>��c��Ɂ��i�'��~ѿ�'����O��iȕ���K���x���A{��L��}���.J\*4�2g�6xߕQe����9�-�:J������C�N�����=pt.�!`��so��f�l�k\YW��F��K��p�:�����LhAW��)�V���FL��8���'���҄���&��\����L��S���뗂"=�'��r�]�[ۓ�K��ĥK�'=y,X8+��]tX�V��c_��Ǣ��bM�Z�.���y4�Vg�`����!
��y��Lғ�mu�?ٯf�X�n�su\-�7tF�xwt��L�m�	��6�=%~���; f��ד�]aLdB�QbH�CG����<U��-���j�\�������� �Z�GVm�4R�BY��,��Ƴp�@S�ui�]~BvN	��u�1���g*��vJ��u��m��ȧ�'��4���*H��09}}������E>����?!��:I��A�epH��a��B�W
�DM��yuwk��c��-��:%e���9����T�7@E#R�F=�3�{���p�a����V�\\1S�.��,9d-|���]M�BD�V�$:b�[M��UVO�zp���X��@o�� z�~���[pM���F���l���76�J�>=�z��F=�����-gT霋�-q~|��Y�g�����D�[�9L�;$߄� \�|����`�DOE��eC�q��y��^HnݍhX�OU��%�͎����l�Z�H��d���/�ଌ��s����F���,u��:!0z ]O�r�J�
;�	�L��r�Ro~'�	����'����/*A�/���eZ7&r���_�s�FXl׵��,��v��T���89�J���t��S��q}-tG��M��\hS��;�x]5�r�1U��x3QE�ʧ.�Z�IJ�V()�V-V�9��� �n�JCG_��O7h����R�gŒ�,5y�b��g�q�5v��m>����h�s��$Iǲ�@l����|g�E�����*{�dqN��<�$#���en���\���ˆ3Ѡ1�n+�b($������vI�*����5#+1���M�%���5�a�c���2�j�#Ӄ��V�q���D���9ۀ .�'_4$<���=E隧)x��Q�6u��(*g��g�l^N��>*2k�z
���41v]{M��'��ȱ�����}����CP3 �ƒ�;��mf�r��9��¶͕����,Isժ�*wi��$��-�:�A��	=�WcuT�ck�8.`#�w��U�L< ܨ��&�:t�0�T\F%��>h��e1�1�ӄ��r)x��?��Sʗ�ew�Q��lH�g�?�F�oU�<��O$&�Y�mXu]�bu�ъ�)6;��uh���'��Cߌ;��0Z�P��bK��Z�s��Qҿ7���	�끺�^'�-�l"���J���=���~M �k��*�>��3X�� ǲ{F]��i����!&����D�e�d����&�MN����QO�R��S ��%);=t�x���J�N?�y�RxD7W���W�A�|jO��w�B���\���N���"�7&��m����D���=�Snuu7�N�U���Y�Z�Y��^G���=W����&jС��鄻�xu����$Xy�W��a�O�W��WR��j2�ĳN:G�h�[�����3����`# ^Eg6�ۗ����MO{��;9i�*b��%�t���O������ae�_����V��>9�>�<�b^��B��N��Ӫ��Xܜ|1��~��e�'09�Idc�&��Pu~`�El�R�I����p̼�Y�o��{[.����9����hZ��N�Z�y��LZ�v�Pl��×�tx�E���=<��H;��TU���ۦ�ڍ�w�f���&���%47�n�,P�8���S*v��w��v�H(�`����Ll�2��"5��v�q2�<&*��&�ҥ�c���s�y@c�e�R�6 Wl�Q����������{�t6��O��D_V�UsE���w�,E*~����Gr�a)(K���s,���&��D[�q"��������y
d�֏��O �QIV��s�@#Ѓ|��n�=��,��j�`�r�"W9q)���{+c�)������$�/�K�0錫Fn��ަ#�MH���=����L�w�����i9D��o+$2���v������3�+��"?�+=��l�D�4R�z8B �F�ߴ6Ƹ�®��X��r���~E"�֢�Ceh�挔�E5����@D��##�,s���и��5{��.�vN[u��R��d�W�*���(��o�Ԑ��#�~ r�N o���bl�ۨ��e"��9-SX<��	b(Ia��j�x���v7Cu���!���sm���(��cR�+z#����̄l�$�V��u���A)0'uSσ��I}Z�dǜy����-T�P��t�d�𱽂'
�s�����X⪴���`�\*t?!��bB��
���
��3��BB�}�;�hh
(5��r|�؍�*
/{r^+�$�-��R�+ŽD�|$�b�����ۅ�� ��}����m�8�Ғ5��A�p��{<!�V�45�@٢$E�Z����K}�t+�O�E���n�kz�*��U ^!�0��(V_��d��D-t��rC0e� ��f�E��aRPbǵ-:�Ba����X^ꋎ�?�6�vխp��eg��E�����fa�?YO�"N< T�T][�H`{��L����0#�����pOGΰ��æ�=�b���C/~r]�n�<o��*���Z�N ��--�e�3���⮉֓ď�)F�{dƱ,F��&m/X��6u�ST�����Tʥ�
�!G,����ǟ؛�]"BX�������C~����r��m\I��s�H��p�B�J�jHD8S#�:]�M�<�d<��)ī:�����:��gj��l������M�"��j�=^���Ŗ�a�9�	����o�WH���ρ;�u`9�ܴ��)7M�P� D���N��S��J萧6��^�'���O�����4�3{�$�5Q��\��	�1��A @pr��&�u~Tq�?p
��Vk בz�8�ml���a'ל1O ���)��L�a�|C��J�I��=�
ϯ�=�
�z���}������߀�q����\���	~ٲ����}�H�H�G��+_|� +Cxy�cZ�����F2[��E^�,�*K����Ͷv�͕4-У��`+�p1+N�0�܇�$�"�s�u�{<��4�eC}sOC_3u1^����H/
�{ұ[�8���g_�c��Rj $2�0LSeI��y��Zp��O|>���Q���O�S��P+�07@;�[��$��Ă�u)����A��C_��1������P��V�H�L:&��B�N[�Tg?/ ���5I��̷��x�7~�Z +���"L����dZYlA�KWi��D(���]�{`i�f�U>��c�)<c�FK����v T^��Z�Bi;M?�T)��4�/$$е���,]L����PN7��Q/�������Aᷯ�7!���� 	�&5�ʵ�.ru^��Z��DI�,��E�ҩkP�I�V�e��v4��-�u����D�(V��:g�c#��3��yZ���f b�G�Q�Rș�������
SFJH�"�.�����t�,b��;��r����5䄬�:� _h��DNQ���>Z�oi8�l�2�{G&�3��"��jD���3}�a&����j�|˄�t�ɜVt
������z���V�Y�K���+2��}/�/��Y����t0��:��fI�m�)�M�a��R�ƀ�Q��<'��e-����%�SL#B�U����e'�DRH7o�#�t����3Iy��@��ˋ>JT,���@Inz�-��J]�~.4[�?&昪�wR��C���1����j�_g��=� �x�*�Y�J�r��KMē�Tn3�=�p�����ȉCV����s��T<\�����3�������w��De�D�9H�d��`	J��&_"�#�	�ϰ�LK-�/�V;�(�\A��z����S]f�9�D-���;��wU�9{��kI�8l��_��w�x�7�&�W0��oܴ|bZ&f���Rrh��B��Wc�C�b�s���<%YRYN���P��^hv��|��b.���C=��*Ͱ�yG^h���XqG5	~=���n�Ua�؅@z����1| ѷ�V�{3OiLk�k#�D��(5�9D/�&;�N+9�Q�۱ә��'�*X��5��l{�g�=�UP�?�_��C72B���p��yJ�|�z�������}�א�������'�������rY?kc˃c�L�	� Y���_�M�XD��A{w�)=W����������Q���qǇ9~ �g5(A�Y�^�i�Y��ω��7Я3�|�����ط�Y3G=�w���w��u�!��aJ��'B6j����1��#p�>C@�G���Z#Lo�SN;ἷ���8�-�3��2��Xn_�MhZ6�*W�_4u�]�#��Ox"ֲ��5�÷X�M�uc��ob�7}S��2!��5:!��壽-h�B
����V /MK/�:gsݒ�\ߊ�ڃ��\*ʍ.匯��'פc��~X̳;�@�����݂j-�W��V�1T­6�Ph�o��i�0w$���y{�$U��0��Q˂ �����tR��_�%����cJ�Y�wEye:��'����UUpYN6 ����@�x�>�D�l	�6�_X�º��?�GH�����o�c��+wk��ry�m����+O�����
v�+zU��@L����w�6`Z⬚��lF�G��饓�z���`�ZV���云��D/VO��X�񸟹�8b-Lb�II�ZXϱ�ݵ�Ro�Ó�W�	���k/q���y�Ӝ�Lf�j�f7�Ǡ�eoL�tgNٝ�"PA�Ox����s�o���->ƯƘ#>"a8�qGr9�Mh�X��)o��T�}�N�Cm����(�z������n��J������
�{x���N��mVSk�t�$�\|�`a��n0U�ᦅ/9����b/-'h��_mq�z��D%Qf�-"[Q�>�ra��(���R�o/Gl3��7'7���E�p��ao��:�o�T�G�q��s�jN�p���e��4$�T	9a7<!��7BS���Ug_�$�^'���0��'��<��t�� :���ƹ�]i�u�oـ���)�G��x����H.��I~��{��9P�����l��h��gv#�@�q����[�H�8^C�]��F�X���yx'PO���`��bE�]P^Ho�	z
p��N�/�˿��W1��x�K�VU��5 �Wv�U�NZ���r?�XfM�1�7���Θ�T�݉@ S������ѷ�s�
r6ĩ�~O.��� d��H��g�C����k�
�� ����'/��B��tXW�-M���ǿ��}�=
���\a���	pB���s?��'����=ZV������'�)��Pm�j!~�B>˜=J�i��Ɏ�K��q����s��br�����y�z�c�R+�8�r����I�
O���fgWׇ��o#�e"�>s���F���I��>򖻸V�����5u�ZG�B�2���"�-i�!/N�LxɞF��+����i�<�f'���~`"ߨ�P�`�Z��n&�완X��ùfM��Cy�+��"���J20�J�&I�}?��;X�NVY�i����z��騿�J�v[o*��&��.�Q��/ə��tфl�3`*��aXś�l�C3���	�������ڥF�z���|]���b� �����h����8��k$n����5����01v���6P�	��`4���j��n��e���2{k����GBU�
��^!cQ镇@�Ed�z;���j"�5͞�Ċ�_�E�|�g�#kLN:����L�=vN��3�T��o�1.��U��2��m��!��-�w�0T���%���}D�Tq��!�Z |�4�;���1���&�Ȣ��(�)%ݔ��UO�a��Ug?��zd�b?�#��I�ਓ)6��Vo߻希�D}Z�<����)9�7�9&���㸳�dوۑ�_����스�*���pX�,2_B�+v�}�7�/�&|���U��b	v<���茐wzg��o��֨ڧ���z׫p�t����M�DO�a|�v�k�����F�x>iJj)��y;DF�U����R�<8R���eY_~�r�lso����������t�%��U���ɉ.���5�_�d�����r���O*� ��K�,�@v��*6G��d
�4���}E�U�eb/��V�~��\�l�VS�}�(�$��;����1j�6C/O�(P\��u��q)=�ܔ߸�2�9�(��]�B��
ʸ�C^�+�3س��v����4G��+�6�W��l1��3U��^��/�Hc(U���lnl~r"��w�G��Y���L�����ճl�H)~L�a�����Q���(:I�����4[
������ޕ)v�A��3'�K��CݒFϓo�?0R�N`��
8����7p%rm�[EԨ�4�����7`�o�FpU�|.��e�Q��gq����t̽ع�">�YPV�se�A1�xՎ6��*��°������o���OȡyG		�{1��t!E��򇌇;���/�,��.��S2H�8���]��o$�?t�j�Ah	��	�~`7ɠ�N��ۼB>��H��%�a�R�C��� U;�o��6�2�����!�MN�\�C�$�i=�_%�-�X2*P��.���Ql��rY�Y0�T/�}��� -��+-��Z�(�e�Ħ���ƌ�18�k&���=���I��?2 �2^'	n��5.m�6������P:M?��!GOf��Bq��Q5�+�p蠋��a��[[\D�H^{�h^ݢ+6��.�p�J�t��xqޒ��-x�z�Ëj-" ���pyo�<��Rתw�6�}U��/7�Ug��&�d�sׄ�Ey� �9|�^!A�w���1W:*qU�k�>��rJ�"��;[𐗳����9e���J�\� ��v�o�RZJ��
�B��wWvޛ��J���IM�����%�/��6�����\��I }������`XL�|V�$���O!,�Fl���{`�7\ʅm�������*��y������.D]<�ܾ�P��'P?���/��ӊo�"`[��sDH�D<��P}�Î��b�w4q�֫���� ֳl�����ُ3�ӟ'.=�G^ɩx ���[�양��i�R���#G�� j��a���0Yӥ߽�/��}����ו�L&K�)�`��J�� �0�(�m�L���w�Gz��$u25_�쾸��s
Yw�?���j��>̓�\b�-
�i����hw�6��ؼO��@��m#�}���cgI!=�����i���%L����ט�?�l@͘Ĩ�[��lom�ڌ��t�����������{��P�6�����������X�A�t
�n-)x&;��jB�1砉(4�3��=�a����IJ������3yjQ!`�{ خ��5�]�u������#���|��B3�HUIb��<b�G���(�^��K��|��O�mu�mGA���c�ܞ��E{]�oJB�\�&���W���w�]]n���0�Rb	�������z�n��&{?z���8��z����L 'ɧN�F��B_e���B�`�� X��닭DIT�v�>ڤcN��=Ān�ܜQ-&Ը�"�B��V�O�&��>%�hy�h� �z�.F�qJ�H�ւ��8��=�MYl�5������Ӳ[�w6�I7*Zߐ;��O�9���Vղ��F���ŧ�������9��?�Am�8�~���FLt ��|��:Z��#�����=��l �_�h�������&7N�Lg,���!�)0�R%�JW����jm�r�J.������d&1�F�
���7I��rT�7mj{J�V
A7�(����� ���)�E(d�m��=CƼ��6�v������,98��c�Xx�؝q��HHr[-�5�6�&;������mn��^�nb���������'�v��w3��s2r��T����b���ޑP�>X�r���z!�e���CN�7!�
��N���!�I�=��������`�t�P*k�M��������<T��a�ܦ�Q�iDDv��dG7rtVܩ�1�i����f����*�r���k!�Ddd�g�0]��@�X������k�z��!��\�^bK9Q�Z��~���72���"s_�v�Wýl����q �fpŖ�	���فfm��{�U��#;?�$��Lhn�Q�� W�	@ѵҠ�652LSnrO�;�	���fQ����%|G�I�j����L	���J��w�0�Ke�J��|�	��l��y/�i�����2�hv�LA�G�Kn��3hgGd`�xz"���e�D)��KnU1�y��Ȼu�40��6eB��4��#L�(	k��8�Ӗvz�kTp+Q��Kbfx\���Y�ss�1V��.�x��ĳEI�;pPeB��8�iD�_?���65'�:��~�*����+Z"�ڎ�fx���p�x�KQo��O�S_��زΠ1p���� �g#�E��.52�t�.�Iن��������s�R1]\�-yMe�M����R������!�Գ��Y������ƎMsm�S��n{�"�Fĩ�_��־:1�!wF�O҅l����?�ٞ9�؏��~�x�xt�rl����;�[H��vcd,+^���e���?�f���4�|1�I,��H��7m���S��@���9ظ桶S�ĩq��L��%n��-�&Q��f�Sx�e��ҝu�>��s�{�CBW7P�	� a�ߩf�������?�?5"�)��?��r�4�<|0��2x���ڨ�w`'��#�]jb��7�֕
��Ax�J�)'r%���$IY��bZ��m褮�'@k;�$�L�0�+���$�p0$�S���XDq^5��H�tƼ�E���XF�z�>����-�ʄ��sP�?ϼ<�^��oFA���/�D�s�z{��6}2kxT��_�m��w'�1F�g��N���啑jP����]��#��b���!?׻~��`M�&Y�诈�wc�����l捓�@_sWz��r���C//|�����+�#���V�[����1^v���Y'0'dk|�`Iڶ���}��#��|Ae�g�Yk 'KS�P��q���-=�C�|ܟjwu�%��e��;�b�O��и��x�ӄ��%��0��O��6ʇ�����f�(���^���X�~[O#�nd������BTT�R�<�z]��UT�?��ΤٖilE��N��ٴ�:�^�0cN��]W���\:P���oV��SPA���ͯ��0�U!<߆o�ݚ��2������_qDT�r%\H^Cf��d)��*�v[m	��7BW}�fQ����|��sr�T��3��՛<��i�?������,���HX�
u���(c'6���g�r�ħ�%t�:�.Vp�:	�VW�^�ڥ���`;�,��b픧�;����OIJ}�40L|q�lm1-0�g���z�(�u��1�l�ꄏ�x��|ƈ�{�H7(��Y7�6�s��Q�E�ʹ&﻿���ãy����r�TM����?�M�l�r�A��]�8�B�9� ȕ���<[9�">�3��Z�������X��q7C i�Fv����@���!V@GS��XP��̔W����,�CG!w��+�3�f�ڊA4�QΞQ�F;iZ��8�2{�� ���ʔ�ŨC����Gs0�Ԑ����&"x3��4W�����ؠ|V�lz�qeG�P�.�N|ً�5���j{Y�A��񻀄�`��&p	�W���������҈��I,;vtf:w..�9��v�5Qt��x@�tXۏ�Z;��#&�矍����f�,؉H:�7��)@�裨,��0�{��M8����4+%����*><Ufȸ�r��ρզ��[���'�)_\�3��xP���f�B��=h	༒t|��Lb-�Uș��R���i�mt�w9�9����bT�0+,5�*�0����T�;�ȸH�ƨ@4��E���\7�U�<�5���/�d�u�8�P����O�~V�}sN��_�m�5��1K@-]H�M����Мy}�kfzQ�}�&ӄ�$ ������RQ���SH(9�Že��\��>�}#��IZ�_Q7�#A~ܚC
���'��6?��TS�]�7���S��|�����]K�]�F�q��6�aYZfc�����g�a����GV���2	�vА���Cl����K�q��#�AР�u�!�t�C�S�!A�&�ע^n�{�'HR�p#�ȅWH�
,XK�t=H�a�L���30~4b}H+���?]I�L�;2ϙV,ο���w`gSl��B���J~ 	��v9|��������z�CJx���9�sz��t]�dd�c�{BT��Z\j�9���TT����p�_Ҽ�eq�� g�Iv�f���[ط��iP9�����)>�(r�9?����^�į��LZࡦ�C�缄�
���*E`Z��А�eK> �S��qϝ:��W�f�g���c`�W��kR1ZJH/��^�H���A7�����:��M+�GIe�D�J��OKП���iwMT)��M\7 S�ic��Z������]���^#��*[��.��O��~� �.��0X5
*XP���I�h�%�GsN��0�|0fX���&�%���/<����<�u�gM�snd���r>y?u�8_r>�E2�/�����4�8�NK�k��.��2S%�\�Xm��X_^�F�3!��"�=���g�ѮB��$��O9�L�ԍz'�br�o6������K��l��&!���M��Zt��7ء��F�V��|�3޻=�f�Vβ�r�BXK@��,y7�v˕Cz��=}"�����MeC`�oIx)��$�$��Rz"�JC����#�%ز1��uBn>�o� _bn����.���ޜv�_�<�
�v'�����MY�����<l	��i*`U�����ptU�8en��θ���)�LS���t��	�r;�P�7�.�*CBf���2�.�9��n���o��Z��F�"�?lf��H`��h9I|�V� 
����[�]�Zg���1���A�W�d��7ن�DH��,� j���&鬪�p��,�,W�3&�=uF�3B���$��"oV! ���
��z�)�a���29�M|�U��Y�mV� Z��z���I�8��m�5�b@���Ã)E͚�°^���?�(U�����W3�r�n�	�K�Cx����� <M�a�Q��۱���^o�5[|�w9��
X�B4-�L��?����W�s7�d-�
#�ȃ����	�Q�����������qK��Q�j���5��u�]�P���0��?&�Z$lh��z�d:B݄��!������/'/�M.�-�H�~g4#�i��5�w��G��_=�܃R�^��C�Je;��<���������� �&�u$�t����C�<4��5)x� ��5
ĭi�'�HU��?Dm���8H9�C�n� z���6�4Ф\Ґ��X_�7��G����*�PidK`�O�cc\��/r�9/<Y|����%_�Ѿ`���:����/��0%.+�S�g�v��H�@ B]��I�[����u��|�P����jD�fZT{���Nl���a�p�u�C�&��r�ĺ@HI����G˱~{��Ío������:��(~Nә���9	�@6z�H�>��R�� �>���e�P�<���6ړ%��;�jư�,a�v�g>՝�)�!J"��/�z��/�55��v������P)w�ާ�\Q���DG용��|����c��7� ���O�z�E[5�s�D��+�-Z8�p���^�\5��e^RH�"�)wr��N:���D�H�?�����\e.W�$���ؑ����C}��	��{BS�eش{�Ř�,)���uĨ���k+΀���x��+���*��0�wV��.�FٸN��$��!xM?=ަHaJ�b�=c/G���w}R`�A�B��#���w=5��i^z*�c"�9���b��$H{�?���!:��APh�r���Se����Ȣ�.�p��Z	Ro%���g�J7Q�e�1,UąX�Ӑ��9�d��� ,���L��cg���w��Ƃ2������g�
<\e�E���O��1��4�PFH���R3��0H.�xnF@`�V��9ܕu��[	�?=��&)��;H���tZ�U��cT/�}QO�i��Ta��G���P��kǐɸ�X����*6C���r?AQ]���?���v���V��'b���!��W)�7�R�1����+뤋_g*wkSrӻ�o�̑�\!�U��I��-6��ݐ�߉�ԕ�ڗ� D���w�?��i��?'cfL�Ba!1L=��.�nw�3$#�gӑ�#a�lB5��T]��uj���e��!YS0p{�����>3!8�	ZsY��+>�[(�-����9���d{�)Ļz`AD}v�!�J�=q�}�L�of+�q~�"ɟX���Lw{��^�&<+��&  Ӱ�u[M��;��C7Y<��Y��|�k۫����o T�
T��~���0�>X=uk*��"*�]V��UۑT s�SDh�6����06�a��)a0�p+�&�1sؼb'W���k�Bi�.��V�	���Z�Y��Ψ�QBV:�3�C�+0�T�,M��V p�s���(d�k{�E��i�����=�D��t1�錠�7��K�W��5���օfN�~}���s��+�)I�޴��B"N��,B���S�Ś�YM�Fd_�#��
���}����3@+��Ҝ�E'jo���w��*�u�w6�ۑ5��f�b��wA��	g`$�f ��X�k_G��Y���=�|m���#B:����������MSy����_;�f�d@�S�Rձ%|�	��6�f=�NâB&A8dpNa���~�M��Xb~��EZ�bAw�
���T�k�jǝ� ��:����⡚^zl(�&6��l�J<H��q�;Z/,8���@����+1����[q�M�A�����K���(	�P�r>��k����'%sK`�:n�ڃ�p	��@Z�ī�B8{��(�E���L�CZu�c-����h���~�>1����l�u0�k"Cf�<ƙ��hg����2� F��q���-�M4j.��;�e�2����Ȇ��d�G�$��	k*��Zz[ẵe� �[�*?c^���W)'�����+J�b�-�ҍkOm�O�WЦ�U4*>��m�z:��^��-%�zÔ�)�IR{�N�o��0H�kNל��(�u��c�-*�z�GW��,�Mk��l�Z����C@��'n<��B]��E1M-���Ăn�
��ۍbM� ���,�1�m��O�^� C�o��8܃�t����2���뙇�i�������2�Mp�FHؤ��UAv������\��cg;�23�*D���7Ca�խқ	?��e$t�$T�A�G�=�{Ƽ�~���jny��4�d�Z�9��@B[{�F;�.'�oe�2˳YR`�� ��Z��$FA�,$oZ"@6t�Z�G^;٦8	U9ĖpxΤ�X���b_5ZʴD���h����;[�
�%3��o���&�i!�ܜI\�FNT��>���a--�c�#�E��f>,�J��q�c!u��;��X�x<�w3&��v���uFef�����;�V�5��V�-d�M�W�}O�=����<�d� �&7�̔�[���Iu�u�)��[ǯ��]�}���!1�{T����+��Ob���W9���޶��;0/�����"Vy'�y�nV�ȵ�P�C��T,�" �9�w%�^Bhހ砘�}�|6c�o"p����RWSY��2I_�}�h��)�W�|G�?.�x������p5'��4��=�/� I�ۼpu��9�[�  ?�db��D4el5��!��� �VX�\l.�x�'E5�/f[<�T>�8�G�� R���zƒ���^��(2�-����A �r���(J��»n���mQ��n��5�d,�w��<�����w�X���n���647q�o��3��g���K!i�us������������(���|hw3�%(�����?��&���(a��񇐉�z�Ğj�yV���x}��[�m(-k��Zvkl���x����� ս�W��{-�Vl�s���"#F8�M���r u-^��tc��aL2z��V�N`a��Zokmmzݹ������N��4��.j��V���L+��c}��9�ǜyd��}Į$�֬�g!f�G|07_��I�� �&�W�PlcU�4^Fy�������kF��|Xl���t͓���5���a��C��޲f��3�G?�tv�n&�L� co����h���J@��J}��m$0ĥ�����0�Ym�l��,��%�W�T��]YN<������Z6�~o������nk*�Ibe�EG/օ��U܁['����B�/���O-8F4����}N,�_U�*"R(gQP�X�*�����C��s�e!����	w�N� �+N�x���yO�'�h5��k�b�f�t�b04��M'�ޚ�:�d�Z ���ϰ�&O�Ԗ�Z~��%g����Q��z_}O�=@�l P�JO>��;�qHqF^P��"I��c��hKy�þ�j�?���F����HR{4�^�xIav�k[��Z��Ƶ��J��gOv����9�I�	Ժ��yL<*��_z9�$��٬b5�w���#�ڐ��Cd����@��B�"!SF�Q�落�G��q�%L1�hN�<4���?�#����}+<��C,G�EvO��7����O@����/?������e�b=�s��w�/!CYS�������,-8H���l��v/�F
ȥ���*�1��E(�Vh�I�1���6�؂����R�g��?��1��Fo�{��9}���FB�0�*B��L"K�}����ęз�����ƻ��5<1=��PL�b��0�ɰ��l�/�)a��)g��_(N�]�z1n�*���F�#Ż|G�,t�M8��G.���4ɻǥ�<���h�_���LJ9��L���S`�\?�d�{�n�0a�Yo��H煺�1�!�.�o"�K�72V�!m�!���WH��]kW�hn�_����(���X>�R���7�q�\����Hu=��� �rk8�?w �Fߢ���aa�nՉ��$6� ����L��q�ঽ<<X%X*Q�z�x�a���g���3}�ݭ�{p�/�4U��?:��B4��9CS���������4z������	4gl�,��y������i�c]H��7?qH��#_n�����Y���k]� l��Ub�*�DH�ð�ExY���1%���an����r!淞�me�⾝�J'#���[d�xq�k�Z$.�$�umrU-�S/���l�%К[	ή?҃IA���x�x[फs'~E���Q�R�֓�e��;c$���3i�:�D?�O8��UJ)*�m�N�z����&���.QD}� �G$7m�XG}Y�ӛ ���"/��!���� @D�]$�cl+<��*6��$��)�pж������:2[ g�� ���UO	�H,�Ĩ�i[��FLC��@�Co06�TxЊ߈���$J/�&��M%��V��>��(�����E���[�hM��&�hO<��;�����,B�XXE�6?o�ʤ�e,t��3��FL��-�a��\,#��w��c侥�`�z�f�[<�Ry#��J�ŷ�T�79R������B.:̅չ=b����>F����.�[�E_�;�;f��>���;���X^�ݿ/��;�&L�Gٯ`�Pd�wY+�+�a�0B'�y�Ҥ�2�f*�O�`}7e�QA�����LLD8/cX��/������\ƿ��5dH���������}q���X�ES��*?	���~4�����uˣג�0���?/C[4i���$��X6�p�|���;��`.�����vV#�K>�p7�ĕ*N�OX�CǙ�+���g���28~x�'�)���,�KE�	S��'3Aad�*G�%�k2l�7u��B�!�4>J~n�O���V�(H�{W���*
���AN
�M�4�/�)��C�{{B�a|��^��~z��s��薮��v-]�a��|�)��Wى����ޟk���&@�3���DN��Ii�!���5���*�/�m����{�u����dh�(�TKͧ�N�a��Zc��D���{�'�M�뾌�aȈ�o�E?TA�H���?�x\�ݚ�����&�\UY'a�~�{�I'�S%.(�`޼�:0���{��dp
�NS��@�M@�ip�?�;D h��=ƻ�����[,քܔ���函/E�磡|?:l��ے!�IW�A����x��P���v��($ ��:1Y�q�qH�y�K/#\W�2�WHV	��0=^���X�,|�{���L������ګ�Ghv���f)��;����!镚 s�uZ�o�pr��g�R����������&�bZ��W����92Cul��.��oճi{�?�
�h��Ȼ����D���y�b][���YiAYy�j���K%�����k�b4H��P��� ~x;� Z+��
Fta�@Dy�v�b������4��8
�EĈ=�񴳸��,s% �e�Ϟ=0�4�8�%�JcRO5$�3@ۃh�9��@]a��!;� M_��`H*:�z�[2���7O`t�C�s���=
�����a,>�ҩ�X�2[��)��K�
���A�|���������z�;[m@r��ւd�_:������tC��RV�P_#���#����/1v���!1��u#���ELX�o�WMs�Ȃ�<elJ<�w˵ʡ��FQ��A��o���@߰��ɛψ�C�;C	��.79^��]?j����I �/�͟R��4�a��M�_�ͮwLb�I	��W�Hh�ق3�!�a~u�MK1���PL�+ue�6\7���c��3<7W8��fܾ�I�xl_-�{��<BJ��U�r9j:>���5@�>�y�{�ӷ����*��W��Z���#,�����5��z��].c&��]D%���b��5[֦�i�~� ��	��\ C�yΰ��v�j���[���ׯ,X��vw٥����=�.Z�.�H�~����4����ڑ'���DhR23��1�d���	��<X�?���J��vn�����	݁� ��W�1&T��B./���g���Qǈ����B	z���ԑN�u��\�/�9��w79춽)��y1H��O�&.5*���Ĺ3�s�w�̶E�gz��I��ʗ >��j@V!�Uz\�B~����%+ns���t������f$'�a��/h93���hfR�+D�껚�{�����������������҇	�[��㡐cs�'��q��\\`u��,jkz��rk�&�
N	�',Qc���::��B��B��}�~��$�+�K5��htj���O��E�vf�* ͠e{�f�-�� �j>\Ź[��!>�R�&Ox����D��y�hmk�Bv��cc-��Z6�=�:%xV1��ޯ�ㅈ6��k��ϩ�b.��f�5�	j?x������3�=�F��l�!)�cL�ג�'��KZt�ܸ6��h׊�U�Hg��!�<ZU���P��Z����U3��pu1O$����HdQ�!�.^���5af���0&�8�n�!S��Hy��jT�u���h�{���r��BBD�G�{�̰�-̄�>���ǭ/���;hg�YR���!��b��k>�1�1!O��jNJ�U	�>ʸPtA�7��R)'J��O�_�(�C��+�H������SI�Yo�(�aV�Xpq;�`D��\p�)e���\�xC�\F���;b�-f���V6-6*���.E�G�iNk'JP����)b�#�'L���� ½�6T��e��6���$��|��L��+f�Ֆ�l�=�S��y���p׻g"+�������v��r����ծ����I�|2�F�V�� ��v��~�G���̷���rkm�����SXf"�y2�䃯"�U���x����;��񟔉��Bƨ��_f�V6c6�ʤHRv�/�L�\��R����~�fa�bE�j���BD�F�ψʅ�oi�|A��7�NxۄX�˓��$:x#��U���-�%��uծ��{9.W ��L��f��� ���b	/r��mR��b�B�o���#���pO�O���p�`��7~J�T`�a������Nճ�B>�KR�ŦC/U�%.��M��l�/J�X�9Q���yT�u��$��qX���<4��ޠ.G�tH%Q�T@S}��8�BU��r� Y�+��8=��8g�+�K0	F��T	�Y$�s��{�ӊ��=&T ��Mm���R������Ůx�`�����7�����8�@�d��?_D0+���{A���ܺN٬2j?a���n��}n�,U��J�B��[y��]�U�7v&sU!V����P�������B#�۱��b�6��<��ˏ�a�(�{Q��lxn�C�����sɥ@�9���:?�F3
��6Z^��r82�i �RDq��S�GJ�&���ϩEH�:�^�[\�=sL��8Q&d攮���c&���9�0d�k��_�����[��g�{p}jo�nB�9f�A%��BP`\Ώ������	9ͩp��or�W��c'�z7�kv�H�n�0*P�ͪ��s�ɳ�Y��
g���<�6�}�}>���gsN�m/��κi4ݺ=$c�d��M�8'���.6�2�Hff���T�kX���Q�S�H���;n�E����:�Q�qT���������N?�B�+�aMQ@X�"lG��*��b������t��F��gȕ�a�`��,a�;�����1u�����WXWݲ�
�h���o�HK�[æ��=4%�_>ᨥ�̈�`��K�v� ��u�f�Xn�w��� #�wp]5��|Ҕ	��^�����Qg�6�l���#���8�� �H����+���=��"�C,��4����k�r�L�Ք�FeQ��I��ш���l
H�I���Z�h�9L��#����J%K*	}� ���ߴ�+���yGN2g[����@��J�2��7���=���ҟ-`vm���Fqڛf�OZ9��c�x>,�9���E�`�祅�;��6~q۱�F�&ő�CR��K���<P�P�-��ùQ���ʱ�%Z�RHM�ҏ�ӌe2�",�N�5;Iq���o�eT��.0�?n8��i���X왴o��8pV��۴)�[�"_m�>�|�<�g�-1�?rPB	����3�V���2�k1��j�%EhYr/!D��V�`|��!��RE��`B���P�����2}sф!���I����su?����Q���S̍��˗�h�i��I�������*�qژd���i�/)/��\��[hd�!�G��"�D���5����86䨯��������9w�O�UQ�q�m�--^�I�>8�O�L��JQs�zU���9G��H���?�^���m�}^�3�?\�	Ү��Xs���ad�\� �f�)v���D4g�h�k3<-Mf�Z����;Ȁ��ls�v!dR����c��J��~����Ī%���<�XjPG�Z&f�$��V8��<-�H��I�0u��i��WC�Z-`�c��\����K �1k�>����~�G��,Lո��~�I��s?U �R���K� �������
nї��+���s�
�)fTJ�;+}�x������'��^��|��=���5Et�������ND'�:����';,�(ߦ�-|� �%TI���yW}�n{��be��wJi��V�+4�8m��"�i4y]ŗ_�/0뻙���?������zk���5�A}t@O��hS!��݄jSV�(uX�78H��L��z���Y���("E�Dtۣr�r����^�?ŮaY�׽z�y@��w�>�<C�ƙ�Yx^�h~�a���&�*���g�
���A�£��'
)�С�t��L�Ö�A)�+p�k��i|�u�}y+Säط�]U�*{�"$Ҩ������V=�Ï:8`v9{��u?οk�;j,	+�_:h�!�qoΐ� D�:.ડ`klkRC�p�ב��6��E���z��ߧ����	u}���if�؍S��>O�>�׈������n��y[���gK�燲�W��F�~������0�������KR*�X�X>~��5;��:�a�"�=N�����Q����| T1���Zl�8��/�Ρ��\y���"F��0����#��Ϥ`���9���܋�y� 2Aڲ��k4�e߸��#f��F��-EYu��&G���m�cM8:��?܋�Z�;�y��	�2G�U���عWPS��MdKUif�o%
�lwԘ ��䫯Cp����>�J�lD�f���Oڸ�[��uߗ\�G�;�ͷ^���A�^�I�������eG��d��fv��%Sb�����X������<L�	�����ٔE����Hg�J#��Z ���'�����:���灢=&f义���-w+;�4��Ґ0|�h����t߹8��]����f�5E"	�T���k]doo�0��Tt�J��I{&f�wj���*"���ĸ�A)�%$C���ځK�Xl��#�;8��R0��p��+��.7�Hf+�=`9\'%0���JnIqT8��Z��z��/�.wmQ�T�������qW_�Fi��A�p�H��bq��rfC]���-ِ���SJ���HeK��e~�*��N������÷]�I�SJ����֧,�(��wf ��hy4��T�^ߍ�S���E��8I.�}�b��
1�J.�<�y�]��AD���8]�J�?���(��OP�u�*�zZx�;?������[���ҳS$���TX�+[7�t�<9@��"����H:n7��]l+\���bi�I�J:_�R���9��\zQ��t��=���1�-��I�Uq$�]�ɗ�3���Nf��	�@�G��?�Y�k������8����Jd�<ߥ	PIe� (�~Љ��[(���6���^��a���xR��R�<�rc�5�@�!N���m�K5x�XhǛ�Q�)�^��M ���W |ǺX`�z��V�m��?�Y�8���ց�@���b���oz�!^}����j���0�'U�U����7��1�-�4����Ј��<��jD&�K�ul>z�Z���H���s5�΄ҀY�
<g}FO��,+�ޝ~���SG.>$�gq�/(��Z1 D/J=�V�}��"D/&N������m��-�O~��-�U<Z�'��ϐC:�wU�dc�߭�pX����^�4��IGߥ#3�څ1Z�df?�ed��/��|��p�/�/�w��j	G>����׆3j��!�.AĖ"�><��!�d�xج/Uϋ��~��Y>�����Ayd����
]*�g�P��|�%���X4��:��wd�t
 �)���~v}���o�aOJqΙ5�֛���PE5��S�j��3>���O!�>�JU>��j,J�x$ln��3"�.E��%��{=��i��Ť~�7����"��Yq��נ�%S�[���b����.�J�Y1R����h�K�P�b��[��T�I����b�GO���<U%�n�t��/+]�W>��v�����Q�~��HD��{õ݇xy��*<��s�as��Qk�NK����m�#��ɗ*��
fQ��_�t��k.�hU�фI�	��<]��.��"?=��Z\��� i�Sr�`��&�-M�F�
�s�@���6�<8��V��
qZ��{`�2np:�B�S�A�(�4\�EH��2�g�J=Vٚ��~���*ZO6��xN^0��1�Ki�n�rg�T՜�����޼��Tzb�#��2W�A�5f���`rO�7L��gH�c�{�� �w�-[���qʜ!Vݸ���(��ظDs3<�M��7jH�l�	��S#�-<[k��e��١W���=|
J�s�Ѫ���?񣯂�&��?�n�	g�ik����O �9�����t���? }$H�U��ꓹt�F��P�VM|�5��8�����p���V����k��>�tc�p�xA�_I�������f�-F4�	O�\3�{XڂG/�)u�>_�ߺ�T��7b|jN��'��⧟:�5*p�-�&y����N�(��Di���g�mw���o3�p8���C&�/Y'~���v(�͊�ј0,U�ޡ�g죨��\�h8�����N��!�Z#�Wn��x9�*K3�z�CzK�}#�c�*KV��W�;].#ݜ�P~��0b$��#�8�8+)sj��i�'𹋣�O�����2@qQ�K��`^�v����;��b�s��2y�c
ߨ�����ϐ���pq^��<��mα������>�ݎ*(^	�X:*�Z�v|�G�����Z�J�Y+��hׇ����q'H�Ip�a�YV�nQ�^�l��Y�֛�hL��yol�W+Ou�+�W����POf���a���S�
�o������"r¶�YB��t�6М�C�A{&����n5=�1a��a�]���NiF-���g�����R�����H�!�$�,(�<�^�f{,}��͜���.�px�s��ZR[�M��b���
Fcs�}R�j
�+�U�ѯJ��ر�X�v#��]���h���M�}�:�������g����R��#�,gۮXD�}ou:�벆�^��3q��� �5F���MWt�*;�1�rAN=�'��]���\-��A"r���ݬ�D݋ �dH�ݝ3A@���6H*T�}t}o��ت��-U�#�:�V	AM))�)��9���W66R�g6�Z��*3O�أ�r �Ph�e%s��8�˖��}��c��"��[(�͗ߤ�M #�K�bܗڶy�i�\:���	��q3	����	u.Go$W�w�0���.�ǩ����f�P��v:i���MA^ 7/}����[b�[69�ejq���� ��u�%���y��'a%Iaig�����F&D-������K�[X��+��D G�iY�w��g$�޲�w�Rg���McEE��6Ey��9���O��h|x��[�}M;���� ���q3��~�L�.�K%�)�((+.v�(��T�����A��t*iܔ�G�����>��T���N��ǋInC|��e(�02*�[�ǟR���;T��c��.\q��/�q��=�s�fX�*"��}���8d��K���ɚ�zr��E�I�#��Z.S����HPd�@a-�0	��ylՐ�D�PV�U���+k�N�U�*D~g"�m{�K�ޚD2�-p����zZ�r�'sQ� \��97lC���X���a�uP�+Ȓ��S徣�H.=e�:�O�rV0�
fe��
�WJ�Ũ/x�tRxf���R?�V��	â2�E~B
&&�G%��}�=R��	��M\��������j�~ۃ��,l���>��<�<a�I!�T��o����T�w~W�4�!f����>���:����x�$�lۭ��x��� E� �I�h��^j#�?|�2N�4��RAT��������݌齳=UZ�p�E>;��9k�X��X��2�%�G���8Xm������0B�QI��s�'�c��N���7r�̍8�Q�H$�ݘ�A�SXZ������aU��c&������b�̺rHY��jZ߇y͋{�����D�K9r�`�C�.s����\;_DZ!7ڜB���*�7qS\Е�����G��h�h��Xg�t�2�q��9}��o�G���#w��\���0��d9;d�+�_/�=��V!�A�^nn`��S��*��=�=�p�������z�M�x��B�+��-wl�d#�g�೟����.�i��՛x��P߾݇>����UW"�sXwS� h�{��5�臿s��yȁH���'��-��FR�cf�y�I�ǔ2�q5�t
dpq��"����5���ct����20bM�ȅ �O`LJ!�`���s�y�a'؃?"O�0f ���EJz�������v��q!�J
AV����'l^���_4��Ϝ���8*�9��+dqa=}�b#����#l�,�(c#��4e�5��gqP۳��o54��F׺�P���F����Ի��!����D_���&Mr����p�}]���~����i����8t��AA����JM�m�7�.++k��C+���!y�?��#��EPkp�Ng. �*���FLҝcC�d@�t�IwI�W�U�*�"(p��f��gsp�X ���'x��H8�ۈai�oǍ�6�'��e��-0�ڃ����9�O~�Џ�%[z�[W�	 �C�E9�*r�~r�FÅ
�V��M��ڐ���(���eUez�'TƸ����Z�����+�&��YS:� �#a�X�J	��0T�eD�G~jZ�ILi�qT��U�\q��y�V�L���l��z�ۺ��S������W��M�b�j�ˠ֣��U�T�](��C_B��L��� �^1"�s=e��8_���R}�m��/���9&����yM�2���B��$euC�@��!e�qkh��9Ҹ�M���a~��m�q5A��x@z	�_�O�nCsM��	M��X6[�����%�u�Ѫ���;�
5�1�e�T��p�����?P�xX~����K=�񾅇�Л[��aپmiU{dD���ꕅ��+��F����`�j����C�P@7�5���~i���)��J'SOa*�S��5��J�� R�d���߀ף�0��	�o��2��_?����+�6ҡn�9Ift
7�*�S
[��Z!z��!'�@֍uS/�xvC_��&1o�cK��Z����fЂt4��J<j�{��K���C��U��E� ��,I�����gKGp��6��C%r���B��� ������X�=Zֻ'dV�����E-�q�A9���A��c�+�i��羉n��]d0��{z�]-D@G�Z�*�?�êJ{�!�$|MNIa;�s��B�1�Hx��y�1�o^PB,��k����x�'b���Fi��Y�C`F��i�'�l;KX����NK�4 �����'���ʘ4��1�Y�>&��aށ�9���B�����;e*�u�a�:��r�4E�˧N_X��Vdg��棢@%�r1�k�#�(�n�P�$S+T���V(���B�	yoi���=jI@2dzq�uG���T"�90tSmI; �a��V���:�R���ȣ���}�S��Ibj�E�vnQz{rߞ���(�o�[������j�]���7��x���0�N'ҭ�����fcl��F�(��_�?�؁���=j�ԣQ[�)?S�6�~Ҫ�;��m[�V"�ڃ�;z�Xg#�6�W���,Dr�'X>�{������14S����:� E����LWxwK��2�-�H���Xl���?Li�&�t}t��Sݰ;΄CJ���F���V�ȡ����� ����ѐ��Ǔ,�g��������εB]�X�}4�q.��.�d��ߍ�t�( ����[/��Ô��Hq��q�*�T��PpFI�d�1�q�rp��^���P=Ҩ�^ӒD�������p�z��K��S|z���c�]����ҷ��F�U�2�Hg�Mĉp��@�6�͘w G�����KD�8�~2ūt.��#�џ���ή�{`#�v���G�8'\eb�od\�sڷ7J�lj-��:�6��	�ꐽ\~q�n�v���mFx��KBF�n(�{4�e��r�Jy��IQ�4�t8�@����k��x��k���Nz#���;�NfH�?.X�/����;�:h��j>�V�]j{$"4W����q�8UJ�~�w���K*3y�6$��*�8���x�B&H�l~�<�y����f� �4,t1H�_p�j��d�P�?*En��o-)�	ސ�5W}���*^%��":��t\zaw��� ���N�^N��T?�_���2�:>�������3���u�2���'��l^��Sx��LlmR%{j:��G'�E]��_�e�|%It�����m�_�SJ�9��wz�O��&>'�!F��[�C��a�n��s�i<���:�o"]ysʦ��� iy`oJ7�r�"��.��_
�_$R2��?���v�4��2�e%s���qJ�I%I�Ӕ�������;	{�R��!-4�
H��I'Hd
��j�G:�j���.h�vw��Uq�0�:���Un���,��B9ꗚ��CƖbҶEY���k)��1��_��Q f��w�}b[�m7H���Q4h�O��Cs�[�^v���JֻIR�v4��GB��?L��h q�4��`lD��$�ϊ��Y�Vn�0��8X��[U9�7�lB(Ȝis��k�����f�~�!�	:=ʼ�OY�#��ȚzWa�z6����P/l�]b�j��0����;>�x���zAW;�ɪ6�ʄ�5�	�����W��PW�6�T��%v�~��).��0�����m��E�0R�}ߞ��ɂ1'�O���cy2+ʲ�Vr��٭zO��ɰ�d'k)�g^���W�jF�B̂��\�!O�ۭ��R�ӟ�
��&J���P���!Ђ�V��/�CхA�$1Gh#��)|�a3�o����]� c��D�H�g��KnLK������=���^=S���J����v��3���JJY��4�w�����"��%��͸�g(��H���v<���Hmŭ:c3���[��1<���7�Jm~�bF6m
��V�+e��[*�/������'�͸8�K�J��?׵A\�|d�'���Ĳ�SAA]eY�#�N��w�Rj\c���-__;�1 �X���P��cj��Kڐ�X��~��$����.;��- �G�IG����v,���s@�T	!7�]+�{�R'�( ��$VBs����4���:�� �kJة�l���A��~�M�;�ˋI�ָ�7��U�f7�;��E�ɪtOR��h��KC-I����_�����\�W�pX�+0�_���L#ܳ�w%���_�Ug��ʮ�"��J'�2@9�Ƴ[���d��fj�Ena��)w~������_{����d2��$�{�I�Z��~]�4��]7�����V��&�֍������ԟ��o#;�c:���u��j�KbA0[���H
��v������,�LC�z�[詝K^N8S�����P���aز�գ(��rv��q$�m�~L���➪G��4:,���:gF�|���?��7Pd�/���uOI��.m� &�Ċ���k�c���8sMΣ�ϯO+7�e�
���`%M.����J��<�gM�t�d������o�g���p�v�H�	�*ڲ�?�"���I5SsKӗXިEJ%6�u}�1Y���8�]��[o�R�������6�о:����&�,Y�
�HX>�������D�䉅�.�'�&)=���B|�����9�WF��.Ǥ����A�C`�M=���u�k�d!���vjo�hڳ���n/�Q��^��^9[k]=Ǝ�Z/*�sE�0����0Y<x9M�[y�!�毥M:�^���1�'���v|�_?�k��8��R0c�??�S�i��)�� c'}B��$��.�q���ef�\L���j4��/�"_��nѩ������P3^E��K�|_�A�4��Uϯ�ݚҤ9�o� .����Y�$n7'q�y,�:�a��ip# w����UՌ3���p���C�y�X�<��bt��ETc�*���F
����n�nu�`��r.�m�T�!� x7s�DϾ���7!#>��2��3>=\7��UJ�3���A��oM5�m��� 	ٛ��[UU:�͎�]a`���Ѿ�9J��{�W�ܼ#?o�H�	�C������a��ϒ��W�����yݘ�R���Gb��E)Nmؑ�n+$+����m���3e x�v*��Ax�����[:�4|��b֎�0�5�/��soG>!�P�|W�i��c��������Χ���y8�4���C�9�Pԙ�K�31m���vP�2�I�,#V��0TH8�Y\&bf=#'��s��2Q��ǧ��-���2Y�Oq�X?��~?H% #!�̢,4�LVe�d[� ��{QS=k��M	�j�s'VS�Ձ3�vz�,NE��5 ���� ��q��LI���a�H�pi�kg�0�kL�j�̰[���$�����wƘ�W�н�l��h�Ġ==�ܿkdx�T1����\^Gy�L����JH0D��X^�~���yGUG��}�&�����q%���ʢ{4�S�k����?Kֻ�43[3�O��~��uv�����/i�r��� "iҗtws�פ�ʥ�R��>���qA�6�M��Zkb�?�}*�w9I?�rj<�NteƋ��X�d	���j�Z1���6��vzQ��T���&!W&ā���(�i`r�1oǑ�Z$��cC�U����ƨ��i_!��$#���&��~e�*���)�β?����h'$7�K�w3�J^O����'�.�.��F���Mf�t�H�+d���T<3y
څb.b�ɇ�Fb���6���O`��P�w�@����$�Ԥ�|P%��YL���?������m�ԻhR"��g��xܘ3��F��n�p��t�O�0�������U�至��O-�b�iʛ�H���� )%�FMHm� 3U�Ѡk3������I�i�4D�>P9�&�3z��3c��(�XNi(�X����=+jׂ[������Ud��s���M=���
J2Fd���* U��2}P�,���O��4ET�'�&[�-���u+d����ڙ#���2�.٨W�<���YJ�RU�8�&������٭A��E�l���)���`�{H�nQ��oz&�,/�h���
�� ��d���c��&�5�񞶧GѪ#�.�Cő&��`-�6u\p�[E�(#�A?/N�2k̒�Ef�]��b��\����N��ϟ���J�a0�-��{sp��&�Ť2����fNp�n��-�W�C��9�iǱc��仂	b\h�w�bs�˖���F�����<��B��+s�u�ul�x��
��4,1	
��x�@�!��>�m+�oM\����=�:C�i<�ѵ�<(�[j�%Ev>An� ����ͯH±�����f�е���W�G�o~S�ky	����B�Z��R�g9wL�e��9	���2���]0��z-@�0?�&���؉W&T"� �qE�o9��Ɩ�I�m�|���h��BE�s^�� �>���n�K�����q����X��?�]bT�� )��$��~rAq�C���!��^��]oo�I�兖����}x(��Lɩ�W����$_�v�xjw�8P�ٸ%��u
���=�S���{~]�׼"��)�u,�n97h��ĹUn� /������{��8�$Y�����A�P=��	�{�%�u�#�L����}�vMytU�]���zؽ=e]Hʟ(�$�"� �^�EN��%Ί���XYDөܟ��S|�b��3��^��]ȏs�ͭ��*�v�ֻew�
�:|Z<��dǸ���PYPc�J>�_C{�U��b}��ƹw�,А����FM
�m��:�S�&#u�6a���z�J^~�YQ1۷�v�z/���:qg�9�wވߚ�^��[���6&#�)H�E�i��=����
z,���{�o#�g'�{8ZU���R�E��h	�
���SJ��'`�E�����F��d��b���Cd�q���y:Qb�l�gC�Bğ�$�f�nC�>��]�9���=3�m�d��}�.Rs�_��S��WvQ���A���V��%s0m����&�R��UŎU>���D�ߵ�]�[�{������dyZ7^^�q�"�4z��m���gK�n�θ\�a���/q�0��z�z�H�SW7�ʧ;Fp�}�s���g��� �1���jgF�œ�ё�w��$?������p·�/Ui[e�,uŻO���θ������b®��;��惁����1�}/c6���'�6�7y��x�M��V�*��X�b`/f�f4�W�Q�����\��#De�@��v��7D��8�$d�t�ݟH���q�� q����D4+Čd=�𡻰�7(�H�=I��M��A��3�O��t��t]�(��Ƈ�Y���6��c3k�*��Ў�b]K*1�l�pbuelBU���酨;!�ϻ���<|���)���l�� Z#�?������FT�[\��i}��/%L)�������Sk����<�c�򴡘�1��'X?[R.
��TT��>8����.��3����4��w!��W�+�b+�Iw�j�����ͦ�V�'f	M)���Ȗ7לp�rm��yL��6�b�����"���D��YPV��:�2�V�/�Es�="I-4�������k���Y���Zժ�v݉��Ql�0j	�%�3J��2���f�jT��P_`TS�^��!|���D���4Jq�N"�ʾ@���%s�^L�t��^��*�Zm 7�
��+zݻj��}��	��ϩE�gֲ��@	SiX{C���(����J���M"��؄���y_^�0-�/��¹b�1
3$sn���Ա�.w��] ����V���!r��%(GI��T+k��Z�|Q�㥜fp ��ο�D�b|�h���z��K>�w���ɽ>ݜq%���4ɒ5UP��h���.���Se^	��U�n]$�!�T�Ge��=%�R��|�hAu28xd���ƘgJ:;HX��8�\���d�) �ڐZ#�����ɠ�ZH	jU������(���:��[�_��FWu���>[�Wv�k���)]Mo�`�f~��Ӈ�Źi/� �%�/ǽ��W�����1w2û��0��~�A��J���meGMAA��[K�'D����K�	tpٹ0��.v�s�:e�ccH�L����;�?�Ɂ�kTqg�������j�Q���7HE�b��'���7y�RI����c��6���}~���ǫlS��y%b�%�-=G��x��]$5G�K])�x�sNl��i�X�6쭷�y��0��
'ٮk�����)��P���%�!l���a��;2��/!J�a�`"�f�_�7�O2a#g*c�� 4�T�J=<���p�St����)��灹C��l���OӀ���)�'{����C"{�h�)P)`c�ߙ���t�:Z�%��%W�$�	lHt���A`S@���W
�=o��_��N�����Xf�������0�(��U1i.!!� v4X/7?�d��?W�Xj�^8�<1�ً1�ܴ��7��6^� �!�Ԩ*�T �s��Z��4+�g��j
�A��G��"F��" ��q�s
�ɇ��h����C.(k5�����,�|�OܴVktB��<�9|VL�N�r<��/T�'z�GR����%Kx�v&&��)�{)�m�X�v�v���'MME��˔l(�T����%��� �x2~e(��\IÇr��� S�-h�����	�h/^/;r3�8+��|9��(fz$����է���αKZ7�vq�o�G}�"���TSxgF�z"M�E� ��
���	�c:#��r��$��`x�Ω��cBYR���Q
V�$��M9d�&\c]G�S�BO�Y�O���e֩:IuܹD�oe�W!̢-��ꥹz?�sE��M�M)�T�^u��Wrv���:�at���'@c�B��H�Ή�|Mj -����*�I\�9WK}>:�j(Tb��Tc�� ��ѷ��9v՚�,q�xm�����[_��IY��E�����(Y�q���ɹ�I6w�J v�Ed�����ƻ9]K&�`�E�J�P�bNN�X��<2|e� ��mYv5.V�d�0��a��3���`ʧ
m��|�Jh^D�ڴ+�lQ:�kU3��Yk�������nrP��A;,4݆��yæ�5=ȧ}pi.ظ���#oG��X�c/�$�c�R�0S"�A��Z�[���'�oū���UeU܍FN:���E�#1�ӧ����:¯>������ߣ�*�h�G��6��<	����i�H�.á�!.^��ԥ�<s��,,#'�O�T�Fr˄ :0��#R�̃Uf³�8szg��;oJa�7�ɆF�x�t[YGʸ힎�v%zbA��8~��j�Ե �O�A$W�>�lX��[�T�`hĭ`;�T��9S��ǋ�|�A�uD��5&	�vPB7P�Z3�Z��ں��_B)�� ��oԨK�Q�)��L�������a~]X�w߾�_� ��dQ�ퟰ"��lڮi���ӊf.?DQ�_�e3���ؒrf%X���t���'��/�����L��]vn��5�l��q�]az�&��01�	�v&�BR`��Y�>k���ލ��XcL:��P��K~����s¬�_rC29��\��dꊂ?��H��լޥb2����"Ͽ2󞖤*5kդ�C+]Rv���lmJ����|�W#��ֈ��o�trCgU-
�^�s*��8�׬k�i�)�L�O������G�5�+�,�#�p^���X�-���l���o��� q���h6A�
j�-���=�s�VU���&V��z!��Y҄�˙'?4\l��=��J�?qM���Jb�e��t��	���7/��|4(�7��}c�#4�ֽ1�@K�#.��]�ڞq�`��χ���R��Sj͢��k˵(��k�i���I�8<+�����6�>D
�5`��_s��e;�/�+�VK�7ygw�js��������4Ζ3߉M)�C Ď}���@w����i5��k:��F%������u�׶��m�(��yw��4��,cҮQ�f1�9q�����ur �?EE�/ƃH�r/����3�V�~�^C�����E�����!�^��������D�la {o )_/���i�SZ�k�R��z����!�$rk�߁Ʋ��Q����T)z�a������v�qJںm�����F�э2�r���#�H�ҟ.����8i��c��W�y��~n)|�i�6̀/t*#w��V)���(���=��2x��Ь��C�vNH���?������l�%�@H>m~hIkЊ))���G�G�V��*��#ۏ�v�h�*�f'Flr�q�u@Ճm�u�/"����*���h�0�R�n�&�i�X觺@b�]���w�
K�. �䋑S&ϣ��	��%�I[Bo�C��4��=F����\��<���}!���WDR@��HA5�ް���YYYB�T���͓���� (|�;>�@5k�m���<G��#�c"\��#^�r���VI����t�t���^y*�]��s<�0���T�T�`��=�*6{^H�����j�KO5֎f^��>��Ĥ��	B���s�.����wj��~���KHR��Lz<d<�;f�ϲ#�>�R���t�Nx�I�a��=E����<�x;
t�RH��! �w�*i>�:nU�j{ˢ;�W1C����:������'��N;7Ϡ�plq�~�Nt�NM3i�%�L�?��#�/:��g�˥Թ��*@F���i�ݨ�>��f�%,-8�/��8S͙�'X��ڕc�k����l�� 6;�"����sD/ɾ�Rk*P	\��G�"�ؐ��[��L� ��f�"���7茴���j%�����8Y�IlW>|�
$�v�	.�u4�2R5,:�S.z�߂{����O+~g��1�eA�?6a1�Z�ŋ"�	���M��#�E�q���;@���J�v��1P歾Z��ne�Mb��� 8�%��"bWE�)fkb:ؚc<Cn"� �	�P���N�;$ݯ��}tE�~�٬U+�m���,b֣�����mY��$P�f������ゝZu/p��&6��g�+�wt9���w馏^g�@d�$P���q�G5�`:��1:�=�QQ�9^�
o.�M��B��=~nT}�1!6�Y��(	f<f�˙b���~�9Z��X�-w�Wgt���,����r���~���*��1�3ݽ�2K�����)����ix+߬�iR~uD�[F�t�Vc����,<ͧ~\.tS&kW�y��+��D�c'Q#��3������yiV0��Ɨ�)s?7:��]���[�4pA^�Y(��[�Zf5�����qA^�6�A��PT���g�VR[�~��1/^w�JM;�䆣W�]󝒯3V!�b�`�D��T���l["�K�[X*�����7��$T���à��X6}t�b���t�m�k;�o���Q%.ĉ~�ꐢ���ܜ$՞*����F�
��g��U���8U��{> ]cX&��m�P�:�Wt\�I}�W�h�
����X�Y�/A����~���-"�\`���aWJ��b�%��"��<.���7�ŌzV�)Gf�[|
�����I)�wR$/l�m�=#��R@���ÿ'te(�ǥ�^c�4 ��(Z"<���ގ��4fy
P���q�� ��)�͇u2F*I��^��!�T�.4&�b����u��+:�7iY�k:(�,�]�7X��=X���w� /͐/W'�L\��j�ņo�zᅂ���2�@������N�W�r�h;�e��p�s��n��h�[f���ߙ
?��/+�so�}h���+*^����vBe~	�ss�9¢#�X�_�ٗ�%񐸐ېP V��v!{�r�3XE?M���	���+a5���/�d�זt��*��f�Z[~P��#0R�^/� 7��A��KnQ(u�+����l?T�砐�� �}-Gڐ[j���i��K��X0�G����L#7%��������:���'L1P��^�Տc#"'2�p�f����-�߇eז��ߤ��u蜀:@!����ܠ�$��^uY�O��G�+�Hχ�|��})#�[�o�0e^�ܻӶ 9U:� q�
��z��`�-*h!�����-o�3<����s���&ZXz��6&��0�S�s�0sK�E�U"Z:�Z�L�i)D~QzIt�7݈���LOpu�����I7��#N�g�I.@y'���k	��Z@A�쟷��_MA��"�y ��f���J`?��S:��L���즲��
���K��jl���$����Zq��
��餣Z��u��/����z�UGm%��ba�b?\�7e�Q7�{�~ӷ#���hgT�r�&���)�S9����
R�r������5��A�`y��p�\	�&y˳�)K)J�U�^{~/Z�R"���|�Η-n���s
Q���?0ٚ~{���ŏ&�"�ܗ*��VmՑ'��W�-���>پ�ʩ}p�=9�؆��<�Xs�ctјz���O��"X�={�s^%Ci��)K��QC����=`����HB?�S�ڋ�=�KaT7�K�����c�B�j���(�z��Q-(��>�uJ0��B꟥���{�k��q�no~�<�.����s@�ڧ(�J��韲.���q�$�OY�l�]G����o��I�S�_ut<�t.`��R@���T��CoZ�����2�S�o9�|�Q�z�{�.zf��&�t;]��͌;t����1�����=n�(��ԡ�:%��4��E_�s�l�	��!�Su�P�N�w�ߢ�ߐ�9��ʋ�u���*?V��8<�ьض/���D�f���Q���͍Ͽ��
����mM�(x�łwR��.�ԦFIzJ9WL�k�jK�KG"d��j��CL��	�v=2-$�e�"��yC�@
��� �A"K���,�=�zE�H��<�iK�w��L��Ém��(x����D����ɛ�'�	ԁ��f��� ����_�h����XY�iVgԔ���:��Ķ�R�o�ɣv��IODa��2:M�X5�/��7$q�ONml;VJk���IV��B'��{��a&�6�M��ڈ�ۙ��vE� �������%��:;���O�)Ċ��g�W9 �$>Bi,�y��vQۑ�S��G3lt8fUDmɵm��?XW�o*�؀\��`�����7ỪX��T�|���Q*�S:�Ĕi�0( �k�����v�
Y��;{��W���� ��²����sV�1��T3�6�޹���»"���J*�Σ)B���d��aU����(P��\v��Δ�V����z��qI�(T ��lwRGB��ע+	8d��9�檏V/�
��w���#v*�R/`�����{��"��E�meUVJ��ۢ�� >vI�~z �"ۤ�wC9�w���_�	8:\}�x�`����6�B����;�C�p�+��|�����zr��tt'�i�ql���N�Gb�A$���43x~^Xnf]�A���B,p9�yd�3~5�-}5T�}��� ������Z!+�ӕ/h)Q5�>����m-w2���1�	z~&`�R�@&4V��©e���H�"���ȗ�w9d���v�w��4_�t��b��j�{5#Ds�)���p���J߳iL�y�8si֍;Ng��.�v�t$(�=q�2.Id&˒�}g�0uN&����.�
`�Ր��""J��v|�t
��"��Қ��9\�F-Q����z����8�2����$I��'U��lR�r3���B��m����H9�;��8��7�Y�5�ڼ��������o�����A��I��w��\5�mS��]����X��5�Aեq}��H�����q&)�
��ƈ��mN1ŀf�N��@��ڒ�#SQ����;�)��M+s��������b6��ex�}ޓ���0Γ%�g�b��:}�C0� 9Ï%��ZPp���t���/����k�ؘ>C���n�n�e�������I��,�)5YdR9P��� ��߇��Q����h��_�2������  md�������K)���-E�yvE�Q,����@��!��|�w���9�D��Ofn�/U��������77��E	�D��p7|E�����3�z*PE�Ff
��3��(����Ę�nj}�~�=�&�b�V��+Ǫ�f�Ta{���
Rd��Ny.�A!1�y����(��&�um�-_z9��y�v���Yo���_��G�(ꘅ�'�p��0�؅8`{�q/˓�%�U�(���w �JQ�߾��������߮���Jq#�,R��N�\ $����dq�{Yqr,������БM�)�������FY�#Z\��>(P�(C���?=9�+L=�9p2��ó�M����,h[�-b�o�f�lM"�-5�+.M�|<=DӘ�'�c�f{R�q���M��["�W:�������x��F�qd7*A+�(�
�ݯM�������g� ���)����ç/�ּU��i4.�O���]'9(:��R�7v����]+XT�@�7F��xN�ڇ;=�ިv��n�B6�_7�s�����j��ns�~х 7yй��k�(�O:zKj��G&��#O0���Wӓ�#<�sH]*�>Z��<��ٶ�^!0}��`���{!h�zZIȾwQ�B��*Z�%N�Qe���?C3�Rv��Ҟ���>�q�=� �D�%���̯�=i̋��B�W<�� �Jı���=�Kj��ư�r����o 32 �'�|�j�M�='>lp�D�{&���k`,�"eb�w�_`����1���ѿL��Gh�e�|T[��Z�R��j�4q�����>{*r$/�<�}m���\U�#K7��TC������d��XR��IE|�z�}�*�};�^�\���h�ً��_�������h�HW&_x?.�*���\XoY?�(��{l�a��X��X�r����lm�/|C�Z◞���`!�|�u��� qR��}���K|���Mi;��["���X`�;�# HS���J�?���)��-� ��q���F{��Ũ�>�AE䶦��j�R1�n�}�UA�3�Uu�F4��_m�H�hd�����A$Ԕt���b�w� �.�+��Ќ}��]�C�\�R�'N��eb�]��3�*V��@[ז��?�Cp;D�'�� �O6
���p2�� pk}�!�@ �ũb� qO��kƳW Өcq�1��<�H
Z�|��Wv�V٠]U�Y��)YV�ʛ˃�=��۵�c<sA���S5�� �TOQ@��AP���;L�3.��_�C���7��P[g���S����f(Ivq�0U`~�z/RDk����#�����0�,6D6]o�b\H-���+"��h}<�H}��ύX�e��u�M�����(���8�۪����l�ޛ�+
%����Ul�TylIz�^�_�Q̞žc[t��ua��`tk��J����_owL��Ԙ�
�Qǉ�#$3���W!C�ǣ�ɤ�f�E��pR��=n"�q�K��k
��������I����	'Qr�e��9�����h��ٱ���bq�=H��?=�~(������;$�������~gl�lэ4?�~�*[����`Rޛ�*��3O9_`6�T���-+����I���,�çQb�Xvw�Sx��~fճ�hm�^���dd�A~���嶒ή��!vU�Pu�UJ�j�`�n�d�������	�%,2�=Ǖ7��esn �_u^}Ù^<1�(���H�F 0�=�SPb�4��ر��9��GJs׳<�$�P�P���	W����~J+��7�!)j�$z�Uڶ��N��O�>o"�1��]OО�����W}f�� ���b7fV����0�Ȩ�q�$�\^Ֆ�My�BM4��ޔWJ��>ߓ��iQ4ָk
ă�}� K�;�
�5��GXWNm@�B(v��[���@(�h��IU{����'���h��u�Q�]��l
`�����.9f���а!Ĉ��3��9յ�Vi�Gbw�di~�B�J8�JD2|@i_��,�m{���Ν��p��5�c�ӑ>��8g~,Xo�&��<c�q>�,,]L4^��Z����j��!9�6,�m7@h�1%�d��
>D3�a�����"G��Y3��j,ï� ��8mkq�I��kC��ю�w���v�Z8j�T�@����|�X&Ay�^*`�������b-�;��ߗ;WD�0�4/���x��C%	4Մ�Z�! 8~�����!��F�bvD��bυŊ�~���J�i��J���_!�\y���0��z�1�u����3�1�B���(2cٱM�5^�H��/��x�b��k����wF�l�_�ɋ�X�W_7o�t�P�x6��E�J�a�����le���p�h�X�{D������݌���"�H,*9��v��}��P@��r��MG|�5��OɫdR���	ʚ�v 2ع����b�W�4M���@��|�74�R�Z��.n���C�y�{�B���@��5�g�JLdy�T<��z�|��9����fhYХl��Y��h�)���2ȇ	�Ksܭ�3��a���� H�aƈ}VI1�h&Tꂢ��Cĵ��9�>�;��ttF��B�;�|�<��n�\�R�A�iZ7e�R�X]R�t��{tP���
B1���Ŕ�2\_./�}.�9�	f557,9J�s��`�gMb�.h�eg��k!��б��k(u�2#��7�HQgb���Y�� DDxJ��I��oO\F�0��~7�8��u~�/���)��x�jem�`>[��3�i/_��j�箂���q�"�!� Y`�JAwv:aL=�a?�
n��D����c[Χ��޾{��8�7���:�v���h���w� ��1���n��k&/����"��gj�07�^�~�xkǲ~
l�/S���/�s@EXTH��z�fw'�R���iqW+!;�RL�<Z�	�4?��T�ʉ6�s.Еv~{��<�N�>ʓ{�J}��4Da�h���i3�r��P�N'��ͷ#]3����v�r�[��n��~4_�G�Vi&b�
�<Aq�ȇ�� f=����3DM�����f[��T[6{��i7fR ���>I��+k�|Z�k?�K�(���Bq���|�)sM��`kU,RzFv3KNrC�:���I|��6 
�gt���X��'�����ej2�ȥ��-����À��+��ӝ\�o}A�]�*�A����Jf'���ā[�12ĹT���h�-Ⱦ�/�Gf�����d��ORoV`G(�?��gz�m���`Z�C��󶫞�}�}�Ngԫ�\ǆ�W�?��$�l1�v�~c#lnw �l�yw;�q��Y��rD�=�{�&����a�����B�n����iC-D�����}V���>nl�VH����Y2A�\�`��z�[�<��ҟ`�i�Oy�z��/��iL�G=��{F��'#�6@l�$��g����HXߙ�sl��[XsI=u��܅ѝW��^�D�o�5�_{�`�m�0��x�s�l���*�O0�zgH84��=�S�������2ià�3cn+ ��N�Nl�ǹ�`�2'�*A����9�CWV�/��]P�f����s�ă|x�U�׻�~_aLa���˶�K��0�OӭN)�˻^��|2��v�#�D�M��Qo)lQ2&�{*A�mc�:���K!NH�볽���t2��s&�/-�*��ܲB�_���=1�'�Us����d�B/2r���4�Y��إ�-�{��)d�F������v��@D�u��� Q"̴�3ލ��La�~�.�:&^1��G��K ��4��cK��X�V?|�Y�p��m>�0o%��ьXE9�ԞD�W�>>Mn�6�''>��g����<D���S�-��,���v�T�"�)�ȣ�-m۲�C�'�[˱��x�xt����f����vOT �E#~a����u!5?��s�Z��[g�J'�V�ڠҀ;L�5 ����C����M,	p٣� ��y��9��\��d(�Gux .������,\�=F�����7ò�8cL�h&"��<3���d�?h��gbq1�}�u�sˌ��*ey$�#}X�X�z:���q�0��}Gdl���M��(�́f�g�A�z����Q��z)�f�,j�]���Oy��{��-��YB���łFݞ��H�F����|�k�́/�u� ���5D�y�4�D�X�l���'����l6���VbV�̀���4��N�mtwOXJ�T��M c�8t5n�m�>�xu��U mGG��F!V$`B�k�5
��8��s��ڧ��*�+��v�0 {�Y
B'Z�>e�L��.���vݢC�h���ȩӰ<�,X��AH�R�k����{�5Ƅ�tI���R���.~-���9.���c����vaR͒��&R���Zn�4��b*�Ηy���t)Ք�O�
,5��)�. v�4��E�d�\�ǕJv�p��W�9-|=�����j���+z�(�GA�H���n�9��r���s�$���"v�A'<@Q�D��tĂrz^�N�9��e�k�YB�EO� �Rv�0�����|�yx�`�A��h��w����ͬGO6��vU ���W}�8��?���.��g{A������P|hhn���X�}IL�M�A�_��D$g�t:	*`�ƹ=���Sd�ٱ<����e6�{Hw��Z�,S�ֻ�t�>w9���i��=��>j�4yc����ߒ6M\����5���]�{;"�^{w�n*�'7Lu[��U�)u¥.#�4�Ӗ߼������eϊS�v����J2An	<��]�uy����XCDؾ	j�&�~��꣞!���h�������ل,UB���c�_��W�=e����%���.g40i�,Gj4��1��@p�ą�`@].y"����{\��t���[<|
�d�s����s�w1H{��s{-���B�?L�����n��f�CY�`e�����<߇E���sz�v�`�OB!�$��g��zcE꟡U1m5���K��F]���\�a�h7�=��v���S�ە=�n����g��eVKq|�7��Z�Dl�	�,aîP�ܺFm�-��i
�`�aڌ�qG� ��7e�^�C�":�VB��ߕ���o�kqCtJ��A��A���q����W���j�C�gϓ ��L�Y���r�T	E�Zh*��/hClɁi�^6}�Ұ�#�I�~WM��ե$�)`��P�>at���4}E�����w��D�N��:ͼ^>Zb��ŕ�j\���*ެ�`�������|��:�&�^d,�~B$�-<��{�
]'6޾V�X�b3v�/�{��|�]/����!�� ���t- ܺ�{2N���M93�il@� 9��D�C����T�� ������X��Q�+ŵ�'d���a&��-�w��힂e���&�U��J�������)fʷҖlj~e9�{�<m�t{�I�H�ˉ��>�S �����\]�J��[�u�Z~���(|JDg��'{����Z��(�{�AAi�>������
��oo��A�2��J��J	XU�����r���ˍ5��n���uuCC�m�,��F�[X�6���2Ӄ@V2��}�*��ZW�Ҩ�����⨴L�ȳbi7BkAt&Kq��^Q��v��(��{��7y"��m����W��J�	������J�X����ج
J�7׀��H��x�n&>>%�� �;��������a/\�9J����@�$�nw욻��E����"�;���f�f,�pH���H�C/�_o�0G,q7�y "�vX�uI7x�������c������[VC�6)���A5���S���*�>Z��Y}��*_}|)+0UU�b�b��lz�5�x�/�i#�n�;N��kh2���n0��˨���j�[�\�>	7����j�Zá���NƖf��7<�y�����t�����Vlr�`�������j$�"i�^�j�U;�8��U���:L���f�R�S�e���"�)m����n����3�9�����9?�Y���r2T��A��^2��~�S<��S���u�l�T�v�$|�f�i���|a^��m�[H�j�'¬��90�3����՛ I�+��@�⌲�k�*3g���pI ɹ�\c`��N��+�j:�[�t��ȟ}.a�O-�D�|Si[/�Z�+��D���x�腁������KW����=�۵�VV�}s��^��nGO\OW(�|���O���2\d$�($V5�O݅�j�O����xub��$	A4}��v� g��#�{7x�{0d:?s�,�\���"u�e����"��2���E�օ��&���$�ַ��נ���f6Z�ClF�ۙ|��tˠ�J��B����_��1�3+�^*�F�W����V��C�d��{~��.���+�,q},�;���������ٱ���	Ǉv&ڏ���J;5^ ��z�l�p�SXX�&˼-)��j��j�K5��./^a[�y��3�ݎ����o}��-F��t'��l.�>!B��GЧ�e��h�-���	�b�H6p-Lϗ���1o1�oM��w�N������u�Iކ|G/D��2�SLg��.�v��D!L��˪��[�p�>�P���<.�	64�<��)Fเ�����Y���@;}���-	�@���sF�Db@�j$�PJ��ǃtRy3�M���e��g�2�J�L��Q�r�6D���Aw�{Q�Z�{3���ǜ�%ݟ�<-P��ɩT�71�b	�q�y��	���!�_*NY�H{��֛܌lX�9�+�.�����'t>�>]�j��~��kRKU?�ۆ�m2�� H/���_c9�cP���z��k0�)ç�N�X�Ϧ�m L�\w=�ӳ4�^�$E0����N����6�LR��*��6���� *�aU� ���FO��)�9I���g�5���g�:�xEݳKcMgoҞ�a3W�|�g���b����X����;`Y�� ��kן%1a0����= �HRUS7�r���G>�� � [���캼e2��;Ff�v|��"�YѐW���q(���S(~>�x��Y�5��ֻ�b�7�i���<�;���G'�k�I?�yW����'��(̖o�B���no}���� tb�B��y�"��ʠE�9�2R�s��� �'�ku����eD_Ge��}��"���6O�a����cy9���<p	�7L8��[��2�;���	;�~�����R �����xp�q��$�$��ӯ�s�O�?+���m���/�D���� K�W�4��䦲��M6�|�H�6�θOS0^��sڌ�����������G�3��^fs��,K����q�iT�����j%���h��̮�쿜��@��ǈ�b=������-o�������d�刕�a�/{���/x��tI�_C_J%L��GŐC�t���/)1䣋{��{���}�1\���n)��p�� qm������m,څ�3��u(B��p�zf78�r��&�m��pl]O��L�'���u^)���;��"|��K�P\�͕'I����������'g)$���n�@)�#8O�m��6��=�ʅ�X�`��[�;XR� 'P� N�	����1����'�b6Yt����Q�\ܱ������%�H��#��Y�8�z6�R�Ƅ$dD�xx������D"��^d�33Bp��2p*����������)�s�����bXjNum�$l������q7_�c?���<>�[��/j��Tm�$e�W�DqH����j�'�`Ec�� ����wa'
��e}�iz)���E>-�@7$c�c��̎�ɒ�P�7�Q�à�}d��	q[�e�RK�UX��܅��3��}���#M����ā���?)�������]B��VQ(�u��j���`�ʲ@�$�]�}���98�� ;�������/�Vl��(#*ǊJI>�H`�����TӬ�X蠤����MZ�3�I�(ľf���o(rS�|��B4�B����e���O���دt���a.�1�<f�jXzSv�����<#=�=MMrw���t��z����&T�"��n�|nE�����Q���B��H�2 &��{���@��CEpG���'*��T�����D�e�F�O*�L�9�_�_tΟ �^�ź��[{�۬y��L�+7����r�����7�'����p�����cZ��j�1��Z���DG�(N_~�d���Ξ��f�d9��1���iX�53��4F]�Ļ.�u:MJ��-8 ��0�B\�s��Ӓ���K�u;�`%��*�5q�}e]��
�з}O�I&����`N�~��V�Wb��N�h((����{|��/�G;ٕ�������3�H���8o�S��6�?5Bq���;�P�����M�b��ܶ���L�=P���B���	���1xw�K��L[A9�ɀ$�;Ri�uҀs����1��xb;��ЪN�̵d����n/sn��|�&P�u�*�IeӅ��̣�(ƱE�O�%;�;��E�Pв�דִ��d�/���+�a��X�l'�wGj@	LKO�Д0�u3Cޡ�%d���}4��d�}sRW(���A룿]� *^%�紐�,2����.�@G�И p��8#��Ռq���Jr�t��z����@0YnV����X�g�]���M�FK�',�t�9JC�(E&8-�@v�׉��G�s`s������*ŴU�2P��gh�����qv�F�pj��y�g��
hS7�.���|yj��Nk�`��X��5�`\�ʀ=�ӥV
Tz�v�K��	X�9H����fxY����������Pu�<���9��L�W%z(�{�e�W��J�Cp'u��X*]���A�0.��/.�iS,	̞*�!ۗ]j�Ix�1.MTK����o0�Hl(�w�2�B��Bghg73�� �!� �8Nq� �)
�Oi	Ə�+3S���[b�ęM����zsx#���ǰ^�2���ez�����Ȩx2�)7M푵�A���dY�C�̠�h�b@s���']�P �r1-��=�J�#v�0~�=
��+ˡ_@�4J���]S�Ɵ�b#ʝ��!	�h�{��
�g<��7�H���[���x��|�R�mpș�*핗��ɣ$� �s:d>�oNM��Z�+F�ٲ���՚]�W�?|ބ[�n���zkZ��w?���\����vE�Z��M�M�L�,�R4�C��\�|�a�ky�)fG�� z2�,ڕf��d�ZR͟)�ɳ~�5���D5~�D
E�B�}8� f)�ۋ!����E��(k���kJ;��<����l�?nx��K�`��.��`�ʻ8���zԇ&�`�qd0_�>F�̕��lʂ.ME��<�$��>��}r�Iܥ͝�W�¢�Q�;��t����F�>����½u�:N��}�e�w_��WHcx�r�i���Kgc��G�[���"����]<M�%l�}��F��l���5l�g���N:;UIH�����eO�͏�4C(��5������}"��r����o�I�}e����UX����T��D����h˰�\H����*�_�"��)JH��S�|}� ���̋fc��r�m@��7/���o86�fm�Bh� �\ѱ��l��{�����-�5�.%j瓣���otF�+#���������u!��U���h��6�����[�}~��S��X;������M#�������&Yfl.A�@d�9I��N�����ݢ/�P�������0�1��ԍ;�Dc�cn�V�&����Lڍ�S3�-���|�r���!��zlZ ��<��n���/����o����j��f|�L0������'Ʀ���0���3����e���2��3�?܂�l`zg}�F}��qB\�7�Y�΋f邍�,L��j��p �<Ct�ξ�l\cЊ�9�EhףG���(���F�M����YD�G�/'z�"L���tfO3X�6�+q-�O��9Ų��EK>�f�nE���lxB�,�{p6?$T]�2��FVn�t����N�j(/M>��DDz�̿��ۡх]����"L�$�B��<5�9{�1Ip�����NrIU
wo��Fr�p?!g	�,
���6y�X{+��!�m��k�ԇL��ެƾ����5P����7����X��xp���/N�q�8����Ϗ	�`8�&�g� �a���u*�.��rF���^ �Z�8��n�����M�AVջ7>�;z2i��j����:H��|BA�3�GyN��5Q}`P��m�4��:�������(�>�w|Vu��+����q��`������Z�����u5>�_i����K e�ه��`ZK��0+ ��m��́�(���ɋ�{$o@��!�E ��hCA|={�+*V?_�}穥X���B7K+��Z�8��
����K�|Q~~�瀀[&�z��#j�����ʟ��:��\�q�ڈ{HsvP�},��[�@��b�^�k,�+sl�2��0��Q�����i{�`���]o���V��B�/�22�����kc����s4����-����Dҍ�����O��I�5��-�t[�Vǿ�eW!�7T�p�;lD���_����k�u���~���v�#>�]�x`�V�l,¿��ۉ'J��������T�]$�>D��J��UJH�껁����KhӨ�V��ɉR����8�8{˽�����EGC���R@��fs
��l8���\�״�2��.0���׋���]'�4��
�S!o
8�g�d�ShuPZY�1t��Pa���F }d3�9�Is /��d���B�w�Z�T�~�^nV׎Ac�8�Zh��<__�Y������:[7�A�Bx��*���`��އ���r�n�'����&衂�vu)u��o��t����������a�J�G��=bV�S>�ϗ�(g9��Ǒj�-���!�S�C�����HKP����C�,Y���M$����{3�	��&1�sP������`ޱ��b�+�v��%%�jL컦��P��Oć�qS\\!�E��u��1 ��ICx7K����<��Ƽ=䟾i�;^�v8]WU`�Szp�כ؈/j�� x�߃���a ����\`f.L��|�|,�'�~�K�_�ע�f.,���b������!�SF�R�BU����a11�[,�+����A�����8)n���o�wʮ��>����X���-�m�E�\o��ECF��<�R�GW��i��@����{��l��~*�-OG�z�]RWHd0���.ЌJwɄ��p:�'̕갌Y���n<�
���oW�c� G��y/��O;���!�DGd̤a��X^�~�J��S�����:x�M���B\�W� q��B�3�9�P�B
��{f+�YW��BPh������s/��]�M1C�Ï㮨6���"4��Z~uo��WݎC�$�$n��m�H&� 4?e�u���Sfq(��02%�fP�A`�͑��=�1(f�Yy>�p�ޜ(��� d�x�&�=0	l^r�j�ޮ7M��03~6gG }�3.p�Y���?�L�,�¬��|��
k���/��Uϱ��Pg��F��x|h˭��![�#����D���p3��9`}i��O��0C�M��g0X�R�s�����!Ta�&\O��.��پ��Y�k�0�uO.)6�:@Q��H��M�(�fZ�������AԦh��<��O(�(N�s�2+��^�Qt��E���������}0l�6QJ���@���-!�F�_�h��f�)i��ڴ0。Wq�̬e�D�����m��^놁�|m��`W.�%y�1��Ts�9+2�$1g�X�X��An���{�Y����W}��4�?�c���\"�؁���0�Q.���˧�"���z��D��DaJ-����&�����2&Է�@�(���15HY�����{��m����/`�$M�SG/Tl,Q{��ƾ�T'��?	d2��$eHi?�)�	�7֋�蔘Nqt3��T�pK3�[V�)il�>�칓�Eibc)����s�vm�M̪F]��+�+j�Π�|�t�����fSk��Â�������y�E�!m�T\
YC��mx�3L�m7�T	V�R��f� Μ$�b6��8Tu��ٽ�0�߷�B��*��4���j}4׈G�N]wW�eޭ�ʶ�p��烕�y<ǩ��U�;/�Y�#DB�~�z,ko����ҋx}��?!&C�+����
�R���;k��X/�*�t�8�AQ�wv�G��XM�{��A��by�k�3���.5��
�M�������?�J��SnP�4����E�w'��*����^���k�	������5��O�,YĒ�bT�H	�v��AsOTȫ����5T��F�I�����&a�����͂h%ɮ�I�"BW���N�=%~������ko�)`�U�9�˛�gl��]ʇtj��*�nt7G� 1c����V����%Z�WӿN%��x��I���?�H��tP��˔_����}�؁�+�k��K&J����k�`�x��>����'@��������[/R������5w��4��LO%��V����i U�C�z= �Z��gf#�ri.ޓ�WϟÔn��C������t�*,������P�fq�>}����KWȻ:K%B6��7+����2τv�RM�	�E���F�q�� ��h �JC�A*u�,S��'ԯ�������	�a��6��L���.��H�� @܃�$rMj�DA(�F�!o)�rB<�;�Ԥ3[��*X��7nl֟^�8�'_�F7>���Z�y���Y7�ደ/�o_��o��j���MW���B�:�����g����4o>�Prc��F��p[�e0��=~:N��v��U(�'��o��,���-D�6��=��M�t�P���ɥ�vaVWzKN�WG��=�q�Z������٫N�y��N�	vn��{��ôe�ӎZ�3�c�Bλ�6Tb�A�;�\�b�)	�X�Z�Q���Ρi��!��⪳n�+�W�hd0�g"���Iw��w;��`���Q��&����\���6 �A��a�3�iG�������2R!�����^�p^x~��7�cQ���z��<�ߺO��;�O�8�D �E����>y�B�@o��|	ֆ�.��q������,} ����V��/��GZ���ҟ�qf�R�G�O����jN��	m�&��ߢ���n���	)��y����U�MNx\aw;A��B��yU�����-2�3pv��|<an��dhE�6!�f(�fP?�^P(�v��k
��	��B�8	���*ܞ������9`b ���C�P�2��?4>�GD�U�!w��L;sڬR��ً��S���\T������`�X���{ǰy$-,񸖙v�4�yG�ԇ��
"�B(ɩ��|_�������a�^����6H�y,N#Q��3��29�Co�@�2P1
{�*�\QC�d���87��S�P�t�額�<�R�?�R7~�2�?���� �"!�9�&҂�a�lIn4d	��˜N�1��P��x<`��A��uC��� �O8��ylι�3��G��4��L�VB/G���sp�D4-�B�L����Y�$���A,���QIk`�x�J�c,;�Ua��;"U��g�j�OsQ��t��`�?����FSFG�刁��Dھ���tx�3�ރ]*KZS���tb�x���x�����ʯi$�U'AP�Sº�⥻�3�p���,�a����iYO<4��Qj��\.�<Hp�������Y�`Kj�}ܡ�f�V�R ���S���8�$��,ys���]��]FP! ��F٣ʐ�f�c�� ���1��t��`MxM��C�_��,�����������A��բ���_s��E��&k�UכO���*N�Pg"P��Z�=҃�H��ʺ��ti{ѡ3(d�Q���v,,ǥ�?�7��!q��Ă��Ww�