��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�8k�)9�k���J�f ۘEN�R��>�Ug:�&�1�|+|��%ٲ���,㑍��kN��`Q2ퟩ��C-,�-��]��{i�Qs�ɻ��"ڀ��vcӪT[_��N���,SƛR	�'F �<�GǱ �d�1JD�·nu��K-:Sl��ŀC�s���Z���g,�r�W���J�m!�ʻ�9��f�د-�����U����R��IFϭ^Cc�x�_��3:a޴1S�>��F4�$�W�:d��Gj�K��n�;p�MB�Srp'�}�����YQhX1�E��>W����/�.�>^�JM.(<����2�:���4�o����g���Ϳ_[���h�7���PHi�������ǌ�] �T�,l�_�S��	���N����Q~���������~��w���3����О<n�K����CD��+V��%�]���<��C�c�Q�Ma�O��
�Va�k�{�&P5��^�����vƄ�>-��w`Y��0ó(��3k5J�����A�������L��<��m�S�p�$�v!)����R㿃�k���w���[>�uZ�/4y�Ѳ	p7���c�喝5﯁ T�T���
Z�
��9�NA\��sM��f�<ft�B�׋��#���;eB��g�K�؉U��2���Tʼ�~�-ٮ)���b__� 七�䤠��ԅ���Dj�B:���<�V��-�W9��wa�8��Dfٜ��B|;Go(����@S@���-|+V���kϑ�4�e%V�f�{a�2N�S{ώ.��p���W�A�x��w����*����o;r������q+�x����=����;Ճ+�`�r�<�#តȡ?[���j����U��!�P#P�g�������T��6�Q'�0�����7c��|�n��y98�+�����q2��l��@�v">�I�A�˦��{ƒ2�jX�77Fw99��"�-�' r�쾷Z��+�UQ'���hUe�_�k�.(�ta����A�E��f�F�:��
��P��t���g��3F�mQX��x0�Pߒq
^H��[vu�����	Ky�\h7����2��������
�w��T��/)����J����1G�Ūk�� �Lkh@�z����ӌ���-v�ϻL�!�[$���P��/�I�P7�(���z�|ry��o=�/-��,����c�c���w��b�sc�$x0dx�I������]�~d�/�/�<x#5�Ub��Y�Sߺ���ޛzc&�ׄo��/�ڶ�U����)>~��P�*�\�O���@��H�)���^�-����Φe�b�g�?Mӷ}�=24��N5�ͣ�Za�n(ID��z^g�	��IP�7Z�{�z�����R�π�i6���[Yc�	�`�C�m����X`G�pm0m����w�g����,��؍�3w�Vy��քo�2n���$�^�c����72��P�|fN�N4~��gr� ���Z����,9�n��?�Hi��	6.�i��"�z||�
\�X���xF�\�\�St���k8B��C>I�7ّ�S���n
 <4��f�P��R7,8�V�c�b'�LK]�]��� ��Ao�1K�Җ��3�X��k�z� 5��1a�w�*'X���B�X25@�d[���5��^�}����H�X$���ӊ�������8��#�C^���X�Ӧ�7�P�˞'	�z;��U�\�3E<4�k'�^:[W�m�s���'��E=�E{9�S�U #pZ�S6ja��b�PW#s4/�Cc�CJ�o6�R?�ӭ�q�6�������h'��;�Se���=<��"�v���K\��c�.ǍH�aK*�^j��9�C�%G�'PH˶�Zt��=�C��g}k�CN?t��jo��]g�p,$̣p9aGJ�	�e"�A�4FI
�c�u:6���Z\)D��b�T����<��tm���ԈJ�J��c���q��y���m7to7M����7�lɀ��n<�j�^<�T��0R��W8��P�ͦ�&�
|����� ��I�$ؼ�>
-�.TA8�t��됾` �ۇx{��8��.0*�k�u|�J�ȡ�����3zܢ�R����wWr��S��k,��z��q[($����@����{D�WNp��ut�Ւ���� R'(���ͮ���Q�k��d[&_�E�A�����W�H'/�Y'��I����H�$��u�s9��5��ԡ�)��m�� ��N ,H��Oxa�1NV��0���x��K�2mv�5rXg����-+QsHXfю� (Ȍ-��6�RS�_�a�+%���Otaŧ}F�&|-�RNh�5�ͽZ���C�r�"2���=�	�*��G�t?<mV��H��������]K�b��ן��$�B8\=�`��}ԼPLdIE�h��`G�7D����"nE��z�x=��=�t�F���?ƶ��!#6/4pnE㺩��0]?�d�g`SG?"O� �}�4�`�c���w.��ׅ�x�fw�F#���{�߉vO���P�:�/���b���\/ȿ��%�2j"5���1\�b�����>���GM���~���}���/r{�G�e۱�$+��� Z��$c�u]�H+4���f�#0���ۑe�z1\���t����>{{��"����[�5	��PBω*ԝ�R�޺g���MHΧ�_e=<�p��J�P��g��'^&;�� �Й���cQM�����&��0%�%��&����Oۃ���J۫��k7A���N����tM3&2B�(}*��ꀴ��g4���TʨMs���ʢ�3����3�q@�ч��O@]�� >5F;q�nNS�9D@��G�r�zO����k{ V�Nd�QZ�)�=skѢ���M�F1緗��?/)���0r�-T�3�W�I��Ï��\2*[��D�G������(A�pvŮ8��VӼԵ%._��wG��x���Xm�J��#����>�Y^^)�^��M�(X�#����o�����p�=���/�ѓI�CU�0y�T88��=�N��Hm��9h���$ �S��#WB�'P����&�U��؀�0��h�p�T��퍛g����t	��3�`V~��F(�O����f����_�&�����&WАݴ�W���S}��b[��^��>��|uϭ�)�����$+O��B���(��Gfd�I&lQk�Xg<��K�u�D�b����0��� �?[}�����_�!��w��?� <I�KU�R���
c-�9��0D�i�������rl)�^�xJ�G��"��E�Q�W����I'����C"�{s��ZC�T�?�m&�l{��P���n�[6EAlN;�۞�|"7*����YY�� /.ňg"�vj���¥N�µ"=Є_?~���q׀	��������.%�L�+i�oɰP���/H�du`�ӯL�Xz�Q�ޜm1���7^�A��BM	�ɐP��oW�,�|�EH�Fu2�8= �L��>��܉�ގf=og�������#���U���S�Ń uz���J>�R^Uq�>3���K�Pk��h��;�Xj ���b�-��baNhi��B3[��Fb������\����J��O!
�E�=U���~��ؙ5@�A,���<�=����W5�KF��2��� 淓���^��� �|����0�D^���ި/�b��U���}��+�V�]p7���r�_J%\X"'w)����[R;¨�WM�]M�lm�X;��Վ�n�͌�-��Ei�0+⟉O߯��0��s=(t��+�)�-�L3���ֳ.0�եQ&!�";�c���؅����ls��EZ����7p����{�j88�/�q�y�]ߡR��{,&�����̩�����vJ&�܁7qv.]�R?�NLo�ָm//�z�ާJxD���k����D�}��Gs�� ko�r4JS�a0:�h���aG˨��OFzݸ�b�h��w���_,�f��~�yF.�h���I�)�1���Y�=Pw�{�Yu��` �R�/w�#�����.����`"�=��|E�4Z���ݶ�[i�y�ɺn�w�k�N��\�ϘV�N�L����QD%ފ�w4TO>�+�I'۾ &
�09Ck��s��EЩ�]u�����bU�0�)i,�b'�=.ל| ׁC0}h��'g�%�:P�z����ҁ���� �����93��`�ߛ�� �%��+�T�F������07_21^�K3��/}�.'鯧�s |0��R��8P���N�78N��(��:�?��tq8X�>�nC���d:�2E��=li��&(��,(�©/�Ñĳ���(뜭�;����X�[�M�G�s^�h�ߧ0����h,$��v�@���s��M�,�y��2xt��7�`ln�d���*����r�Pgi�|��j�^�?+���:��L�b�jы�LJ�"Ԓoh�zO��SW@俈F �	�T��"�jJ��\U��.Jc<��,=� �B��^��k n��&@����D6�����m�"�����(
�n�K�[_�ߞ�c�L�6��3pv�4gՊ�2{��ZAk	b�W�xL&�f��qM�u���yplh��u�"�������Ё�ZlC�2)���.�0#��4��s�B�R�>��c>-Z`V�b�J�i|�Hw�|���h�������I5-�G�$���
x��9�"=�f�?E�@ �d7擋�<F�7��T.��q��优����Fx�g��av��F[�Ѷ���)��q.#[$��B1�Q,V�zN�x@��azڊcS'�d�<\���n�|�*E��ը�w���&�`����c|7\�0U!� ��v�����*��-h��O���H�Zi��M�����D�+u
���_�"�H\�x�ZfƉ�e��Y�Zc���A4B����$� �� �Ⱦ%a�ў�9�;�d�|H��=�4�� �J�v���!x�`R� �;g3����ˑ`d�X�B���&�8飮W̳:�ĵR&�r�!iΗ��oX�`	0FJ�'�Y���U1�?�V3��H�wm�ҵ92�jR^�È�B{��gL�Yb�|*�~���$.��Ӷd1��/YbdˏY��
5_h;���K�Ix��O�z�E#�1���czR5)�y�\1(x!���f�_��ݷ7�'�d�s�-XT)�VZc�W�qľm9����S�!��V�*�����v;�$�IUN�=&H��8�,\]R�L�)۹�L��e��N�������c<��������F}�r�ZJ�����;{ǐ�}������2�j��A��dDD�������(W�W���r�y��<��U����Q�����9�YS@��ש��뽢c�9㔻X�o�1��y�2A��k�q�<����`����#a��k�����lH�K��n�*l�w貒v<4d`^�]+�����͌�ďOVq�?srF5�pq�\�pzW�Φ3>o���g�'�ZbR;�["ߦf-�F:S��Țѐ��A'��[p1��g�Ў<�	��N2���T�Q����zF��. �N͋�Z�I�$���=�k��`�y�wcP΢������Ҏl��PT���'�Rl*�w�:y����us΀p�;7#�ԯ��a�6	�T%�+[3~3��4;˷8�=>���/JF�%i�]1�۬L���J&J�vSm���?}>��V��ʨ�f
�/k�=�;Q��鳽B!�i�%Ԧ�Y�9Gj�>l^j�k��o���;��!s����r�� ���Wsh;1��j��q4��55"� 1A ൏�o�E#F`Ua�J�ЁqV�E�ϰ8��
������ߑ�A���nO�FI{���	� 
��=A���f=kӨ4?� -ʏҎ�<�1��&�-����46Q�҅(�O����Ԃ�%�F��e��X܁���|h[
$K�s�]��3{+��r���9�,��S+��Vˠ���L�� *����h�Z�6�
V.���r���h*�W�ɸY*�k�tE�+�J���)׉��PK����
i}����)�N�� ;De��k��@��YT/�M�8���v2�p�������y;�}R�&�CȨ�O�)����˛vpS�@��V�:��67F6
=�\yc���Q0�޸2�p�kxm�v�ОC�T�e��W���q�/%�q{o[2�4��T��{c���]�AK��e��\��K��l��, �Q��07������E��Z:=�	�+�6K1��A4P��������5r�CJb�b�H��H�<Kp��%���cofٍ��\,"��t�N�~���G(�q�s>���P�߁%�F�p�p!�a��s�O�'���E�%�]{��RۼI*�Rˏ&��tѺ�F�	�fsȱ�Y�#u��Z�T[�3�2�f�����s�����ɿ��P�Wh^{�ĆMv{1d��W�A�G �FH��ե=�A��W@��k_�K���6m�Lai�������:���{�v'en�Z�/�(�@>2�827��8£A��)w�7�Oܶ�x��h���@ͫo���z1'G��A�vJ��!�ѕb�V�&W��WU�z�`��@�$��X�!��m\-�y�'��?�`#�һ�8�F��(������1�Q�DN��h�"��N�\�J^1����0��*xR�:�Qb���%yW�W��&v�g{�H� >���j$�o�af�[��DҞ�a��a��E�����q����P��纆0��o[��%��Բ�!p�ɸ�%Ɵ��*��Lr�ز)��P��i`$�H)��RT$=2�w�O�2�?+��}nJ$�4,��\�.ƹ���ބJ��p�e�vg�A�q��:>z��£�����3\F�X;Q ���v��IpP�	�Q40�n),'����\ �P�.�̜JyEM~}�ə7��kj�O��A��g;��m|��Ii�H ���W��,�k��iX��l���,�.p�~�V:�"�KuE`h|f<c�ᢣ|�n�}�$z�~!N�=ڄ�����s���W�Ra�^ܤ�##e+-4i<�`�$� -'휝/U4dW&��g{�X�����Wgy��/6��'�����:O�=�~�U-��*a����*��C�:Qpb�$8FT��W�Ҁޫ�02��b�	L�7�`<f��������QC���daS+]x���!�_���ՋՂ0G���	J'vd��@��-���U,�CnTq�M�2O*�x��x=�,��Ab$�{�e�����T�����*�
o�Gy(�N2#�ϱ����?]�h^���LW\���-SN�݂�91gu�S+�/>�d�=��;ՠ����Ѽ�Xs߉���u"N�R7�SJ�:|kW� �}������F��q+r��c�yX�vp�UA���aG2G%��q��#��E�2�����3a�d�ǂl�7�����Y���F���w�eAB�zi�� ��_��	*)]5�W���u�h�Q'� b�77S����N������猭j�l�S����7���IN��!�8�Qd X[QC�h]�������{���%-���S$�����\A�#���<!8"5�H}�'��[���<$��^��k�H��3
���Ra�w�є�����w=��N`�8��Q*�/w�%��Q��f�Vo�U)��.��ͅ;%��1�ՠ�96�m��:��e��8���-Goj()�^��c�f}H&&�jF�5:,V*��<b��p� ��M��M���J[W`T_�+O~wU.v>��7�@�o��_���ױv~��Z��7i�(�y�U������gB�A$b4��&2߳�0����[#(������(��R�E�b#���� !ȶ���M�{'�ӁA?1� kyL�Z��O�'p^A�4�=������p�1�(��v�?����~���XO��1!6�Vj��X��"�y���ey����K�ն�'�dòs��]����6�i�,n�g����#�e�%w��ø1T��rѲ�R�S���l�]��y�̴L7����Q���
�S<l�IZ�S]&������5���0�ƆߦUQ�e��+�����9�Ɲ��02Edew�5��c��Q#j!MǙ��F{J[��o�7\�V�{fN�[f�aՒx�eH���-I��K�Q����٬F�x�RL w$����N�b%!#2a��o���h�
B�ч�H�������c�~��S�O@�nL�&~m�R0H0]�_�r0?˰x��u>��-���H~ub��/e���r���&%�1�C���\�6��O�٧���IUX�$�Cѽ�ձi��*u9���:�*��җ��!�gl�F�3(� ����i�A,O٢�����w�
Fie��j�C�:/+s��Y{��\��ph-�/W��;�a��Ĳ�UI��ô�&g𬠽b�e��Ͳ�蛐�	��z��k�ۙ��{sa�䍙῾�V񮹸*�o���E��N��O�2����I�k`az�.b	������,��Y�Q����ǾSi�S�+��N���8$�2�XL>�=����c������Z�u��L��0E`�~�_�D��;���~���FʉZo�BԳ��N�k��{������z�Wʔ�j��[��!cY�����S�mU%WJof4
��`-���62s�h���n�q���n���ţ�KBT���z���ܡjt��KR���(��c�/�������$��'�ժ�!�D����t�]���Ei���J�R�L�ka�
 �F�}�g1�Eㄞ/�,+qpv�;� yU��"��_# �\&Sԃ�u�4�?״}��qڞ������o���x�#��.b�Ҳ�\��@P2��b�!�����pj���x�ߩq�>���쩱h�E�'�|VQ��~m��QBJ�׋J���Q����+�Ⱥ	�D���A����+O?��/�!@Qs�̯fJ��[����\[�N�����4{p���@7��g�,W)�v�����p�v�ox)1U[Eu��Lsǫ���EA9Q�O-KR-�� W�Jf����?*��W�>�T������f�_=/>`P��	����G�7O��p�8-igRf���UH�S�`ԱП��=�Q��ν�x\^�'�8ʱX}1V�<h����YXeH%˧�Zh�R�9��������D݀�x^�Q�y��/.�K����K�H�#���W�	p��v�@v�DSZō����C{L�b���@�лT$q�H��dZf�2bE�k�N�K��`c���
@DQNjf�:4�7�O��ɜ���������oE��� �����'�S�SRz�W�m%��x�l������+�x�%���P�>�i�y�eM�Vrm} mԠ�L�&$������Z��`�Oa��J9��&��cX�5�J|a�uZV�o�^챿B's.]>{�%Z��R%Ӽ����G���{���4���~�',�m��#�0cߥY�~�宲n=������#H�)�m�ϻ�q��M�>��������v��C5�
����V��?c�s���j����s�k��Go��,�Aֶ�n�xx�<yQ�s�U�S�����@@�#/��$&��;��<����<�	
��?��'��l�,�I|��Y����V˒(iU�*3m�GQ�x�	Is�����R��Y	�}e�?����'�1���rآ����_E8�+\�yŐ�k$�:��81`��=���K%�#��8��\���Ǝ�.q��0�h�7�����r��]'�u�M�K���s�iVze���.�~��!�XT}�0��k- �5�F��Ve�.¥eb��{p؊�54/��oW,'5�E��q���)� �2z��R�`gL�S��67v�o�L��|�(���#�Lo�	�7M��gksyh��xUg�PN�>҄����C0PZ$h�J_����R�#<+K��^��ei��Ir7�R5C(}n
3����De���s�<�3���|ykV0���ZO��P��r��G�P�_�@{�o?龕���v*�#%*݋}uK�`,i:2z����$7���FJF�v0���JG?hj��{ɝ��=��{��tו����(�v�9�e �u�s=��ͭ<�Ĺ�1�&�Ya!�X����mL0�c��E���QQ��˓)f�L3�������6��3ܓ�;����}�_���� 	
y��-�?����$?�Q*`mYS~w���d?�K-��	-DN�� h-7<�	掑���L�R�}��q���Z2���`o����<*�lLH������]��3��*�I��ך�苦���.*`Y���t�.t��rf���<�4�s��hK`�!�^��R\���.%d�n�5����w�,��U�Bi����]@X�t��n� oX8s��|�hZ�5+��)~���������@9N�!�X?���;��J�(��ŧ-9Yׂd���������OP���I&$	IFp��>����{Sk��Ӯ ��k�4�B�Zn���������X���
�@_:�MG�a��L��}cV���ۋ�qk4����_��/_֏��IP�#A(���1��E�'�2<Ƅ �u ��N^)J�ͼjjj�Uvcy�G�j���{�b?r�>�d�O,쮇��	�c�)����$�2\sm��^٘�g��I�N�ۥRE���!��I�1A�ݕ�J&���
�!3/IR��+{��������I���h�dk/�Jw �ﮮ�kC�F	Q��n�bR^��� �L��TW��f=}$,ޖ4p<y�,��zB�}R�]Q{�;��j������1�섑&*Iy�~�>�C)�.�`�9�q�}#}Lk�ﯴ���U���/V,R2�4߷���H�|2%1Xm��T.XK�l��?잔i�����f�z�Ň�ȑ�R#�����g���c�Xƀ��Fxgo�����6�q�նJ�@֙���GU�s�y�X�;
�}�'���A�$�Us�jZD�.�?��nC�H=l���k+�jǢr�$��Ըi��Ӗ�%c5��b0Ci(�k�>���UTj�C/���ypi�h���)��zche�k��:�`T�j
�K�?����sw��k|�3������K������j���ō�Hzn��{��qJT��`s�r|s�1M�T�i�V[���xm��WVo�v��<��������j�}��lI�b�G5��j�,w�9��f<KG���1�_a�CFb�&.C�Ȕ~�ެ�i�M��$��3��<z5b0jy;jpo��Oа(MI֚����u*E�%��5���u%����K���� B.8�M�h ��|Ǩ�~c�~�AA���Zr�$�2k&�h%�x��8�&4����@����%��:�_*�P�B���\H�KH�D���eh�<�)^jey��]u텥��ҤGМ�E*{�2H�!����M�\����*/�n�%�h�#T���Ʃ2$����"�"xf�p����h���_�e�9�X.��1�a�uq�n��R˹�kW��k1/w����k67���Z�4� �u����6���oD���w�f�U}�W��U�P�+k�ܢ�uvbyF��F�-T�#�����Δr�t������������Ϡ��ꖳ(?r�lv�ɕ̽=P�K��w�#Y��zXS"qu��=��՛��:w��8g���甦��!�P��x#��}�P%m� '��<���x���6OM�Z�#-�iQ?�M�����"��T����8���ݑ��w-�f�K��-��ǐ�n���
%ZL���D�[�~֎+&���[�a�lu�J^2gl>G�aq��5;��P=�h̎���P�����\�>�}��?=d/��m��f����
�Z��4��.Hw��e+�I󔵜�m̤/>�wXb�ԫ	Ґ������'�^ar�D[��\�=�4�����-�Ms{��q��3Ҥ����%Z�9}�X'�j.��݁a޾��F*�E�wC�x1+lpv�n�.�n_�.�������6	{��)]:O�CG�/>��2<���kKh�م0������c�[�#���d5��C�c��z�L��lf���&�Tz�9���r�I	��%�)|Fw6��i�[��3H�>��;Br�m;�֠#O��`���@+�Td�[t1w�e�f�XH$s��P�n�Z�����+������qc�&ϖYr>E��o������x��V���?�+pZC�i@���U=� �+x�������x�x�|����}�#M��N��ы~��a}838SjM++�܄@�S��Z�U����q��\U"0�m��5z���EuЦ���_�q}[�Y�gh֐�R��u���������,x�l,�:�o��������D�c�C���%��5^,��M��<��1ЂE�k���?�rڻ��j��=�O��~FRQbh�hբ�
@�h�Ӵm�]1Y��<:��hl��`,N����S��;��Z��VŃ�ñ#�����6 *Y���=#^��f�mX��O6�
5ot��<Qr4���Z�f�gg��l����IT�@%-�$�GGF{�J^�<� �yG̗��b44fI�=�Ǒ���q_�ؾ���Uw>*�>h��g���$�&w��^���0`�{�jxPȲ��$�뎕H�ˮ��32�-~�ŭ4���s���-tu~3ڀH���(s�������qB�7�形����"/����&���:�rU6	x���Ň���<X�����?e���E��<�-�W�L�oFZ��ةY֗j��晧�,ۿ���6����̏�ʌ�z��v��q��(w�Si�C�2�'2����!3�'S7% j_��?�M�@�e/z�����^j��i��rtd���8��R�c.���#��r��Z躷kz�7����FߑO�r��4��6Q�i�By�9P=|O-��+v�h����O��Nf����)�	�s!���S�m��}m��2ǥw#����b߼m��\�m�*�$az���$�5���A�#I��q�SОZ��,FI+G#A�ٟ��Ѕ����o����JDM!K�@a�G�0+����\�H���A�y.9C�ON��G1<�[y�F5���Y����:���/#�䲼��{�d�W��Ĺc�%Yn
�5��	.�P�P�y��O���v}z*��ٸb͆�X��z�(q\�\��1W�8������)�H�d�mh㱁��g'�ӛ��K��7o�5�,>̠�)�x��;�e�lW�U���.M=-�S��#��>{�El�͠F_���]s��w�&"9�c.�\gI�}�~����݂-?��v�g·����g�5T�]�5V�b�t���BN�-�������Mahz0^��A�5��fÔ�s��D��a���Z22"�k�2~U����-RNR��� ~>�xÅXrFk1s\�lf+t������_����Vr�΀�E��>�	p ʲ;�Ǫ1�Λ2�+�)k��G]�C�g��}��-�b�Q����h��`��\��
3�/픀��ͧ��k����.D�ɟf��x�r0[F���U�Ox����[�x�1޸�b�O����a' W\1�����Ȓ�%f�H�wSn�9P��\�e��҈�2�2�����^��ä�������x;�	���aM�(��K�ح�{�.�,����'h��[ ��p��Z���᪔�]�ҷ�\Ph_�{����xX�������^���U�[=�2�9���P��9�}�Zw;\�*~%ܹ<����VE=\�sI�L<���/���B�~��D��J�Bb�Ͷ�{H�li$uD�F�J
�64VyJ�-QӇL�+EB�@3�}����wZo,����w,oY���x�c��l������G�G8���(�.�}s�B�y,�c��o_:ݧ��"��Ur�U�>Z��$��Ģ�C��EZ�E��,�����	&�_�3���2y�{���R� �_��m88j���i4hʺ'�S�!���(���Ј+Q�̨�)��FG�����Ǽ�ћs��{=)���1��\�t1��J#�O֛�E
��,�0#<��O�,�pJ�������?�e��q�_ip��s��T>��9.���n�*��ڀ�Z�XbϷ�·�h���6��A9%�	S��,�~[n��|�i<~ A�sX�lH%�U�vjdg�y16��Ee}���婠J�u�FI	C�P��P~S]-pa����!�8����S�Gv�y	"�����+pZ�J懄�ǱwA�W�.��1�����-�A-��*,�:\=��Q %�`��h�_�Q�ʝ�Ý��R�3�?�F��y*e/@�)�U�x<���g>����y�7H-#� �`�$�|F![�n�;���)���fפT�b��q�\H�Շ�H��.��b	�c?l��W���T���&͕����Z���ʟ� �C_[1�~��앇U��Ԕ�
�A���PvU�d\X���t�	p'�����Ȝ�����Q�H��ʵw�aI�OCWv�!��<���^���h��w[	��HW	�kt5��;��}����US�������"�( �L���[�(��C�o@˚E>~R?NoǶ�$�I�����ˍ<���'�����yLE� UK=��9B�������N-��q�V��ך�yG�7c/79so��y��Z������2�տ�E��B0e �L\�6�@ͪ���_h�JT��%�V��o�<~O�N9� ���m��g�T�M���Wd�j&?��I@�`�/g7�J)NR܎������� ��2L<G�U��_K�/�Z+=�d|y�Q{I�����Q�I8�<X�h��z<��c�����v�	�e�����	���Ɉ��
<L�#x'�B���<�GO����t�T����u�ISq�MD�dD:p�=�[�{b�[�,s2�O�b�,��|O⎟s�vuF�z�b�~m,*��ܦ�$X�x������q�T�y�'Ɍ�\�T����,��-�0�t2�V�(.�E�b]*3�Vl�0�~���i�A�b]��ܻoC"�̗���%du�L�`�"�+���Y 5C��%�#�S�T��4�f��
F(�zU3vo�Gl��3v����NZ���gT>�r0��Ӫ7.��ACc��7��F��1D�4f(�p&W|��q&����(�-�n"�Y��QnFO3KgN' I�cZ�����54f8��~3�
��i�Ͻj�<<GB�%ř��.ՖU��D�I�>]�ɪ����:
�L�
��~U����h�$]�LC��#�� ��V��a?�l,O\ӍWS� �@��=��M:�B�g��I������Ż��3V1PQ�����*�ա`S@�P5�"�џ�?��\�bq� �)�������G�d��繓��$\䪦U!Cǿslq�q���A	�$�Kd�+R�s�ՑZ��
���Tn�b(أ� m0~�帵��� ���b���!��������� ����@G���QU&��,�]�w�OA[��ڞ݈�����ttI3AU�7�4�����D�2�AH�3$��+J�?p/��kWQ���~RICVY{�^h�M��E����h^=���֏om_#�@,�?�!;+�2��PRMi�5�5=���j/Eq�=yf�ă��{�rB�=�eT4ZigdP��ŀ�"��aA�#':���6\Ukf:,�|�,8�}k�ye�F�����?%� �����:T=w{9=�G�uy�x�H�e=+��FF��g�/U��������cr��G(�u6�͍��=�:��J�Ԋ�czУ()w�A�^(�=��y�d��8��s�"��V�^�_xr�H[`�t��J(���6y�)�y�)Pmip56P�	��2����q���?j���Ʌ��9�R�����������b@e��g���{�D����
�h���Gy�8;@O9���IQ�D��bA"W��#���Fw���c�v>�m�=BJ~L��* ��N�����L�h����/�����9���%�4:�ؼV��	�}"�_x�z�s�������aȩ�{h�����)�ȍ�Go�E��A�*�`�N��p�6`��%��Bux���+ǎ<1�Zŧ���iY�ةd��HGzd|�=Z� �!	�.�9�M�#k�ϰ�;��nC�(E<Ί��9wOPh.�$�@l0�oF��L�v(�}A��߹�sb`N'��.k�Dv���sM{)�VH�d�r
��~5�b{�N�a�@"��.�f�����{t���|�31_�@ت�K���1�	�M��l�������6p�I�vdߺ�����M�=�!1j��_��[�v1ژ9|��]��̀�8���ԣ���d��q�8�4���D�5����� �(C�M��G�_�Q4AD8��<�&��_�+��7U�-2���4Ҧ?�a,	W�*r�(���J��"foq�+~eER&NY8���l��P�
�fۯX>ݎ{��Vce�������P� �)��|oV/�
��"i������CqG��[�)��N�`�W#�z?��U���n����M��������C�o�1�s�o6.�ǂM��G�N���|�b`��u�\ r���c���%��^X뮶>�x�+AB�ﶠd�{�TnDx��t�Ӄ�0Uo�ŏ�Oj;�2�X���NxL�s&��86V��kv�S��L�T��<�P}�U�J����p��Ջ�~!J�5��XgQ�e|�0.E3�?����7�D�&��}���C'#�"�18�h��:�C�A����LXG���SQu�����+]�����fu�]!�D-<����Hg�{8oC���!��=��:Dh��,a�Mk:��~'���e��JzW��uܒ Q'ܵ^I���9:,�����}Jh�V���G�crv�fr�{��i�R��س����08����䉹gg�J�� �y���.Զ�x�AL�IS�������?��qg�?����{��2��_Ts&6���w�K�����竝�5��J�B0�Z=�^��Q�?Lf���}�=f=ˊBnN����WFm���q�J_HKoa'�Wz`2�=�����m�<�؅ǹ�p�n/��m9�j?�a�n�oǢ�4�C)6�49�����i� Vn�l�%TH�r@?�:�V;�������}��?�9/d����2a�_���h/���ߊ�=���'*l��ܽ<w��q4Bb�m��Z��7�X���3x��M�� ��$�PU:�%�^�e��J�f��F/C��&����_���	�i�0��8��a�TH��Y�	�%�\����d�z����P��D����=)yu�,����0�;zڧΚ
��ЃEo}D�Voǵ���k+�^〰��ZB0^y�D�J�Ζߴ�[<�nc�����{��Y~@�f
\Ҁ���`����xm��V�+B(�ߌ�ɶOl������ʈ��{ޭq�o�Ye�{횂=����`���G��a�~�LV��ϣr�U&����\�K\��O�e����P1�6������$G���1�՘Q0�'27��ʱa�$���A�#_˴�يF�����l���'�&yFR2>:���=����$h��%75[F������Pنt4��h���dP���%P����9'�<��eB�0n<Q�q�,y�'U�x�;���&}�^7�_�59̠��h�L����,6��Q�,��(��'C��#O�9xI6y�m���?��5G���"&�=��1YI1�^��:q^�HF���S!�z�RɼZ;�+��3X)�Bd�~d�4$b�ʴ�WHƖ�A��O�p]��xx�\�l���hFU0_P]+|���3nB��K	
/��c�y&�U`�f���a��7�F`c�:|�;��)�ɽ|A�2F�̷ =������Gq:��}FR.T�d�)�/c}ʚ��A�eYZ�~A:���+���]�O������Sh���٣��`��6����(Ӣ�٥{/"�80���c�/��ȴQ�dW
N	|�j�|F��[ل�E'YdwEp�/����m��C�#r肌8E&�+����["lM !:W�`z���j�7E��<]�@��N{r8�~$|�G�G���+m}��� +�>�Sa���zHɼ�N�H!�Y+L�(����'����Ǎa�K1�\V��?�K�C��ݯ������ſL������A��*,ew����h�(x�`Xjp}���.UNq�*�uN�k��NM��KZpG��l����)��ɐ��L�t�9v�h	=�0���m���m����)0��9A�R��q잶��~S�s�+�0�!���	��,)���;��)�9���얗_�s�.��}��(V<�uO�i�����"�ꄲ��39t�ݱ6����d��J�B�;��\����t�F�]�T�ϓ�y��uPھ��V�3��3����a�nQ�ŉr<j����E�#�3�bA��%�8%R̃7;A�e�R���{sǹ'�52���
�����m]�)�|ٵ�Vt[g6����zKr''7-v����.��K�o��i�I��2|��/�AQv3�ܕ���L�e��B�.�(�{q���AO_"�xB��h�׀!�(4	y�zE
0�˜�f�ޤQ
�4�Ƌ����+[��7[C%�#�
݉y��I޲�>�1���'F�t����!P��[����x���d���\]^��0-�p����EBÊ��=j563v�Q�Ǎ�����d�N�Q��fcU�)�ߔ� RL:���p9�s�]8�-/��8[V��A��x`�*\�0_6/� yn�Z�wȥ��DC���|��<�u�j��u4iz~��ӯ��H;��p`x�@������� �O2�<-�[m!�j��1�Ô�@���x2�P����T��
�c�r����2S�erQ&��}N	�������1��㝡��+�H�׍�`.B���÷��V+�kh�$�"��lUc�BR���t:��kEO�wLd;���"]�!�������˚,#��Hg�i.�"��K��,�%�Y��S���u���>vxT�ɵw�@TGI�`էt��72��4u��{{������*�����T�(���	�+>���`sd�At���~��APnD�D34�Mθ�}h�o@�.k��3J{y:�;�6�`�ٕ5y&PmG�s�Sr���1���ߗ m3�9�r ���#��rRMlч�S�Uqs�!���u�a������`�'EY��+�.��o��BW�W�f[��N<�v^va#@�6R��U��m ;�)���8?ؔY�),�_c��E��:���q3ZY�8�� z\��~���B�|�.ke��@���@#���0�9�B>�]+wj��Q"D���|�N�a-��5�`I�9��VZI�X���)�>�.fK��ۼQ��@.J60m�O�Ƥ����@Q}��HCo�e���{�-�8J���0�o1��Ĉ'���s%����
�[j�o3�r��[��bʏ�u� ��a�i�ϡg�ɽ��K�@����֬�]#ÑÌ��� �z7�mĞ��>�J�א�W�[ه�iTY�V~K�h�����ρf�?S0o&o�M<P�y/�E������[�D�Z�:�%��BNY�5�f�W��~6���t���v�C��)�3ц���܉��K�=r�����R@���\�uEXC�-��l��T�$���D��k����p3k]D.�r��*g����`Q�ihl�M�iBև�[R���扱��]؋*G��{��u�_jv5!�#��0��f�X�>�O�
@h�=��{s�Zg4�k䮬��šZ�2n��Kh0/�I�?�i����a�-(#,�9L�� k��jd*:Z�T*<�3٦�_�>={�%�@ߏ�4��ІU?�N`���|74�]��r�&q�q���2*T �OW�ῡ'-�/���t�����jr��.s����D��<~[t�')V��S��I���%�H��5�CaCٸL$ˠ8��@b�;b��ɺO_:���j��T��?�2�o�+�N!�y����)U�����6�Fȩ�_)�l35�E��Q�ݿ��3��8n�J.H7���?��`�������t<�WF{ف�T�7�����-l�O"|Wj�7a���τ_M��Z��鑼c,uߕ�n�����{v��m�=��@��"p�v�:�>�=�LW6�F̈��]~ B��U�<���<�L���.���ĳ$�x�(j=�l`]L���Tb�fq�ь����^y��&�j�l�	��t���z��q\��:��5�;��(=��{�]聴��^�T>����2{�����^��^��9�	R���`��	ǂv�H���C�q��֩�xX�6A�a�RL�&6B��H���zn!�%"7d����cwwM<�x��<*`�A�@�uiy.ۋ�?�"��1hǵ&�1(�ͪ��I��Xܻܬ�5�)=B-�7�H�J�2Zx0<({a ���i8��yۄ�|C��_C� �JU�ч+Dm�R�H�A!R���d*�f��>���G.�Dr¼���� ��s���A&y��PV����"M̏��*�{q]�����7eW����S{�aO��Z|��@�
�5��G�6{����
7[���N~�~)�.���f�n�*�O5Е'�ϭ�A�����D�OwJr�?yda�7�B�B�׃r�8��p�eg�l��bOp��.�����"�z�(��֮���`����`@����s�<ZӇ钊����Z��P�/����L�-߃� ��,��čd��:|u�k���CV�.a��`���S0^����ƥ@��\=g~QV^UO��S󂑭�'9>�(��L/m�;�������0�~h'��H�h�1x�}�]4a1� ,�����:7NS|� ;Q��zG�г�^���t�.�_c2~*sʹ�E�Ɂ���'�3��t�7g��m\��t�ɯ�x� jh��c�f�gr���[��c�4ޔxa�Ͻ�m����8dw�w������S*���}�JZJ*�8�@]D�{{�,d6u4X�4��x^=ø<�b+�#��¹�G]��ES�gB����n��@�-^���N;�r��Y�{�a�v�l�����+�(oYe�Y��IV���&�+C7��EغMEj�h�H jh�Qp�Z���I7�g�V�5?��i�R�6^Fͧ�vb�Q(�A�lz���R#wmc�`%iU0P"�4�,?I������I�ga�=�I�x>JU�7w�,C�G5؇%���cH)P5:�٭��X��N��dJ��h��z;hC�13?�O�������f���E=.^uت}(��r�q>_��&~�����[lFF���۴c0��Z
J�<l�9;���mɏ�P�9�q/��u�p�n/�^=s�BcYE5=�/�`�c�N�`�keʉw"t��_����kq}�휷N1�OG����j�βU��q�
�WiZ���h$խc?(��r^Bx�йO��:�Qc��+u��V�?މ�r���h֛�J���y%?]���4c�����# ����*a�v���ܞ}���-��E.+vW����ͦ���Q��}�؛S��xN�R����f>�aW�0P��Щ����:�y���-6��t;�秪&1-����>�C��x&�Y��O�z �i9���ӟ��
y�� Cs��X*e��R�} ҤY&Cy���o+?�eVRü��<�0�9�����=�R)�3���4\�2n��% `�@'"�,��F!�
Λ[�{6��Ȧ[��'�c}H�<_QUu�F�u�c����G����̓t��jKW����rw��+R(�AeT�`�Q8r�<���yJ�����\�=i$�~��?`6�ww�xFH���a����	dmv��a��B=��j�0�l�m��J;[�L܈
��n���hD�V(g� Ǖ-X�7N� ܾ�9
?��������)�P"��Y��aXB��;��ԃ	�취+1��P�:X���r�~�kQ�J�w�c�ׇ�J��.�OB��1����#��H�mm��㐺�mW�D�[�\�SY�q�Jx��f�t���6Ǐ��S)�R����&n���,�6O`�3��o���!�'a�Q��y��h�y�/#��J�_�e�zTρ4�'�����3���U<Sk��J͢�9����D}E���1���k�������Ҕئ�r��IJۂj�N?R�UZ9+C����9.Z�6&�ڄ�P�	t�өI]�É�u�g��a*��꽸A�!n|�7���s����Vm�7ԧͦj�<E�`*�=���ʱA�	w��^r�78N��籱�"�ն���i��� /�*�z����,��ttK�2O���O6������z�y���X;�2�s�p2��?���v�:�҆:������Pe�q�&�#��:bޘYI!�����$ݛ`�$Y-�L*�u�m�ý�)�o��P�������d"�-��u�
��� �O ���4��=ք.Tv�@F�����o���$R��S����V"�F �ڊ�����B5�rgOl8y��e��2��k���<<d({J�[9�Q�9'`�n�)�|�<�P�&�K�܏L��2S[�e�����,d�q�Ų����M&�l���;/t�}���u(��hoʊ �"NW�ZM�\6��/�a@�Yd7I��^R����In�ɃG�r�4���{�s"�.������v���i����$�^����&>���^ʐ�N���ܞ`�2a�9�����]��t���,M}�M)+� U�+��ߢx��,��M��S�Y��	0��0��ʯ�����4�4�F'�Ć�=q�cNl��c�v�wǏ�̟9�L��gKe�"GR�\?:�m��\�iv7�pn(8DUD�6���AaiY�.;��HV>�v����������;�v��y�t�ά�XP�d��q�/���밅hh�'��;l�`�jg�5�;.��2HJX�C�}
�|FM�B���)d˸	�I�M"wP�tuw�)�`�Ԁ�~O֙Ι	�=��+��Jd15��1:� M�pwQ�2􎊔��N��	YHE��*׭:��m�V�5U��oox�0r�{��~(��󉯂}�����(W�ِ�'#}t�*OCJ�>X�����Cͻ2�SZc������E��Xz�r�>᳚��(���\�P0���W�+���M�҈z�8=)nT�闠%j_'�A��X7Yp�tud��t���g��k��b���^�~�N�����f
W�9f�ٌ� �Y��-�T�9j[�ya@����OҙI��d2��w��`�K6-�tf�T�׶����C�֗����fA�����ڿH��y�	qڽ�����L��0Ӟ���0�S��*E�>�k�H��=5�f�ޞ	w��\�Վ��TM���W�	¾�K��%��t f�H~|V���6���zCe'����H��Ѓhm�(�@����t��#�m˵�����@@����B�^�m�|�;��XfWD�1�Ϗ&L��[�[�o�� ��@8���'7i�Ek^j���1b��3LXѪaG<MN��Nb}�[�z�YW��w� �z0ٝ2�Q	DD�ɱ߸'b�xL]H"4�0�]�(:�@��w��e`a��<@���<b)d���O��"%�!��<A�!оa&׊&�q�-�sd?�{X�;a�~��m4������.��>*��mF@Imɻ^�O7�]	�_4��9^�3H�n%��i�'7��^K����0�|�NģP�ݧ%M�<OGX��/����J�2J%��C���Qj��Ѭ�������!���(L�0�#d��u��EDu���t�?<-�G�a�ww�u�k�[k��!ap���"���li;+���UM�K9�K0Ѵι��_��7�V���J[_�,q����ǋ���J�f�CsV�="�	��5�)B�]�mCzj]OLue���	�k�bX�����p����2�rҚ����ƶ������<�8�yͪ|Fy�a�Z�4�;�[B[���䏼i�7-�݊���H��U��� E�#M&'Q&����L}�8�'`;4\n!W�@�����^Sɠ�T��������~�1˨���L1E�'�0,�c��D���x	JO$V{�f�-H-I�Q"�omq���/�-��$"+"�]k`!����)���|F�CKK��>(�^����i����hj����Y��~4�˰���7=ݨ�޲�ʰ�!s�����N�j�j=G!]K�b+~�j�Q��o��S���`�~�0��w㓶P͆�����\�~B����E���Vv�V�ͅ��Oo�~�(�ȝ�Q\���9C�ٟh-i��(�(R�jݺpue����Yfs�/���~��U����_���jX�X�Χc&�;'4��=��a;ȊD�1=mN[� �������?�>��۠irG=%� !�m��{��a=5�Y�G�#�N�,�xh�ͶH�G���chشߨ�N�)>j�C�YB���) QG��w��Z�Ʀ�i�/D�و�(De�^�"���ROk5�Ɖ�dT{֝7Av�ٍm�hZe#�"FL�5a���<&��sL�m��v�:joE�t�AО?�:C_��l"�
�-���A���ȁ�	g�ԅ�B�7�ѠH�cd
]H����/��A��J��d�"@;��7���69�cJ��E�9�i~�-2��}�x��"�'|���z��x�H����Y�)�LI��řH�Y�����Dx/2�l"��=-`�@n��\i�Q�W�-q]���L�A��H�1��4*j~c����չ`�y�/�����)�\�\r�Wa��xKI��9ٔ����9�Po\ŻN���֤��Tq���w1F80��9�#�y�c�,�L�V�8<`c��,�B��k�u��� ��}?�o�q��U?�rӺ�q�wޑ�_�r��!��uk���#�0�穝,2���|= cl����?F��^V���2cх_$���'6O��
��2��}ӂ�W7�"$DPL�p�;���'so,}�{l�J���3���SY&MI���L���r(aı����P;�_��-����C��zOT��d���5Sߟ�s�}��ۏ~4AEOe��!��L6�w��r�i:*e�rS<Ҫ3�3��B��C�{����;����yJf%?9��e��=�j�Vy��r�U ;}krc���Z2z$���:�\��܂1�[º��h,-*O7:|A�o�t��'�c������1ۑ�v�ü6�Ha�`	�,*�E5�}�\-�n�&W��b�>�V�??)�6�yt�p���u�?�W|�x�!I��
�ql�n��V`�7-��E��#'&��a�F��LC�m�j��`��Wxg"��7�nN_FEv	9�pn\u^
+�K�4��j��8��G�j*T�'E~7䜫`�_Ȍ.��Zm6��i�}ޜ�V�S��� ���=J�f�g���ev$:�f*�o���~С">U�e�.3L~?(��O!p2�'C����T�Ad�p��X:��H0�b��L?*S���u�7�W�G��`���3`iMr�|�m�g�\��\{m�5Ӯ���3�u\N��۝�g�M�}���K\�q��p�J��?C(A_�5(�yPBڠwFXA�3U�����)kGG�t���R��>]Z�&�����N�S5P����JM]�����!0*����4�@c~��2�[s�?��΂�H����W��
?�'?�S(�EvF��q�,�������[C|�,Pʂ3{K#��a�c�xn$�rOC���1�<��������0TH����׏9������H�^7�2���=c[�|�]$�".�EY��1l1��*�H�r�u��,=�n�I�{�i��X�W2��J<A��5og�4��7Q�礽g�"����8�Rn�]�3���u����X�ns�[7E�E���C:���S߻�4�%��96�&�TOX[�]���Z�/R�H�Y̦��m6 -S�!��e�>y¼"�J�H<g.W�t��6>���
��DJ������	�B�^�6Є��1�	Oi��W�t����J����+�C�#���1u���*�����M��Cno�J/c(�R���� �����ۍ�}'�D$4�$ �B��7+��T�Z
oeiΚ$^����?��� �=�����D�PF�p8Á�w��^�|;8���2y�k�J�&����?p��D���������
���Ώ����?U2)��I<řQz+�zZ)����2�R���%�y+Whd�Y{R��G�k��1���e�,�,��z�����YCF�N�H�?��{�F��7Q�R���21�ы�靏u|i�n�ں�̼��ƛAU�dZq�m��T�(]��*g�O�rQ�1�����#e7�.���Ҋ�EG�F��N����}G�Jr���T�4�Mw�A�a��O�K����)���H����M{f\�ޏ����~bG�~6�KU���l�4������eϢ`�+�3nDe�迱�{7EhKY���U9m�(pņY��5=l�h�`M�/��C;�ey|���}������J���,weZ�@��m�Z�u��Nl㾀�%�Bmc�<�Y%��FV%�&l:�kܟd�^��o�;����W�X�H�R@��!F]C ��[R-9ذ+`���p&����1r9J�hg^=�A�h{`O
�3��FҦo���_E$��� V^�]�ho�`�Lx�x2ˎ��c)i�7`�0ӡ����׼%��G_���s��C�˖f�M��Xi����M��H�ƽQk��YZ�������U�r�4TTS�7�Az�r�]O�
�pN�G�̹�Ŗ��,lFt�y��1Xsë
�cϭ��ٳR���;@T�BQ�RQ�d�`+g?sԢG��=R�#���7H��q��
^�e[�<;��aL&�F&�ea_~$#QܡgǑb��ˇ�2y}��Ut����^q5nEt��ɼ8m?���+�,i�-�Ȼ��J�pM��Q�����|u�|3'��2)�X��cBafYe� ��v�����4�8�=���[�ҿԄ��8�w"�8�K��|췙`�˨������,�}ff��'�$1����w��_"���َB5	�xm��G���YY��,H���Rz�a�EW���Ǻ���iGK�����$Z�l� ��A:���L�0:��t�t�-���F�0�(�CYJj����J=A��Й���{Y6���N{�K�lV�5���l��_�f��Yצ�M�aH�u����j�5|���7�ar��T͈��;w��V�?�D�g&sQ��>ki��R���������8kgq@w)a����r���Uذ������>f,ue�7���ې�P8�3r^U��F֋�9��L�='�Ye�������|a�����i��E���f���h>�=�n�r`9Kƨ�aKi�n�]%�n�蘣�C�B����Q��ؕ&�r�m�x�N']u@�p�q�nv*m�qD	���}�?�2G-�X��-��QM�O�,�L��	<��UG��=/[2��9J<��������� ���fd�뺁o�+�J�f3SBL�w�̬��ݞ�������b��(��� TH���J�>wQPR��11���rxT���.�z<õ��_KMZ?���j����CnK��K\���	S��o@a��A�G��i��OH*[�en1�3v#ޝ�������[��OQ�q�*�(Y�$ҏ�$ߊ6���d�|Ͻ��g"�ُ_s�<@xu�����l4�[���
_
�w-Ċ���+�<$1��w?d�b�'W�'��D�(�p���9
ь��Yl�dK�^���تг�\�w\L�Q+<���@�N����)��E���M8YCιw�<��>YpЭ]Oe���9;�$�^U�<	��,��޴buC���h��q��z��������ܻ���~:��)z�%�{��.gsϻ(�G�/m�|w��CXr�Mw�+�	�*�9�k�v���R&�����������5�P��@�>�_qN��k���Du�9Y|�B��#�Ƌ{Okhw5@�Z�c���b��"�%�K���E�pb�y~�H�����L�%��9����M"����9D����S�N|Y]����� ��$U����g���NT�u�(�=�X���<ֳ�nO��=�2���;��\LmV�	�C�*l�OV��-�?�0�tv5����K�ą�r.o�^��0���t�+7���x�?���+�T0����4�Y�}�k9�>�>W3Q�\���u ���c����s��$C��5C�nNUQ���1N�=��>��rV�ǝB�)K��7����}[��<�EzHsb��GS &p�Qa��*M���c˃�*O�f�~�91��$F�IQ�	&���+pv�p!�sS#��G��ǆDj���N0�����>����iͬ􋝴)^{r/��*�+}U*.Y |�ez�1��lS�b�I�T}��)�:ZJ���`8HL�վ7��Q4���[.��$�>�K�1㚜FI��ϏM�;�J-��e�r���c=5𪌊Am"G�I#�xl0��h��b��Wtd��k�;����E�H"W�F�2��,�|-����oLx���=J���Rbb�-t��O(�sJ�
�v�fM�7a�uG��(���D�)�o����4�L	ز�����pn8ç.��1��c�'x.s �W�#)���Y�q8�\I����3a`�GJ��S���gN�/��sAy��q0���{�Dt�U_�K�0C5�	C��S��<�W��zJ6
���V�Ӱ�˴Ry���6,,�V���}@S�O?���y���*���t/,���^gC���B�Xw��\(*��LF8@Ts���j� ������k�9�{߱�Lb�gWS[��H�����s7�I ��Qɠ���z
.��6�潉ݲ�[��up�)?��,��1),$٤Hם�fb��RA���ˡ��C�Κ�'���F�֨�8xg89�@ojy^��d�&���B�M�b1^�J?>[������8 !�]�*J-���-����;��,M2JgZ�ev�5`4��9��ܴ���iۧ �������a�B�t|g����zV�x��-��4�8�/r�dWVA"y�<�g��c�؄Y��sڙ�2���"/�K�ۅ��	����r����ҽ�9�� ���3���˾���2S��E�C4%8Q)(F�ti�]��)m
��*�V�Y��<�"�mn:zbI/�$3�9��ѥ9�l�����Vx����w�Qrr�r#�wD<��{m�u���ֻΗ������܇hh� �L)��3]MH	��Bu�@�Q)x�@�y3��Ac��x�Ws�ѓ[��4�1�zӟī�/��^�o�dD
���$�)����z>�V�=PU�Wh��qs�D���{l�������i!����M���Nd��OlH�|��`[\�k�ȿ[b鎩 ��x�CEJ��s7ʌUćbժ>[�bz��H.�Yb�	Ѥ�7�|�{�ίf�� x��Yu�Eʅ��ںw�aI8�[�&�b�����c�o��va�O��`Q�+��|����{����{��я( �z`��ya�"�I�\.+�:r�z7�\�PѼh�A\��6q�~%.y�YK�1����H�w�>G��������N9وW�SS�(<�Xd��k ch�!A�ir�d�K��'��\�^�4��Eg󫫰�q��@v�����(�(�{�RW�GB����A����Xme�%~962�e�7ĎwnV��A��~�����V�%�Ӂ-�����t�����'%�E\�:��CS�O��\a<�d/�\�����rq�!����	\�B��S�߅KŘ��L����f%f����>��08)o���s߶l/&y�Q�c����M�h/V�����ƥ�a�U��H�|���
]&��I}"z�\c$��R�dR@E^���3�*E�N��V���i�et�ޭ�C��5�0�-$�����_2��NOU�櫣5v���عҲS?���ʹ�������Q*�o��2������#t�7s�3��Z�rin>i]�c�p�,�}?�o�n}���ؙ�������f�WL>`��JvB���4V2���eS2��c��~g� �=r�J��/��i��RۍþiI�qp���5ײ�ݾ$���2�K���X����G�ٲo�O�C`+�^G�-�5�G��������x���ڳ�~ܸbNH������ �	�i�ɷ����4�������E�&+P5���6?a�����hj}i���ʜ�R:δV����c� ���,��P������ ��w���f9Y���QC-�1ޏz=R~��X�C�y|ڞ�=�Yc�/�m�Ip��N5�/�5HL�L��v���1請@�{���uG]7Q:�XԈ=<+�d��!�Z�]��#T%
�%�Ż~R���ɟ��g�[��¬�b���0��fDN��%B���s$��<v�X$���Zl&0	�/�Ӹ4����
*ͤ�2"tHu���K��R��©Su<�c�>�>��ЎR�������:��3�4�@<�uF"��L���9�%�C�	��H@�JCk�M���iv����~>aF��5�ҿD�sW|��;�6�gw�e�@Vh؛��uRKם�=�iT���S���� G�ŜN$W�'��i]�,�8�B⥾���h?���xً�7/>_1�S��$oL����Ƒ�ԭ��'=WӤ�c�92	w�`,wQ~�DL�@��u��7X�j_��L+.�,�
�k8�X��1��'2p����;�.�8�n;y*�m_o��r�3y�o{��0W�D��}�|&�ܗ���+��^����Ʌ�
���ܖXYL�s`���qa��Y�?_�|�h�We��$Q�9��c���
1;���od�:)��E���.�^N��`�=�+ H` �O���4�{[	,�n9��J9��޶�]kc�,K���b��2*��A�T6b>R޽�iA�B����0l������i9U�.��2E�l$�kz]K���xk a[mّE��SD�,#/Ҕ9?�rB�\��Re����T+Ryj���8\����P�7�܃0�W�!|E�,t�[Y7��7q�"�qdT~&��n�
�GR�k�zF.oV	�^Ha'�.��_�d��2-�� ����C���X��wI��E�w5�A7��u���W���2�"տe3���/)�o���wi��ֈ��$Ɩ^��#pnK�����GPm2�2��,#�z�F?�{C?͗ZQ�p�����>4�Ғ�_l%=fpY�)���_��_�Ŋ�Ym�k,��ǎ�қ�[u�=w��k������7�oY��������+����&����
��r6�Vh@�"��u���8$A�C��!��B�+o�b��#�����M���z^G$O
�%w�(�|��%,-���d}z{��P�8����Ն���
d�?:쟍]:��GF��]��Y��"ܤ��3�Y#���Z��dǰ�
>�'� �B���
��L���o���K¿K�b41�d��7��İ#��)���?ء�l�1
�n^�4�łt�8�O����'�4��Y��m$z�~�����3�����u��e�P��ӛ@��9�Y*iRy��DF2�ry�72R|��R>*��و
��5;���ۮ�n�c��ΣI�߀��Y��S8Ў��H!@�N��~Lx�`�uA�aWI�-�Vc�@
(���՞>�3Ot�	�s�+�۱+���R��|mPy�Ͱ�&����5�4'���������3�֬(Q��F0��s��
,[U��	~�?ڤ�7Ϧ�r �!)(���@7"{`е��[�{,�
�{�k�(����B<��j9x�b�	�7�$�k�� dԒZ�B�N�&��O-0�����f���$ZCӣU�|�y���jBn=�3v�I�s㻦��E��LA.�SE3���J@���躥���9�0�F-���՚��vĨ7�e4щg�^i@(}�X�� ��$��<�t< o!��!������x��r
����v��b�g��`���T�+Q<�	����xO�8��SL`='!��x����~��6Bg��f�̽������£���ݑ�<����Z�h�`W����c��9�eKe(�ɚ��O.R�j�a���|
���<���m��-�V:q�F����z�KU��m� �3����5���ç��6�	��˷��!�����pg�)c1OeI�h��AUݵm�q�q�ȓ�@��b�Y�d�'�����j�{Z!o�l]�{�F4�Q�و�A�QV����R�!5.��gR����̈́Z@��1����.��G}}�ٺ�Z� ��eb�qc��v[���G#��OM)���'ʈ�� �����!#�7S�����0�CV��3�� ����)�>
k��8�Z�a8E�`HMᆈ0�z8-�$�{��Ї�º���K�Tbv9�����*�#�ػJ�����L���+�>�p?yR�0ߏ\�9$��B4��kN�4�j)\v�Zy�M�B4J7N�E�p���L����!�
U�a�n�K�
�Y����H�ヮ(Bd�Π�F	�P�-�q��_�hi�"��� :�I�9���:IFQD��^���	\NpLr,��~�S��3�a�7��zON����ר��<؀z���2Jw��R���4v�G�̼���N;�u�_�h]D�	�* �#v�q��R�]
4� �dm�Y�4�I�A�2j�`�nwX� la�l�.I����Q���k�aʒ���W!�$�l�d*Ү#0)|㹯��ER�l�8��Ud���2����1��$�Q�H>|m`�K�}��te�����30�1�M���p���]_ �N�J��o�Ԭ��.%��X=ϊH�k����L�H�zHo�{�J�HE���kΥ^=�h�|���oA'	��d��X�Dd,p�G�%ig:�p��4���\��[�
��(y�D��A��Le��NĞ�,�!�YSTyl~�֭�d�y�
p�[����"��<^���}_����A��N�+���WQ�,BσE%�"�_�O�;�u6�Y��P����+��+��SЭ�/�]91w��o83х5��]F^$��h��G�$���x�x?�,]���)��*����K��:�)��Rn�C45�кTn���s�+?�(;]U%�K��r�j8~c�jg�Qk����:�������0��mU_��=�.���0Q��b��#�U�H"z+�H'Y���o&�wK)����������}�?��h[T˚���'=��(�]�h0��l�	��}�h�,	hMj7����R�YQm�W/p.*��fW�ؑ�5�ᵲ�M���S�c"k����Pa`l�@�בG�z�JFT�7�E��&4�./�{@N}І:XB��_J=�Т�ܑ&3��P����xUс�7�	���â۪"k1����*��Y��m���V�%Q�ITSjS�V�?Q�JCibs��jFoS�z 0��;���C9�i[��A'x-��$
̳�������
zBJ|R_��Ҋ0�%^(3U,\{]�P4=#�D/��n{���ƨq����6� N���m�����:
�b�O���QX ���L�⣏�ʄ�$ �K��e��1� �����D�ڲ�:""S�<UD�b�gw:"�_��hW�1�鸣� q���;��P�E�u�0�A��_s�N$��Ƥz�<~cڷQա�V(A�Oբ,��헨L�����I�;��&@��c2��1Q��Wz��*�C]T�j�cB�99����6�36�ξC��ֈ��:����+�b�-�~��v{I
 f^"�窵Y�U`�lq��y�i��^�Sѩ;����'��]�5h-.S�����b�U�I�_���b�}�ؐ��!�+d$�E1d��쬗q�ݡD����2���X�4�����+�j�#5b�g�
m�fk��"��Y8��2DW���)�����o=��8�
 ��"V��=�:օ}���5?S�S��F��	zJ�q��7egE�Y�ׂj4�N-�S� \��82�x�~��4���R�c�* �,��l��[�,�h�M�^� �|�+<'���4]4>%˟"���V4�B@�F��z!bkӍdQ�h��U�|����Ͼ��G\F�3�i���9���/�X��N�:�+�S'/�)�g�n+��Ȫ��|r��mY�-�ǰ�Pڤ�~i�,Fy���y��`�
~O�2']V}�����%Mt�u�p����:(��S�1��Y"$��woOh	�$&�3��#qYSM�&J�^l�v��K��)��T���4b1~�N��L���p���/�%�&�����}c%�H�Uz�aK���;O$��)4�M.3d�p�
��/ޠEAL�YEo-�dxw�ņ���n�����2g�(��Ck8�7���!x׽��(���SpP~*0/f������'d]@����Ü5�DM�{�z��|G-�	�X5:2;"�c�>��v����G����41~+��E[�$&<.рM�ǅy��64�`zxM�P�ٝ'C�0�nF���'�� ���I��X^�>�mZ�p#����C8���>ty���
0ϡX-���_�^J}�D�a�[��Ʋ�������3���-aI��������B��a���
��*K"MXqXq� �a3~�߱�5�W-��U�W�#�_��X��K+Cޣ���$�=
bl�}h�H�|2�G_� en����J:�	�9u��>@�i*"��6OV_G�=z�������}��P�:X���1���Vgҍ���fX��\���E���N$��p���\��t]��$ф��˗y�.5W�A��z��hw������A"��4�3�H�;t|��oj����vŢ��/0������H9!���*����� z�Z1��Z8��+�����7��D=S�����l�-%M7�J׆�P�J-7)�ѠJ`�5���}����ֻ�z�@��$�wb�U�1�f|W�y���'��vȃR����KQ�4��,�/ʙ��g��g
�=���l�]}c��}@.Зr��
7a��6ގ]0B�9�|5��Ha��j�g������O�-���,f�2�)<'��ޔ=�#��m��P�G��Jvumn/^��;;H�Kףl|R;_<����b�O5�W�Ϥ�
{��[r@륜���d����]�u�8 �%�4�Z��AΎ��JZ���S.A+�i�&�$�k�}n��RT���]�����~=�ޣ�DK��>��wD*�1��	��oaw�j�7F8i��24�X�B�l��� Gp)�cm ��Ab��h���4٠��Q�8;��-��iA4=0��Ώ[�6��Hf���x��lV`�t2-$J���`�"����]i�Z����ۮ�ɝ��3nh�+t5��%&;!j�������Ja��9>���/�x�/�M�0�`)}���6�5�ҁ�BI�%8O����K���tX�Z��s��h,}aU�].X������Э�/M�x�N�uI
9t�qAO�؞@	���(k6gm��I��O�����U�'����@�0�{� ISYR�D��1i[�h~��H���[�v��w����[��bG���5�'�9`�E#-�T;SfaLf�E�'��sʕXf9.@Po��cgJ�/J�=5�y�,�Ѯh%���6�Ż�j���B�Ȕ�>�ץՓPg�'J��3E��A�&�1#�Z�\�9n�XLt�h5�Z楴Z�m{^�J�kxŅ3ZV���(�YC��gע�`���Yf�;�X�h��ݛX�ik��o�w�$7��~��5��_�6�P-�Uk��߉��� g*�ϧ'�T{U-<�^����>M�����eF����[A��SR(.>r�A��e�����ӚϙN%<ȕ�ݝ�N�i�����>1,~�i�\V��I���lX��$�D��QF�X(��w[i�i�hnW�y -ƐO�$���w&m҆�s���0*��+eT�S�dx4���1\{�&ȹAYC�BSd�'x��U<�e>��B�ؑ�R8�� ]����ZC�$֒�� `���ΐ����5���hC���a�+$p�p����S��r��ϩ�c"R�?� �0J�ɳ)���d&���rK��\qȖ�c���D㣽&U����g�_7V��8�7M�י����A�������)Y���ño��r=U���#��ĹB���������.�ȁ��K�f�_D�V���#f<>�
i�o��j�mS��L�;� {� Aa��}����yX�<����4�/r9���P^�k�*��'gm�����(,]�hg<gߧ���P|	v�I%͛8�Ǜ���ܜ��LV?Y�����(F��$�"�βm��|Ӑ�⍍���9x�N�4װ])�9KҪ7t$tH<��Y����5�.܉a��,�R+n}1�2�84�r�w�ºd�t����������9͗�A�QB.= �="VY�W��,<���+���xI1���=]V-]F�wZ��K�ح3槫��[�Z�~8��Z��\ӫ����@��S�fo�Uƾ��E=����Օ��;y5��f�������H9�$�t&�,F^r�I��D��Ӿ@�ٖ�:��m�D����8_�0l\���:`b2��6ۣkH�͝(��į�uNp��e_��6o����e��f=��0���ia�]�y�O��G�Q/��G�%�(�3k{ ���L��GKg|g�O׏���wA�d���AS���ێ��Kډ(<�5͉�@
:^.p��d��1!�g�kt��ٮ��U�D0 �~�[Y]45^g����s+Gb���s.��?a*�'�&�>���a]`�Zm�����^����nR�|$v�E�[*�&'�H��{Ļc؍c�mo3��¶?�ɞq�U
�p�[��.J��k�҆t����}.2�"/O�C#��[�dЊv�QAG�(l`nn�����^��F
K!�97,��n�yL�A�Ъ�C��%�Y�(X(NQ�)�3�T0��¨cW]�����u!��ޤ���E���ضԱ�_����{�m�,�/�������`A�h+��������\��Gyu�hu �굉�w�{u{&�^����B�}r�.T���s��z-I�J RL^�7i�"{�p�{�v^�ՆaG
�l}����G�:FH��8@��R���K��v�ӑ6{4�z��m	�}�ML�C��I"��B>����������8Z4c�[�nn����F
���w8E!_[︮�_y܉�,O�B�]A��l��?�C�x�O�����*�Z��V��DLHF��<�� ��J>tO�U��ݢ�����Ü�����\&�´K�A� u� ��A���|�L
��[o�ZO/�,�Nꥆ�	�?Z	Q��(�YK7 l1�JH���Α�r�m����t
]�gb��TӀ�=,Rd"s&]���\*�ZZR�4FI��L~ug������n�.Z@Y�Iϡ��z�T��4sM/����g�R�����0Z�L�V'����=�|�������g<�Ã0*�R��k�q�;x[�ϩŋ=��qaE�����$,�x���ǫ���k��d���N�e��{��b_���-X 9��� ����b�c{�?�:Qݔz��7��Y�d�z���=
���C-�D��Ւ�lrJ�{�:��,\��:�5�Ȼ��G�Y�nqQ�)z�b���F���rϮ�8�O�t�Yl/o��b7ܘjhi">�z��'���e,����	ST�� ��hȨg��uP�۴c�SBm���h~�]�����s�`CXS���J�h'd���v�NI-f���,�"���z�,N^�͊.X�ufuʠkVap����v�#��%�~*[�9��Ìb�l���E��7���U�����C��=\WE�Ԛ=�PĦk�h�OH9耘S�~�|8�;1�F�E[����gF8�6�~K˦R�d�?���ka���J^y�t=k��~�ɺ)�^FYWG"�R��U�0۸�X�q��/����m�p�л㣐�g�M��Y�����"!�fť��|Qq���N��Q�{e��2Z�¢�	�[S�&�4I��F?������C���ڴV��N����� �������N�{�'H������5K%�{�K �GuI��R<k�G-DZ�N����0���58i�_��9�Q���%ISFS���Jm�G�<",]�a��h�.RЗ����)N�EVߜn�^I[��V\�Jo��dҹ����G�t�/�X��YN��D�I~��y��~�
�8���}�����0ލ�e�U��@h�ˍKI4��}dEn��7\"��bʈ��@��=�QA����"7ӥ����&�+�Jy>z�v����-��������,��Q�b�5��A�fs��|�:�6�Z�oH��ZkƧ�M� ��P
���=m�O�T �i!|��[���Ȍ~Z�˔��Y1��܅ҋV����q�ĸ�s�^?9���ƭ��8��E� bR�d`�s pK�spV��[��A	O�)�{o_��Ot<�<��]rsA�⿃eb}�_�bTi�<�Z9�%����Mn*U ��T��?�T���Q�L������}��g��
�Q���l�h xh�t�ǘ4���ׯ76|"�9ƀ���V])F(�w���L�!t�PA�_������q_��<M�?��X.�����(pk�v�q꾱��6zDN�(��) �n57�Hho�c_�r���$�fCsI��h��z�����,k��Q{�a�p{�k$�|�1!-�fD�-�^�v^�YNC�3��`�e�a"��Ds�|�+-<�ν�ŷb����ۄ��������oe@��.�J���fv��9f�� A���tIO��J��9aLc7�ѹ�����p��$�,���r�����N�ؒ��=QȢ��V�?�BѼΦ-�Z�e���j�s6e`��d��K�L �0���+���*/5�ON�i��O�ҧb�Q���&���L�R	,�^'hZ���Q�E/��}�$�m���M�
���!�3��H����L���U(�KѰX��)����es�{[�V��C�4�A%{�O���y�Bs����d��?���j�<?���	�Y�Z��0���6U4����U���G)�n�p����=n�4�0��N��P(KZ�I� ��x�ᑿ�����2(��b:~�,%����?��,b�S;=��_qN��5�m���֠v������4�V�N��ݶ�io\��C�QMR%i��.�ګ<��3;�sD�i3F��:қIK�=��)�w�oST\���[�]CTw��H-	Q�"�;/X�y+6��k����'.⊽��چ�J����9���G}^M�V�X=ڤ�X�*R��}}��ݛ���Ev�Ʃ�%l�5:1$����/�τ��T��S��O���H��.E�o�0�&x��=�)�{�\���>N#y��/oV�6�s�Nd��r��f�K�˿�N����-��z���8��8Gn�l����L��%4c�,X��zb����7�̧�1HTG(�)H�|T��7� 8V9>��H�P{�UNy���M���m�`�F��h9�«y&'� ���I����'��(>�˴A~�Z`o0�����(WqP�)Qc�����A���X����V���@^x�����Z�����W��l�i�<1�tҪ�#��ԗM��Uİ�s�Q��L��֋l=fȵ�_Ѯ��������Edԥ��xJ��2��9�zC����bC���v5��-�ʛ߿�P'���.�#V-"B�S��8WҼtgb���D�@#�E�J��ŦG� ��%��-C4���L��`��%%"�5N�M	��eR#u��k����UhoY�Tu6�xVq�.f��A��'p��#�"�B���PڄT�2�m&Df2f�B-*̘V��h6��]"��秡
�z�xg�����1�� v�>.%�f2��I��\�/�[B7A�Έ�R���t�~���I��n I�TT����{	U6���D�\��Cj�B�~)��^���F�w��F�գ��	}g�m]j��ŭyi7���ߗ�O�T�wi�J�4& ;������0��$��xoc `t�1^�Bc�x�9�ަ-77' ��ʂI�c4	��s`/e��f!hA�6�[���9��Y��/��R��YO�I�<�4�K��R�^S�ʲL�O�QqXO<����DV�R�˖Z�>1!��B�Nx�[�q)�a|5�mL>�Ks!#F몝�H�-����;I|�'�Qn-:O0��i4V����|�NuGg�S/Drg׉��a}�,6e$�dH�=T�p���=�_MU��c�"̉d�_s�|����S�O[�)N�j,��u�|-���b�@��R�[֦�{�f��[��(!{L�.�{������'�؋�@��ޠ�����܀�!�_1�ia�?��O�3QVuV8��7�	��7��d�"9�[k^���U��])T���~no.)f,"�zDe���1�g�n�@���T����,�A�j�������L4rTyDIT��F|{t�O�&�\rI�1�)+֑�V��"͠�H^k�hW���P��s#�4p_^&�;9(N���<w�~�mw���D|�
�aFa&����E:��T�D U��J���q�WRݓ9����μ�#�%z��T`K@ �e�t��#}ǽN�M~�$�T#�@�5@�o��{]���x:
��P~��K�����x�M{�bh�	�JVn:Ya����^ݡ�b{qB�R!I\5VT���:hsWʌA8k�	��^N|�@�@�C Eݕ�*NL���[j& ;�mm��W~�G��R���%)~7'�by��9{���P[&�2��D�Vr^f�a��śZ���{������>QLr���;�t��T���.\a�S�E�q�,�!�;]�B�G��y����X
�Z�U|( Z Et~w� �ޞ��zj���dwI�L�����ѩȚ��ͩ}��#��֙�����aɖ������?���05Q]�ȒwS�SB���ξ�v��I���EzHY�Y��KiF����_�ȃ����N�&|Hd��k�r�������
و*�ǵ�1�R�&�¶hҤ�Y#:ii�")9��k!()�-�c-�lb�K~�؊G�y����֥�!�������Tx�ZZ��uw���d\���/���ld��B��Ly�+X�˟�a~�r���g�4���fh�`x�ڥf@��r	u�¨k}�8f��dn7�c2�瘺���b+��Uk��nZ/�����!?����!�U ��-X����+=n2����/#GN��^tX=-��)��b�.�f�"\)-�\Z���p�#�%rr;����@J7{������('ka�
.*7���بӊb����`ދ?��"!t1[��^��2��{u�C���1(/L�,N��-���=�9r��t~L����ٕ�NY����}z���P�i^s0I7�b��tt��D���~
����fa��v���wM��ǲ�q�\^ϟ����~��F7����o��
��H�h�LB>��7Y����1�2��A�1H�L;+��$;.�B�ۣ��4�O��ۤ+�8>3%�8/�8=ީ��~PH�b15c�#�{"iZu�:<+z�樻��l���9y};xs�t:��S�]h��n�3��:?�+�9m,����i�Ѐ�ՈU�M��1�h��a�T�ֱ�P��������)i��sK�fsx����%�����F�����V'5���Ev|HeR����q͢/)�)���s�B���*c���V��N�X�C�MY���m�A͘�-ex�4%?��J$��_i#�~�*ҋJ*�e�p-�t�1`*����7��"Ӱ)��ՊT�&��S�ٍ���!���?���ޖ�C�e�^�;x��L�esV 2Ե�q��Um�X�-���V����H �n(	��8��t2U��߽}Tr�auX����NBh4���}l
͡�֔7��"9��N�è����ܾ?Z�8M�G�:�݃Cz
FYȕ��n�9���W��ݡo�7Iyn��]@R2-�H����&�$_����H�S��/E1@"���̇� ����Gd[�³���4��o?v�����)�O�R�P���]�/��mw��`�.ח
5g�V$�s=���o
0�:>t�%�ĺC��Z,�	Eu�*>ɟ)�����
^��I��Q��b �E�X�?�"���f_��ab�.֪H���)�P\��yM�?�|����4��y���7ЯEj-N(���&M�e�r ����X!��s���gT�xG�$-e�48��~�i���h'�� 8��`z5��-i�!�5�\`O��=��8jRG�=�Т��w�1ND>���҆־;My�{�y�P��Ѧ`���� n�T����Ιl\,����z�������$ͧ;)�ҿEw9��qn/�ȉP�$�H�:y]�z�|1�#�ޙ�&$�ᱣ)��[`�k.�6�pY{�ľ\v+%�At�1c���d�6���L�}�`�Lp�y|><n��}��ʄ��5��b�8/�y[��": �I�۰�����I���߈'ׁP��N9��&pa!��D\�L+�כ�dW�aڼ�u�t��|3�t#e5J<۝#���}��J�/�Eq�Rx���>�j���v>i�B�&^~���%�k�������[b?�W��p��v7�@����(���������`�8͢���IU _'֣
�n���g��7_�t�5%��,��8j<�I�k���Z����v��Z�e���A�H�OB�#�֚�ߝ�������A�!��ǧ_��z�w�pd5o��e�_�O���-�����OlZ�0C���Es�W������ӂ^�d�����~�P���Y�}k�4rM!B h2����`pL>#�x@�TtzMAOSڨ8����G��1ؘ�L�R�W���Kd�:�޶k<�A��0�������^���7���\�<�J��/���v�%u�<ߔ��D�p���b�7ۋޡ?`	�&��~�΍��( <˭�_�Q����������Q�����@���}.!�`�	���h���Ȼ��rې�I���2�K���F  �M�??��8R��%�=U�;�ѕ�߶k�:o��7������ީ}8Y��W��,o��]�Zn��F�����n�.�����fJ�rAZ�,��	����,e�L%��b�D#:`�A���ұ���5��;����0{xi�^�Ҭ9V�Z�K����I�����6n���`�.R(�ث����U�=@��HCt�*Lk�6M�����x=�²�E>QL�M�T�	`�Fy�`�$\�
R{�kP�%���e�h�����X��~E.C,!U1{{�>�?��A��עzʞfYOH?WQ�Ct�|&7�V�UVe&�y ��*��Dl�s�ѓ�l@�uT�j�Zy�݈�}Нi��K�ҋ�yJ���7�����mP�+�1��P�v�'&�5�!25`;RHR��?r�!�qk�a^�RT�1����)��qa���g��c��~���`XF����5;2�!��A������ `���r{MkWS�g�Pr �D+C��_"P��W���u�%.�/0'+���T�g/PS��>T:�=��d޾�`�f�w��fh:�zFS�2Ԟlס��vz�6�u��͉0
L���Ģ�!�r�1$�peÞ$���ě�<<fEU�
C�Nbi,{�^�@�fG�
'�b���{�#|P��q2`���}z��>�O�,��"��z�/����*�l*���W���YtA2���~�o��?y���	j�C4�<n(a7���2�k<����K���e}@��Q�pN��snA���߲%�A)����> ��膂����fM\���B/v�sQV�k�l��`�]�^T6��砽�n[j�������\��G���/Vk�� ��rQ�w��{C|�����E>�s!���[+�1��d�����dLA_}/�c4�A�����a��:\Hړ��o��'� �w����"���8'�Y�oe��0ʛ��$\��O�����1��w��h��:hN1�W�`g����=s���.�����q��2��NH�snc'p'�@�i� �Yz��S�ߴ@=l(��ϐ�c'��!��TGz͏3dҩ�ʄ�-8�,����e]��J����N�����d�٩�u�s� } ����
	p���4\�kۜ��ƚ�������r�pz'>�L������ �	��ثQG�S�%_aK�0F�K\�@?���L:�fo�Ή/~����Ǣ��a^���u��bթ��iM���y|�QP+xT����R4����p�P���N��b���R0����n}���/�
|���l]O�3���q���g��1�/F���\���i��*���s7Rsp0N�~�RZ�2�9ǎ�$	�8�=_���8/W#���' @�
�	�ztA����W��$��7ܾ�Yy��}�0��2�ʙ���Op?����gE���_�l����9�n.��x�(�c�F1r'l?��
转���6��J �˪�*�0�?]uN -5�ϻ��<��]��8��9�;j�₤ǘ�C��]@[8&�yP����/���b[S�2#|�~o�O9�@ۀק0��?���E�k}¬#Qq��R1bF�K�r�$�S�,ơ4�4���`�oXu�1q	��<Lh՟6�!O�&�Q��}%=����$�Sk�M���m�]d{��<�y8���y����c{�>�|()agk�(~
D������z.���A���Yv����H�q�������j�Ѽ��=(S���Z�]A�-H�+0�5~_<S�JR�6�yST2��h�����t��8���3_�_�Z�FD
w�u�7�^`Υ����g@/�\b�"��s$N�Hh�+�&&Z�R��>W:��vr�36�K�(�w��}Y��$g������b���pW�ׅ�@]=���l���e_��)��|hA'3y9q�Bc-����*)z4�r����bƴ=[e��ťS����2-��8L�q�6��M�,2�9T�j�*'w���t�0��?I��i�N�S�Cv�?|�1{Hy�
��'�p��x�?k�_˙ŵ��/��\>����g�Fրg��SUC3zV�f��Sm�I!�/*Y}����Sfw��5kE��������Dux�NUp��t����r��ۥ��H�ȭ����R��k�m�����d׌��y{�V.e�HҀ�g�M����}V� ��Q����qw� ��ũ�^d��a����
h�p�1W3:1�@���LRpur���t�.4f�?Ɯ�[������~y�>9|	dt.�{��Hޅ��M)�E\�x�y��%-o�LD����:���ٶu��B|O�9yP#��r(U0�irx�R�c��Cq������ęcF�!#�7����U����p,k㜔04�YT��^��ɛ��Rn��;l�9$���fPy^=L`ԋt���$�a���V�=;*�xV�M<3����/hg#���4{�3*��Qئ�a��q&�E��@gD�̜��/���F%*��$�iM�>G���y+I�����u��Uō���E�{`���l��qV��?�)�Nl�L�J,S�|�QfU���9�zp<�\;ь�����
�$�@�Ń�1v���
�6��W�s�˵$��_�4�)t�N ��1:��
Д&%�(�a^�dA�|ï�7}ͧy ����]@�ƈ�\"Ҧ��}nm����r�(���s�>� `!a�4�C��.�#犑�����	��:�bG���Eb>����t��o/7O�󪂕�H���>�����"~?.����в���u���s��v�M�`��b�I���w�_)\S�v�)�_�#�w�!.�����,��5b���\%�B7�f�4 �A5!���{��(Mn������ɤ]���U����)����؆�*��)�$�~���kz[jO���z�5�sy���t1~��pά�-5��%/��agP�E�ui��0c&�g��O��\i�c�jeZ�e�Ra��(��6w���絪����ʙ�'���?[�j��d�pM�?vН�BH�ԛ��ϛ��+�d��R�ĺ���xV\�_�P˿U�g¯�w=��HYpY/Ɠ"y��J� ��\1��M�iҾ5�V�nYܬ� �2��ň��Km��z���d��n#
kp��I�Tw={�:���J��
��r��Nr���yLGD��e$-��K��3PR�Dn"�Mh��&';���r��s�#�S�ɗ_B���Y����	(8���>!K�"��̵�`�ˣ��v)��cy1/��Z�f�I�(���Td������Sx�Դ��6��������8Su?Lj`&�3�c�_����1୬h z�8����q|R�a�C:r�2L�g�;	��Du�U["�U��g 	#�W�~�(q8���n0�i.Y8J����F�Y��@�k��7O+%��sME������x�1��`A�T�HY-���Ixx��E���eT��e�Ml�](�K93��2��bќ�JMkD�^>:��j�	�-�/��� ��3%���(��)U=nf���⍘v?�kKѹ���0��z��͢�� (�N��ʬ�,��.$�W���������]5��z�E"�S��{�iR�@a�[^��%Q0�l����ѝ8��~(���.�e5R����7�t�f1��������RH��:�z�2�u!���k��%��UQ����Ϧ�3"��G������I��f� �K�>du���ɞ:bld���Zݓ�e =�5��*�^��F%9�Ͼ.' z�(�O�4}	&�Kf��
�xt�ê_�Tm-�5��݉���?�Ǩ��הu�C�F��R�x-��7_V�h���rm�g�:�G,d�EU!ᦿV��+����3�����pB[�zf��u�+�r�D��ߙFBƓ%(dO�C�t�~���q��P���u��|�2�z�� �i/����F��)?��^~��D &��7a���jo��QwW�磠_3Dz�?;�S�Z����HT䈥��� J�u��`���$=���׼��7�_V�R쏞�v���sb;e��g"E-U�8|{�f�c�����"^.��i6%z���7�Z6�y�j�O�0�b�a����1TqC9z��@�xH�&���5]TH�4O��m��Tf�l'q@��#�W�½�>��8s�����#���]\�f���vw��������-�uI�9�r��d����)�.��\��9AE π�J�lf��*h,�T>��P��-��C#,���\��dO�ʯ�7�A�͘��m�7C��9�;��P�ZFpw�}م1�Ko���"Ϣ�#�#=��o�x�\x�iN�uoF�A�P6��I�Uʻ�R���//�&��󱲍��K��&�>�(
��5ߢ>1�/���K�F�M�W֣ճi�4RD�2�~$�jL��2�`Scq���$Y��Rш�v��H"��/^5{��3���i�5�k��I��+󹵵��L�F� ��-_!#�6L3
'��t���̾�-
��V#�Qp�>�i3�a;�$��h����_t��o^a��x�_3�8G�����<h�~ �Д$!w����L��5�=ut{�X-�_E?!}G��}��H\�g�y�p�'���M��!��&Ye0H �ʔ���θX�o#��������BaUJ)��3�Z�
l#t�G�GE�Yd|$W�p\�xL>}|�3�>�F9��`m�T��x�F��hv+����"4w�g��I�}�(/��G?��!\ ഛ�����y��W����3ݔf�>�1[HԚA�(�����<�?�]a ��V��ʯa]E���e����G�R���YU���-��+A���7����h�;y����~�W�7��'��A� #s���+�����N
МOe�se�w�XPJ��i��-�Hq+ZD�~(�x��HJv7�Z%@���ts�xb,�.�9�n�d�A�6_�AM�9�a���2�+a���I9���h�B]�6�:�%s^���P�p X`P�&i�x�3�j$�aS�f��}����A�W�ő[�&s�"�"T�j[�Uc!�_��ǵ�/EVe|�߼9D{��`e��J��=�z�3�6���������f�2M����,��VW�Q�S�])�"2�&����44=s<NH�&u��8g5���U1C�n
sE@���D��AV�)(������x���Y���X'��x������4�,���7�t����P =O���_�C�X��ņ�� �NWF�����)����׽��/�}�&R[�Tz�����L(^s��f��f z�h�CT�Hֳ 4�zI�g�����&��Q#�A�����/�o|�!Aw��N�T����j�fp�:���������n��#I��E�� N-)vE�����k¸�,\���!#�'%8tD7D�/�畓W޲�W�E��K���f�&ᯣT(1a�.�BDUQ�oNыz�׊����6����t���q��Ox�A�Y��8{��� �d�K+��1d�^��U!כm�@�	Un�T�u� &���chcF�����	0n"�d�I[^P���%Nn���	�/���Y6�qϏ�W�O�#�����6i�D�*�P�\་n6;��<�o�?D2���,-����{A�Q8�V�{Y��[Bo��Bt�o�k�~�޻�S9ZNWٲ�μ<E�H�-�#���'���#�﻽dY�܉��]h�|��d�h�4B�����&�B�U��R���Ӻ���<�ַٝ�M4��}�P����H˰�!��;��9�Y����s巎Vj����DPQ�(5���k��$^�]�H�ܖ}�ɣ1�@єi4��܃�o�;L�e�Ε-�ɼ5.��΋��W�
��]�����p3ܡ��In�-R��8��:�%Dn���ҳ.�s/��sr��af�hM�0|��jec�+l��he�����j=-���y,�u�,��$#�V���	ڔ��*�9��K?�Ղ�6�`��Q���s��*3UU���2�Iq*T�� G�~Q����|����D���%ZT��O���}l��#�Q�:������@���H+$5�2\������s�Q��o' "���_Ó�
Ϡ�W�I��D�a���sZ�����y�d2Z��+ �����tK���Ӧ�?Ƚ��%-��ʐ��Sj�P���2/����?��*s�Z�g���z1�������=�����,Bv��,a^>��AY��@'&�q(UD�L,"���|�V���bi� �m���#+�m��3�X�2��=�e3�Y~�&a"=�Z����������Ut�a���+;��%̲7G�޳�n���&Q�^�&j>]zf�W�n�����R3WD�rn�@4�lA�	c3�&q���1�D�I	S~�Bx�<���gY	iS�}4y�2Lj�ߋr��wm���塧W��CV��O._��S�"�Kxq�?�K��b����?��P�$�A'��y���!C�Ί=F��3�2��٣��~��B�ˮd�M�M�4��X��/U|b��ԟV�Uv������R�]j�T𬰤]���TVcsD٘ ��b#�)Gd�uD諸.��by�1��J������>��~U �ǃӸ"{=z�3!~�FcL��H�H괗B�sr�M�� ߈W�$��I'6�I�h���"���N[e/}���1�$"Da�,): ��0�"�Ŋ�r�ヂ?:���Y�/u{�����2<=�d%v��p�H\Գ�Z��r����gD�v���RZ�.̓��[� ��sM�陥�����s?3f���tx�z`�0����W~ .�Iw\3��)[���[��1^��A�<�V�����:��֊ԏH�S<]���:��s3�13���o�CAw�'��p�9��'
ղ��C��_H��+��Z̳��g��ˊ�����Ѩ[�:�y��#��TΉxٻ�/�����>V׊�������-���,!�T)�2_,��4�Eӏ�~���Q3P��>�iavL��e�[��p߆|�]����9���	�3F�N�),-���
=�&5����ǃ#�Đpx���<��)�%6&<���&[��7`���6'�Il`��7����9�h�M��"Z�>��:/u���c��,��~!�P4Çe�E��G���MD��:�7�ߦ4n͌�Ra.���#�H|1��.��'u�Pֲ��,?��~8�糗��	������Q^��銌4�P�w43̵�͌J_���b$��� ���Qҹ�s��1'#�P%z�}�G��x�U��������p'���/Z[d.�MI�$�U~����¹5\ۥ�t))'��,��u���4�@E�#���N��¦;c(�>�f��c� WD�^��&w�P�m�	�q�1��@�7eP��KNjp�/��m�J��̒L�pf��>F�-P����{-��9;keQ����+p0�����I�"���Y�ry+&ѵ�,MY����~t�-�ʀP������r>��z��Ċ��91��>w����J?N�7%�s��.&�CH�w��2ؔH�,�Z�0��!t���gbiJ��o��\Y�,f^k�F���
��<r�9X�����Ýky!�l	�
I�dqT������Ov��;���6ѵ����G����7s(a�v�TE�<�?��
��M`��P�.$8 G'��=ҵ(S�1�J�-��V�� ������X�O�Yy��n��N���߫-=ʍ��URm£5G�~BGt��B"&���Y��E���$�0ҒN�w鎬� ���e�8��2�{"��[:Ё_w���Q"�=-:uDr��K|%�l�Y�:�@�qu��F������|t�ܤ�������L���X��&i���1@ʀ��S1
���Prr!J5OaǙ�1ћ���0<{�{����MƱ��~�x w�����G�n����>�ѣ(.���<k≫c	%1U>H��Y�A}*B���fB(3p�#�:�\�J����4`B�9��J.��)7�	�t�7&'Df6I��B&6?�W�e�2*U2�R�e1(��w˹�ɲ���4o����3(�W�ϭ[P��N���O-�ͪ�Z��4 ;��Q�yX��f��%�{+{d0Χχ���)�����(E�B���y�5��D�������!�U9�w,��3Nl|�_�:�6p�� �♠�IA�NE�	9�r�tʵ���r}�E����ԣa�E�f�(Θ�����;zJ��r�S�Q�	A���xĥyLX_r�ڭb����*4��ld(zJ���砦�z�+M����71��9I� �@�$\�I��/�d�Nͳ �v�i�Ӆ:G:$̴SU��`���[�s{�u{'���O��ϕl�Wk<�0�G�Rh��8#ˤ���6=
��Cp�J����y��ePqA6�'[k����v
�_��'n�u�)_>Nc���Rmd�P�#"C~��P�5�X�����ߖ'��9�Бr[��gcF#@�넼�l�m����贚��N� ����h�;D�ʧ����'��@�!������t�ZX��;$N:��`�1����7�4�9g-�A�	�u�^m*�%)��L�܊@[�S'���ŧ��3{��V�!��r��X����-�i�,{]��n8IH˛������J���ؐ�@p�$����Y�+h餌�hDh��������ט3�e0Ⱥ��1����b[FV��qk��t��{�}����D��
�5)5(�����&
��T���*�wC;�u�C��ٛ���w�5$
E54���l��Z,B�/ &D���x�h��ef�F��鴱rңN7�g�~[�:�( d d�v�'��x����6h��#��뺦k��%�
nX�~��Q�
�p��+j�d_�8�%M��c!qн��T�V�AW7��mq
P[W�|�"<�:�V��[�f&+5���������P�X�?�\f�wd4�w;�3	$χ�m3>�\�$|��6��%2� �)ܤ����#b�6M����j�<�.�{V\�
�2�|��@i�G��e��,�!�d�`���D�h����p��XU�*��sK�r~Q��X�˱���m�_L¦nI&�
��n�%nS�3�y�P�8����@���h|^��MX���
yǐa8���8'*m	(R,��EX;�e��u�G6AQp��23����4�|���_r?�t�Uq�ԝ2m�Xx��	��u�坞�;0\<
B6K�����(T�/Ӝx%޸���p
}�n6�Ā~���� ~�7��!�y�7���V��GLD�#�n�`��ra� �Ҫ<����Y9A��@���֋Cg��,�c�#3u�$�/&���p^��|���4���r�&e\;z�-��e��΃�`?�%^��H���j�/�a�oAZ�x��Xk�eB�.Z/���	(�x���[YEk�ف�����N&�������'�8���hv@�A��a��3Smd!I��k��}f�K�B#�Z���G���$�C}�!�᱗��{-/��\����#���!KՐ+M��s���SaЫI�
7=��*p���[�>l��Ls��C��R�E
o0b��]t�7̂��t��ę�$.�G#Zh��_j��O�]�S��#����[!��0<N��$��DKCg� �/]���e=��_�� ���g��[9��nW8���J�ړ`3j����N��</�+��qfI�X�FeFR��x���6�P��Iz�R�nM~+��5��ߧH��v�o�`Z�s���{��U��e�'�W�Q�r���i�GE<>դ�62I˾T9���W�Dz7J�̖�f�O�#��Fu�־4��%yr��C*�'H[�kf;��5�-��~Qz���]����;��v�?=u�^�V.��3�:t�P��Ҍ܀
�.���*v����|-��O3�o�R������XD�T�'�P?��˭�[
�ǥ���Uv�7�V�)�#�1��z0̓SO�oZ#!֙m�U0�2iR*9��ZwQ�AQ�+^I��D�QD��Z����~���bXT��I�Y~h+Ȩ��[��K i	5
�08 x�m��>��77K"�;t�Y�x�o���bh�
V�ŶJ|���d�>�;�iB���L����a�J�
@\�i����,��`�y��"<�:�#-�g�}�s]��{Nb��	_M�0��.|�D����Ū��9膵Vd#%�Y6�&^����?� ��� 
�yWn	2|��+;]�6�4p^Vb��(7-��pPsߓ^�F�z1�d����i�Z��R��}Y�9���[�,h�CT�T+	����ƴ v���M|��.,�R�];����;JÃz�hj�u��A�dm��9��7���Z`CO���yqZt�A1�0�+G�<v�j,������A��{g��
2�8:$P`�������7N�8+|7���V6.Ȏ�a>��.h��8�cQṁ���;�)�ogKL�G��ȷD�_z���_�/p*#� v,C@X��
[e��;���,�C�P�`�n5���S�ezwyc:H��V�E�gx|,�T�Rc�����̇�e�\4h���{�b��X��;��]�x+�(���;������{CUJT|����'�W�_�\E�\ϵ���o�2o!~�h�K3h�2?:��e*ʺ�La'�T�wOMA����S��7��c#�Y�Y&��5D�[��&?U�iR���8�D@�����d�`ޙ�����Sꆕ.�â1��W)T��Q�N~��1ϛ����]�AL���?����Vf�g�0�ߊ��PyQ�K������&��a�����+�[� /�.i�{���Vj��EG|�g8�%�2�^H��W��ΔuEҠfe�F�x@܆=``��Ϳ��K<�[R� G�B��ν	C� �@L�� �:��܇J�J�K;��*pr�ml��v�_�U��#e���ʈ"�v^��"��|HU��;���L��FL��)�ya l��i��}XX��Hx��5m����en���}���f�-�n�����DЫ�c�M]����7��'.N�kG8����}��x~�\:���hLϥb������ƙ�O���������.+�<x���XP&mv#"
�O���Z�>i��љng�5n+x�VG*����z�QG�č��_"���v�8�&��	����.����!d>"'��jP̴5�u�U3N�t�M���(��[-�Kו ]5�#�!�m6�q��צ� �k�aW:w�� ��ba�����f���[�iz����e6r�W�r]-��(�Y�dJ�q���w���$,u��yt�5]�v��ӱ��&Fǋ~3.�	::�ڰC��ѳ�#�1�i��TP�etvXcGE�� I�O�\>�	h�4՚J�&����̫�OV����\���ۣ]ȓ��;����	�p������<Qں����+��2�����ٍ��θU��~،l���h�-Qj��,(����5JS�C�D1�Q6���@���2��dF���}�ԇᶻ�9j�&m1Y믤�7旍�L�_��� ���>������^�M@̽C������Bd���7m�iwE�Y�}`��$iI"��"���+l��ζp@���?�/F��Ѷ�sI�t����f!�7|~���\7&PL��ɒ�]�o�N_Wb�j�)q����	�f�"v<a�DQ�Z��0&X@x��[��I�5���g�k��mO�1Z�N��l���j��u�Z!�C/�f]T�UYo�М���G6ɸV�g�]aB����J�#�})���$hAD�;#8����R=f|�LH?�=�!��e���铁yd������@b�/���Mf��r�Ό�by��~Z���]�.d�|w^Eq'w�2K�4S����@�w�\@˦(5f��~����N�8��϶�?\VL����L���L�>�d^ hl���>�"���J����䍴f}�ɰL@�ٖ�FA�R�o�at�SK|5#9���#�
8�%�����f#. �&����fq���ߪZ�y4񁀏���<]�LNhA	!$���M�*�*��4�L�����d/��~��S��IB(q�ݹӑO�沐�*��Va�P#�8�)k��G�x��+��Uq,��r&���
*���֛��{6�TU��:�^�>��h��)!U��y����X��U �G�+�	�4�`:ā�o���b"x��6� ��,�����e�u޻PF���E�a!���s2˯_��/`�d��9a8lxT�6�XǩOe9���W=�b��ɓz����5��D'P����]�i�Ї�����X�G�P��ݍ�a�&��Di�r~R����������a����b�w�D��
��,��f��%�L|���`�k*E�
�����@�����?"�o�� �\�����t�v��qb�Ow{ѷH���͊4M��7����w�<�Q6�*�h�`|�L�٬b��d<�a!�e�NةT�S~�1%�6c�,M1���wα d=�0���&�.���{��(O�!���h�-�Jܜ������T�Ya��/��&f�a�~<��}�L�M��?b�ŴUsd���1�'�����3I���ݰ=�ܓ����\S���ճ��-�6m�%P7�Ã|}���J�Udj塕<h�qB����S^W�t���Z�-�`�����B����s��e�7�<p��`������o��"�1�P�s�sB"�@���E��^ʈ�@͙�3�US�Vb���l��� *y?�-Rp;�T�$�f�S 
[�)Z%�VAA�C
���<M��Ч�Nwϭ��.���!V�W����ʠ脿���k�����{�N�S
���j(�,�>�@����M�;`L85氽w:�|�tk�B�\��� �ҭ��eV����cS$� {JrS{�/x*ɰl���A���k	�Umc63L���JVՊ/�0����U�����ז���#����0K�9ui�5Y���nYc�\�F�=ѥ�S��ŪIBS�I�%f��7���ܹ��Ʈ-������KP:Ɠ�kC��*g$#���UDC����TlZ�.���n��!��	�Am�\R�S�@|ψp��t֩�+����D��&����Ha�#�B.9d)��IҭSv�P"���]����vU���1��a�B�8�瑄2�� G��d���~T4v��E�)� D�P
b0od+�i�R�jZ�}g`��
��Kjhh��W��`�a��gA??�ٺ����*�۶t��S��8�c�i�B�Y�JYH��&���]��ځ3�\G���bR݈�a��o��\ X`U���T��~k�{��(0ߙ#�,_�Q,�$��r��]~<]����8����s�3���XxEߵ� v�w���J�3�����Yo��3�@⛎dŕb��%t�2|y��{���3�������>�TR(������u@+@�S���F�!1�#�M��=\Q#W�����W@ `LWh�XYq�Rp��+��zld4WG҈0[�~�gN��v�̀��
LM�w��v�)gn���_�	8�ˠ�f-���և7�q|V>��W9*K��gpj9�����X�x���'78�V430�Q��)��<U4�@o�4���&�V�34W��.�)r�����/^Y�v5���5c��
O�%�p�.~��&(��$f��B�l��`;�ݧg��}�a�>���*؂���\w�5�5�jM���IT��d��䝴g�b��H�АO�����F̢JS>�+^�[���1=�¤����n��5)i: X=:s�}��R�#��QL5-{g�߷F����=D�}
��f���F=�B�K�h�$Q�u��7��5�/R:�X`�)!�T��,*9�W��i�x������֤�c#������T��E��'��Џ�w��O�f��b�pt=Dwa�TR��]>����+3�'%�B�:����YuL'����3�ƿ�����]h��8: ��[�\w���M������?�曮q��CQLΆ�	q�$�?�AR� o�4{vm��Cs}���>*�j�l��z=G��(���7e�!(|�W<i�wq�NY�X��+���BÙ��Ѻ���֞%�WU�%oש}�W�b��h ��P+�#u맕�^y��BO�$��eT׺Z�(U���p���kmGȸ� ���)�����.�5��hr�7��}��f�6�^��XZ��bl��'=�]�P���>�9ˏ�O b�W�<I
r�5��/��9����,�K,2f�l|�����*#��1�R+�&�n=���Ģ�<۰�VІ07a͖�����w�j���aJeF&4��T���G,�[���깺n)� 瘻Z.tͮ�Ew%L=���.;�F����2��L�[('U�qN����un ���z��c���O��Y4qJx�OKg�:���+~K�<W��*��\�Yp����>��. X�&�E�AФ&������U}��!��h1$�b��&��`u>
��b﷮�µ�2 b��N������/.� ?'��Ȃߣx�>H� �l�6Z��kiB����n7(�1*$]c��6��}� �����i��|�1���FY�2/]b��u�bW��-�X�\���)�U�s�w^��n�v�eQ?�P-����{����O"n�Z��0r��뷰
��}�8��}�Ç�`I�]�$��Q��y�4��7s�����1r�:ų��������N7g�� ,,M�*�Ќ��xM��C�{<!:Z�PqMB-*ڧG���}�b��p5�ev<��$q�\��S�м�cF��\�B\F�Jc(�ҏ[`�mK�	:��N�9�4XЧ&�z�b�J����M��M�<Ś`�d��\>8=z�&���E�9�S����Y��H@�������
���d��j���x���)���M�R,	���j:��j+z�Q棃�6I�S�(�&)�GbS�/Ry�kI�N� >D.�Wݸm}���M��&�����]/����3>>9;���&L��m��_b/ʇ��r�B��7����c�
7e൙9?4�OF�	��Q���*�,3����͑jXy~�x7V*��F�^0�JπY�����XO�S�K5sߙ;W���R3V?�)J?L��4=���IV��(N�Ϫj�iΥ��9��T�K]ȥ�=�;�(�����e���`��g�����w:�1w�.��K�������wf�\9t��Kw%v6U�h�m�˛��*|6���0d�׷�� ��R+��@���h�E�L;�?�����m��|B��4��;��̏����'�g�n�8!����c��L��?�xbD�2���uZ�x�8��u�uƣ���^-9������E����A;����33�>=K]\G�ˌ��͋U�(� I�	��Y-�ŵ�£*�C����k|������v`�5��F&�p�?�J�P�+�����yF��I6�̻ o��L�7����-_�y���kQe8<�&xu���=��"61�p5Y�C��W�X��cF�!��CdU��H�����3���-��� �:���֋ɫ,I{��'ܯ��R�"�"f�xT�C�J�̋f���#����eiW
��������-�0fx�$��0����Q�o�K�s;�+����V	�ۓ��[2<�"$��G_���RL�@I]��Y�m���t����B�UȻ3����
�XX1/��AZ�׺<�_��9x�x��<�i�����uI��s��v�Y9{*hG@o�&��$  xe��e�>��A\S�ͧ!mw��QY����p&�b����ridyjA�o�N�/n��w��5�\�x��GN��x��A�����J�l����w�;Wڂ������WA���KL����0P�0�1�hu��Iv(%7'��&��^(���]�h�cR���C�k#�4�D`]��q15�].������nM��̜�+�ݿ�6wX:���p=�qv����%0�%]��r���܁�����2]���fd&���@v�^� �R�L_�E�s�"�U>3^�G��
����il���x���,��R���_��6��)��}T�rַS]����YIP`5���$y�Zg��&Ҥ�-�C��28H�ɕE%c_q���6��$<]e�t�W�@ϛ��[$an����ɤ!E~p�5#�D睩?#U�����JK'��s.B�}�q�b?�ފ�%vw_���8!s����䁲�uTG�\��b��L��k�u��1h�&�e��S�5�v?�Z¬���.~kc(�
���ڑ��ݣA�]��d�OV> ;.���|���/-u-��G" a\C'B��c�Oc�����
@�1�P^+�5���B���d}��(?�����~1�.l���5�
�=3I���9L�!!�"�0��$��DĴ�\m�ɱ�Q
��+7"d�x$`����� O��8A�2�צ#4`�;/�#�9Y)^Hڍ�l3������m����"f^Ɲ��Q8��IrZ�{{��.�9�=N��R����h���bO`�{���~�Rꜚ��_�S��))�E��{�fq��TP9FD�-B�@3�?o�M:��S���玏n�a�����.�z�G]ɀ��-h2⭍c�������x$F��<�.�<��Q�~j@C�oU�j��������AG#���e���N\�PƉc�J�;ʪ�@c�Πh����(�)h�����f��a�UJ�zEjmg��cj��*�D�U:E�]9z�ӖC���$���H����Z�Q�}�0�n�e�֑$+�u�^Cz��Y��w�v��J��O谧B�~$C\(}�[+�l�(��/��/Z��*J��B�]eX��l�8ߊTm�����VW5I7Q�L'�*�7��ۜT��Q��9%@:��Ì��9Qm�8W�~t���n/����hC���XL�d��|�e� �S�H9�����T�N(��E1������@b�0_����#xl�܉S�+}8Ӳ0RS��[,��ھ�=e�'t]�F�!9�B?���F�^�A���Ke�굋
��Q�б?bd
:�8��t��#C�����~We��B�����?�VSlnr����]�ʎ=빙�^���V�ܗ���M�P���R�����B���z��^�ǩ9}�d	_/�Qc*$$n����L\�������<���`�Ih����/��o�.".p�T��e����;3v��ܗ��4n�)@��b�(6����~�ɋ�0]/ClиyL>M��I�e���������,��Wo�FzU3�1�u1�MY�5���[ڸ����ǘ�2kL`A��q�G�fm�����p�GW��]�5�S^l�x�~��k��+����)���O���3p��[~��r�J�I��G�)sg<��vW=b[����hAR�|�S�E�������{��g�r�ӈ�"���5�!^���Rn>/�u���t�g$��Jt@GA��F,�(���6�ku���л�&RS� �P�Ж�x�z8z��ң+z��ҊkA��BE�o�/\T��r�F�&t^����H�M��(�ٹQU�WJm+,B���^{�@�l3�ؑ����v��YA���e
+ʀ��ct��M����d����;n��d_��=,+>s�-��X�S��uO?�NW��j��y�R%nx�wE�����n6��~ؼE济��<�7�Ҕ�e���
{�5�g!j V;�pO�=�c#��-�g���"���1FEy��Z}���m�z��DRwĿ�X�'�\&�*Vu]Z�6��w�)�Һ�[��H�t=�Z���9�QQp]kJb�����ڠ��+c������>�9��
:U�[�,��OXF	��e'?OI#�3�^7Ι������S��C��P��v�����?ko\O��S}b��Ɔ�M�}��B�ť�>��t�BQO�>6�8��,�\��M�
�#fKt�`������r���sp�.��nPX��Y�5�, r���{>�P� �N�
�,o�_�u�I���Tf= d���iie�d���'^0J���E��I���#.���p��>=�n�\-����D;����-�\��,����� �VV�uce��zICvmL�����&��W�A$�$�d�}gĊ�����x�o3`�x���y
��Xぬs��؟is��.^ �i
���bY�X�����Ev J�`���R��}��{�bj6+�����͜e���͕�b=Y����"�����͌�wZWKF�T�4PA�"�ғ-𤐻���boi�<f~��g��~#u�wN|�j��'@Pk=�%�"Y���WUV;_-4���<�`0� 		�uަE=!��F �Q��c�t�����(I��	�]k�#S��/>��K���\J��4�񯪉K���;�AI��LN%q0��܍*>D��)%�ϰ0�QP�?r�ø�={WNvx�%M�����#2�~�ȮV��\Z�U$Շ�3C�7�j�\&�G5�>��A���SC�y��Z(�h%C�ޟew�]"'��nI�e��,�i+-��zN}nl1���ys��'E:9�H�2@�o�9�V�.e*-V�?xh១�(l����u8�_S@�[$-���K[��6��ð����)lS#x�\��z���2��5����JN�v6YW�%cT��{���
�� ���!6�u�[���^s�x��ї�6-���[�<��<��a�b��,@8i����)����;j�bϼF&Ң�:�~2J����#R�����f�q��s3B��\  �.���f�\[�tU_-�.s_�Q�i�J�.l����7��Ҋ^�-��n��X4��l+1�������xĘ�z�)Ύfy������F�'�dcz�J���TG�`�g�q�ou٧h��]�p�ͭX�th��39��&�\��H~I�U6�X���7|쑙S��O�1���ZO�Z�^d����,�;plD&���Tb�E�"�p�3����K�MK�l� tez~���:�k?�$ �F���ER�F]��V'�,.��[�*V=Nv/|�(�c��B���a�,°�V�ۭ[1*NE:
쇄1�+��8K���c=��+��x^��rvuw�A�Gb�厼T廼�ϺWO�t
��e����z�*�?N���Ŵa���D�+�w:7�n��<���&UQ��ė�E��N;q���+o�J�7"�u]�_x9ck�ң������1�����Rv���͂�&��؈��s���;Cֳh�/y��(B�D�['��#tĨ5��I��!���ƧyԖ����7�����{�P�kk��.&�YO8��i��d�CQ#���Y���h:�k�=ȫli�mp�W��f �	c KS�ev�~��˞�Hh�FZe<�7���MAz��S0�;녂> ��}�%�<�p�[���`;��y���6���;���yc�L/���S�y���D�p`����N����Mi&��CT2+t�=,��m4�u.HK�& E񱘪���j��j�b��^��������)�)�M�M/�BԟT l2����)��|��G0�t�����j��P�`Wr|�I�'�k<�=�Z�B�2�^��`}{.����f���ǙxG����/�:��x0�& R��ȇ3C�	�W@)dyk0i�SI� ���S�?g�&�s����9GV�p-�wψ�P�}�i�w����USF�R�����T�I"}kk*����Bt�ɈfX9����2$�]�p)�R!C���+C7/Q�#�%A$_-�����(+�(�����}�x�e:]D#`L��]P��\p�� K���q�e��+%�5��8�^�=a�f(�X�&�q�p�-|s(�x�M�HnxV�|�iZ���*�R������k�-����r�����6Kw�3���L鶄�ُ&Z����O�s��W }w[%˔���'r�iYӲ��_t�t54&�$�\UݝH���R�ǧ�(d*��A7�Hn���4��<�Ù�(�Yw y���f�����a[8)����l��Tw����/{Ud��!���+ a�������l�2Z�����Cq	"΍�����c�T�"k>�aL���p^�5z�����10�;o/�l�V�����.~"�h��d�F�����H�F�>��x��a����+�yYNݰ#�Ed~����f���1�a���I�u�q4^�M� Fԩ�v�$gN�s+��ǹ�Gy�dl�+�&Dˏ��x/���2�'�I���gAOK��ϛ��I��b!0�G�)��������G()�'�1t�G^-�{�<�f��� �
�P��J׉�a�����N��xq�q��,|4H(^`�ހ���܍9��z(�\_x'ILT��,\��yrA'�����g>_���w���մ֨���1��7irb��ak��v�rN����ʔx�#�n� L|��>���m`�8`��A�7@�cR -�������\<u8�&�| �?AQ�Z�*4o��
Q*�M�,�jr�/j+��T��\�+�t
5�wPw��cSq@���90D2N�����B�Wb��&�Fr����������k衞�M���D�B]s�<�ȝ��nJJH�(�L2��Q7���0����os�V�vWp<;�8p��h3�\J��/�n&G�i��=gkܡ]~�j f!�Vdoˆ]\��4��p��)yJ�*�X�WDc$�C����c��Ue���i���`2�;�.�)d���訏-r͓0��^�\B��L��C�E�}F��iP������F/�2XR߀6/F�̵\x%c�����3�x3�w��r�aq���	���qm�-;�$�O�@����ҿ�"]�伱}��U�����ߋߦ-߈�����R" {g� zF��� �I �c�UtK��؋;V�r�R��li�I脭_w�@�OݸQvqW��~O%p��x��<
HYIB
&�e\S�����w�`l�������|�ov��8���($��"���8$����C�IB{�Ð^֫h�M����8��MO�\z�A�uE�¢��;��u{($��T�p��n���,����.�vj���<}g��m�SUqI��i�'�B6\�xd'�W����8:'V��|@��l���0#M�Os��ڨ�%3�8�BL�>�{Tsb�v6:�l��&:�Cת����ݗ,�����cI��$�;Cp܄�#L�����+Ӻ��������fD�`j� ����-(��c�igF{�?�R/׸	�m�~4��F��:��^'��b�e�|ə��s�/^6b�>Y����48�m+���-6-��ů�;�鞜B��b�mQ�/.?]�&(\�X��;�!�3:վ�m�����n�N(��׏��<Ғ��>`�C�{T�Xmn	���AbޗΣ�:�Ƕ��j��Ax��.g��Y
#�ߎ+���p8�0r��و��\	���E���o)�Ri�@��R�Z�S]tN��ll�,I8��-�v�8M��n��'}�T�#Kc�jb���&墨*� ���h�'Vj�L�p�M�B��u9�}u��={4��>�w68 o�Rr`��6o���\�̴��õ[����$U������������!�A�]���E�����>o���_�$�����Ӯ��J>������2����2H�����^^�ٯ��d�by?`���r�g�Q�̈:	�o���zT���T<r�� � ��x^�$*���c����Lq�+Mj�UJ6�����_��p1���M�$�(�x����ݲY�Gi�p@���奄R<ރ�d�z��a(9yw������+O��J�Y<QXU��s*[�-��a�m�ۊ8�<��*�"E&`�{�~�\.b�Xn���LP�.n�������]�����vXdȿh��RW��"� rI���*`w��o��D�z��f��?�QP���p��cj�Y�ť3��NB߰UTID�L"�Wβ����_���Z�V�+s���4�\J/r�E=���y��ܝdt�*��k�����2`e飽���hJUq��%M�7R�`c�.�����OE�w�6����cZ�b���������� ���*ׁf��^$��e�zs���<�R����abq`�3�t���R�e�&�	���{�Q��>WO�2룤�E��b�����C���T``09\EV���h��&N��ϑF��
���_>P������t.��L�NP�x�/e,Ě�/�4�B��e����}���/�ImH�vg�j�Qws���
����1�.���=tұ��ɾ�".�ؿ�����β��!�]S���4����H���^����/Yh���`�7��og��$�)m���|@3O��?y����H|�yN�[��uٌ������5ҍ*8��'�ft ����krբ(:>V{�f��(df+%sZ.����b
�:�齦Aߢ�.�jUe~ʪ���F�0ӣ�9�q{*4LE�.�C�?�q��h��!��G<-:B�,�yM*���������Gh�y)�A`�*l�w�R&����S��US�+Э���bX�ЈE2�aQ�� �����ρ��lQ1z�%�3СMz�6��p����+=��� }���T�,�/�d��_4���^���s���lfB��t�{4ꕽ�~�ֺ$�ϝ�M����w�lA'�u�qM3�X�m����I>���MI�QL؆�
�v�S;��kK(��v������#��r�B'F[�v�0�f�i�y�}�,���D�Rz�î�*�UN��1!�	�"�d��@�1�������}��:�F�ZN0�xAF��Y��bf�2�W"f���X��������k�&�n �c�#��]����>ۘF>�0�&�jU��!w4;P:��i�p���\T��3�1��U�n��0 �P�m^��I鹹@��G~�F�!��6s�J_*&)�L����~���7�)|*O��C`Ť]�j���>����&b����}� �j�N=a)'.Ҳ��W�'�۹�L��̵�s�=�?���2+܀G���`�UDY�Kz]�'RF)��y��ZhY ����R`�{.�҂j�V�>��B�����+/f�m�mkPk�]7�P�3J���)�7���3	sm�	��m-"�Cp��%�f|n���~鐅��"��?�ܳ}P�5\�%{�~A�Bl��z�����z-3����ۇ�D�y䁓0�ǃ��K@`&W�S^��4[r��UGHK�Q�	�V_r+8�K�9�cr��N�;�ų��A���?A͂�U�� �r���a��� �Ε�^��%Ա�D�7ݬ;17z��8|�Nsl�(�(\�y8��\*��	�Rw�K|DP���y[�|��2��L9؜��`o�m��\"��Z�9̪����$I�n{6���&*��"��C���@�'�8a���	p�Nx=�g���@���.R	�	�;Ξ��TI�7�H|wwd��yx���:���6cBB��N��ɯ	 O�/}C��}���������ݖj��Q�/�/o�R�]�)P��t�:���.ʮ�~Ҫ֐'�����N҇*�:-wb����O|��H���P��!P�*n`!���'& �C��5 �Xr�8�0�(+��((���<���
�qx(�
�3�^�\]8Mھq�dY�4�HS�aF2�!5EU2���nً5"C1K^�5	~���mi���9Z2���T:%4V��v�m��X�-v0��� {0S �>��WDG��!���O=�% �f�&n�td�a��pOK�ز1l&~A�nZ�`��t�b����#�Kt�W��7+�B�����5J�=�i�ܕ�W��+�=�.x��Ǩt��6E`��v:Cw��Fa�W���z�Tp�����_��QR�G�F镑.��H���`}��O/����|�
,]�V/��z͂
W|���D�e-�Pz�bF�QgU'M�A\-痏4"�/�O����xS����q�Q�������Lӄʳz�C`���'�W�Z������K����C���{[���C�e��lf[h�4�[tt�1ɍ�������Z�
c�y-�Rg����	ʒ狢#zYE��6�V����C.f��D��(�;�����n�O�������D[(��bT�US�}�%VEv�Q�j}>
�|/:��X����(���wEhΥ*�\�_{�6�ʞ�b��g�ϱ`���
|<�g۽MZ�T�����P��z������~	���J�����=1]�q%8��]%�����X8G��W�H��:R�_�q���Ku9�`_�?���{0ŷ���eq=����>���H	�8�h޷�Ol��y�P��ص��*�49g+M���q&�!*	�M��M�>�4)Zq�	�q��Y"�;2K�A-W`Rd��M��}��8���y��SavjVȂ��VF���]�` ��'���(���C�aR���c�i����C4jAA=l�& �ړ�Hh���'5�5�V/$�zTH<E���1�Z�?4�u��!�[�OW��#�3�U�Q��`��H����*wS�\˓o���A=��zƦ����_���1�Mk�R(:^��*�w>x{���t�����[A:�w��b�v3FT���Ķ9t��)0�޲n{�tc������9rjl���(�=��W��Ę.D����8S������&"�[��J�'�Q�:���e�,��@R�q��P���JmB��c�����
��߶��傐�t���ز�|�P�zkHy��<g��iuznc���꫕"|���R�M���J��6���/��r��1����2@ԅF�Wѫv7���;�Zr�+��Y�S$��v%�sj�գw��3瓀�3Ul�#�Z����(�a$�"*r���B�K�ӼY��0��GJ��>������_��|������D���
��A�D����2���i�5�BX��߱5ov�B	����?xf_�ĩ#�9�����/Q=��X9��_�O���7P2����hъ�3��T��vI9nG��##�����-oA��|�(��HM=6�J�r TA2g��rh��G8�@�~�ǢEV�Ij�}P��۠�zqjj|Q�V���d\2�b�{6e+����h����������d�!Nk��@iڗ����r�)� *�m �2V��DF~�^�U��`�-~Q
k����A�E�fLR�+4�!MX-�9�4H�pzk��e�U���	�����*3��Vd��U�&�VB�$�GD�����t���rr�
0U�GLj��p_�}NQ�����{�h��[����v�����+�I�(�Z�><�;�]}��Y��Tz�r��Ȱe�c�05��}?9��Ld$�{L 0�D��?(,��v�W4֧n<����I!�R�d,����� :�E����[Pu�+���hF�xɭ���v*� ���ʽH�Q�-�}L��r-<�dJľK��\e�ͅ�1R�&��O�l�[L��tk��(<��ל#wD��h��q���$#�lj�������գ����߰�6�k�G}�;K��������b�3k>6o�C�*֞�~��ȍ���P#/{�N��>�,����xED��E��n��������hb1�1���Yc+'�e]	%�OƔzr�&�w4.�^���P�)v����z/*�pͬ��G�����HБ�>\��;����
S5�q�Z �K���u,��"M$f�=���.��7V|q9���7_���d��G�-�(ރ�As4�Y�~B̚f���PYfX X*L5v��wD��%��Lq����X��v}$%�����M���/���9f����cl�#Q�6RbSgm1C�g�]N�_$'��<#�{��qm���5�i͢�}�y���V�,����X�V;��ZQ�~�ke�Q5cByA}pF���lC�l6���	 �n��݈?��/��+rV4��q%��{����}5�����;]��
M�Oۮ;����cI}��\���%��Ê ��ߢ��!��U���@$@jo�`ϥWLZ����q'�9�W���`,��<7��~��L	�$ӵ���h�|�>eFA��y}�G@��7�(�AЧ�rm��bs�v��8�[T��ڼ����l΁�4��+y�u�$g 5�z�'S�U��~�c�f�qq!�~V�5,�Z�1`��sU����^����^�;,]d�\M@��ܛ�@��l��/TY��By�(�t뙣*�!���
�v�?wʰ^ ����nP��P�]�#QF�����fP���o�قz<�����D�����q����%�u��h{q��׿���29W��'�y��֨R��ll8 ���c]��w�r6Gh�=�Ep�u(V" �C f�����B�]�����X岝�#j���O�,�oס�D;�W��m*W��eaw�'�y�>����8_ �Q��]�ڠ�VąG��p���g���d+�E���h����f_��~���*�);�0G�R�w�]��P�tKpJz&�fG"�£ ���zFXL��?��K��Q��AJ��'���:���\��/"�F2�J#�7K��6�{����b�r��*/�/NSs֩��Kg�U<!%���{_K��!U��=������̍��a�ȏ��b�'`e3ƕ
�L,RƏ�p:�P&�F���r[�����W���)�s��9ֽ�v�z��Ӏ�͌]f�P�M�R͑�-��\46,i�tӟw�Ǻǥ��O>������ξ��S�ط��԰@��-�I��J�فX� '��x]��(�m���S��R�́�+Xb*'�J�`���FTr=�E�b��@�e+H�DP�����=c�4��	��g`��x���u�1��Mi�1���!��"#d&ޙ�!����)֝p}JJЂ~�F@z�xeV���� 4~�������'i9��΃2ʭƣ��o�s��ƌ
��� 3�mčG`F������K��救���A��U�rT�bML]��֟M�͌�Y5�ؐ��'!B��\�I:ɕN�5����[�?�v�>����M�6�?��wB��]�	�<�B��ž3�t���?M���LPȤ�oT�JD��Y�2^�fgk�R��9�W�k��Q�aCWL�abN��&|�
,��R�BDN��yIH.�4���-+*~���
1+���1<�n�?�k5�I��St�	1jP�}N�E���_��WN}l`�V}��^cz �>�(�����Վ�cB8�[��U�m��Ϛ^1�C�/�X�dW¼�ǯ4�4��ذ��$��J�:��.�^�Y����њ��`5����;c�j�W�a��1ꭣT܌�q���*����O��n4U%`�sC�'s n�^� 6�Ck��W[
�����ޕeV�#}�&�9B��MP/�lIx�Q�b����L(����F�J�oiȋ��x�+�m0�6/�'Zm�Ox�~M p=Z�(_�v�9�$_m�i�������s
"I ��J{�:'�{��fT*p� (��W)zG�߶�	���N�l��� �R���;Ղ������NT(N�F��q����|q#��y �L,��ni�P�\�W�N��ǻ��)q�!|���u��H��P��Zx�֭=U��p�vPz����D�E�jC�[N�x��0%�4�z�1ٲ#��G3<G��>A�֌������J�ԗô�����I�CF���c�~��X���9���"#�e`l�D�Z�& �w9�qfL�@�{�L���"��`�z>�q�B

�I1�f�SY'�7'�5���s[���'�}%}{�/ЊX�k�L�Jp�c�*̀�'{@"�����؆jZ'$u�[�f�o!XD���[�*1�1�u��M�E����̶���7q� �wT�(e�E
F���:�m�-�R��)�����C�A��$;]�wZ6�P���57ɏK����j��VFx���@k��2�d�T��c�8�%
.�i���JNaw��:ee��
yf�j�1��q̫[,��7���T��\�:�����R8�z�̣;!���T�̟[&Y��-�ukؽ�������㙊��a�<��:���*	%��;
X��Z\U68E��/��N'�l5/���>��H������dn3����m�5D�%�Gn�1D�����S҈Se���$�Rkw��@�us����H��&��
<��o㒻"m"��Ҕ<wPO45(�f��8���v�Շ����`�k�����QI\�0����K<�@bd* ���O��tuV�Tb�j4K7��Af���X���D�I��t�;ut����L�/K���d9�SR=�����[)��x���`���35N�N��� �������b��h�'�0�%)W�n�OK�%��7Q���S�S1�W,�>0�m�R��[4Ò�Ǯ�8m�6[��j�cRkn�;��ƚ)N����|E9�U�/{/Q�?���+~+���.Y�:�(/�M���/:NW�>�󀀋���OzS#���eZ�t}�떠��V�2hn -�wIꦗ�&��9Wn�"	� E��"�Ӫ��22g����~�8�Q������O�;���m��/g�c�"L�	3ܤ<A�ո_�cd�۰���onER�"�π����z����3�j]�n���6ϻ\�o��)�"�D�淜�zin��Js@��n���d������h��q���&�"�;��b�2g|+�`(0N��bJV�u�D�n����������$^Cd�劼��	t�<$ Q���|`2�U'a��Y�?F�wa�e�D��sxE╆"¾ ��x0C^2�s�m=-��qh�W��]_S�����-#[~��O�zͫ��HGS�7˯D1�F��%C���Kl���f�;� �������P*��շ�0`i������y֙���>�^'[�l��:�PF����=L��u��p��{���r��������M��8p;N�Tb*���'�gʢ~�r�ԧV��k����o���t�˪�#�u�$�Ŋ�l���(���^;8S��z�����c���b~�/�1B�� )<�ax�nC5�T�$ԉ=�������y�;��%��mK""zp�y�$_���kk�EQ~W����]~�<���n
�O֑|�V\�T�d�*��YA�c�2�w)�g�2:����KY�g�6f\f+t�~�fx'��L�7�z!Ɔ���!�_p<zȟM�ɟ\��!�E4�w�X^����rJݹ��@3H8!�E�9=�?I˹<��\����%��W�e'B n.��g�4�e2�vy6ͅGD�v!}݄���w��'�\���z����8��B�I\��U�P�hБ ;�d��d<�[�����kSjiF�"�hD�T8�a�1'�V�"�blx��$�j��}�L��b�č�p�wP��n)�����
��D�d(RHC�hN#��n����7?�-zu��N*��Mu�c�k*�W|��[���-Ѣ�V(p6^p�$l��#��~}�� ��/����B϶R�y��r9���J�N�U��zbG�uG3c�v���#��r�C,�L�Fʦ����,=�z�����n�{��y H�9��I�P}�gۉREY��~@��JܜX�� //&�f�?N����:�m�ۻ�)\��2&-����M�f��e�9<qr�/�εz���=u�?(����L���56�(l�iߍ���Ǔ�?�T$h*���H���cZ�c0h�i�J\��qYZ�k�P�|%q��X͐~@"mʹ1H���۝�\Q��i[�Qj��ǣ�u/���q'oT�}�jo	��W��� ��ʉ�˄SL��( \�=�{��>���l�p̽�ʱ��ݕ��K[�Cz������y���¾� %0.4+�9I��p:��c��#�֯� �~�����LD"�n�����K`����{�3��+[�3x�@r;��⣮^a���v��c�/T�$c����P��n}Bf���쪊0��s�G9��!c�>Dz���`��} ��l!���<�6��ǲ��#�P��\;�������o��Ft��Pa�t[Ė+��������Z]�O> �\��A��v�˝�[W/<`�.�8�ԧc0���~3msVm��u2��n���z�|�d����i�q#TC��,�a�����FR�C�;{�$�|��0�lנ��ǛC<���?-dUp9�ՓE���S�%̼qkL���7�R�w8Wb�Dx��TQ��ү<xi>F�2�9MS�+V���F���d7�\D�E̺�v|���׋��{Ÿ��S�[����Z�E�=��y���#c
D��J�;(~��lx�f-�G�����'n�Շ��R�ctE�.��¼&9�buZV�L灋G�J��"'"�Lt�]�0��T��)I���T���~����L�H���K��+_ �g���$]��˿�*1�?��$Y�Ⱦ��-:jA.'-��[E塎-�������G�!hN�x�����/쟌���sAV�~�/�!s��)7��dVؙȼ���&�jj��}��]���?��~T�G�2���n"3�#�/摀�L^j�zT��y��Ȯ)Il��	�V�	����']�2����'����:���B3�e��:xN��==��a����5��托q���9@C��̕�}�8z���t,T��.K�J#�c�Ӱr�:�c:
@��� �%��x�ң6�
��w>�̰,��I��H#�jKe�z(��U���z8�u�xp_� _�'��Q*z,�ȐJg#L&���-�A\g��cu��Q���[��t�K�e�f1B8�M,�po�D��n�W��~�����VA�t*�����8�����6�a;V뺂���2��M�N`)���>��4��I�>��γ���p��{L��L<kB��Z���՗A��&3b�����_�BI\���R�8�g٨j�����s�R�7Ͻ��)ق��?�A��y˓G���T�(�F�F�IE�A o�>Zȏ!�$��w4$��+�)������2gf����P�j�Iv�Nq �G�f^�eQ����HWW�Q��;2ŝ�*U�t��m��h�r}�h��Ǟ�Ƌ>,0I�4]��2�^��w��ɓJI
���ř��ұ���w�!�bZ�r��W�����@�0��_�^��Bh�A��O�>s8ڣa�ё�R�����?��?z�v�Đ _@���asled��WWy�ֻڞ����!i�2Fn�^�qO �n����Oy��j��mJ}xMl�D%}C��M�u>�go~��~�k�^�����S�^"�4RNU�eW���͝��VH��)
�̈́���hQO�!X�c�����D4mET���'�D�7��?EQ�J���fⰇg�x,0�����L@�������J��y�S=6W�W	�.Ӧq���ۜ&ؾB��"�Ҿ�o*�C�
9'�|��6i�8䱐��<��S�s$h�ص��1.u�:�5�6�)�&�@��DY�]34q��ۧ�ȵ��YBF�!>:��U��Q��I��.&w�({2d�TW.b�mp������YT�������Ȧ<e�zX�G���&�
��=���*۱���Qd7@��_�	Y�!/�� qY�ѫ�r�%!���Yd{ޮv�9�̑�7��I��g&��Nj����>�t����>�D�pYEg�2��"DĲ��O1"F��X C�,U�M����QX|���(*�����d%nn��@�5#��K���>�$';��7�����0ޞ����k���ލ#4\�K�8{Lo�pȡP#]��?��w�k�ʦ#:�ˊ�|��|���mk����cG�����T-��O8`w��y�^O�`/��*9G�h�~	ib�7{X���$�q_yE�6UJ�R�c7�o���?���s�]3#�p�'ŃD�F�RF��>B?!�>J�E��٨>�1������K�B2��+�ۧ�_�h^���C�\��4��Z��ӫ�d�6o���3�BR�3�F���9�Jz)�AO�m[M���Z$�[0�Lq_h�3�����yo޹N�OvfW>�
H�n��L{>��x�@S!�]�k��V�/�˺F�jt�r��-��'����fEr[�˫��z8B3Ql*�A>�D�<�Z�֤l3{���
dEE�i6�^~$D�ob����Qx�sB�u���'� ?|���>�k�oz�׿AyaqU���&(JG��D�Q�j�Fn�1�b*��i���)n��s?{�*�[)��s���1W��>�سw+���i������'�-
b+;ÿ���lwm�'H~SԒ���>:�s�����2��l$��#�Q��O��!]��'�I�x�o�ݜ�t	�����S�������\EgF>��� �G�N�N�T��O� ��v3�8���	A�~0��%�9���z���-���63Zito��X[�K\���φ���.7�> ^*G4}w^5"��g��F�Ǣ9��`�oxJ*;���J&(�8Q�����,��Vw��z��Gň4�a�8�K`]�ص����B�;�0����B��X��`]?u�k����J�����ՙ -|�D��ir���!�#�*�~�w~�& ���54�ߏ`���R4��fJ)J}�k�.�=K,2/y��Q(��� t��ӽ�1S�yP1q:g��-%�d�Uz���tl�i���1~v+�P�����|��#y@���%���ݧ�mb"v;�{).����y�9XN�8�^с�jG������]��e(��O�����R��.j$�M�ƨ�����נ������_���o���ܮ�z	>NZ�XKn�Ut�u�P` ��D}��mJ�6YK��H"�|VAQ����iU�5����Zz�4��B���5�����{�d���P�|��>]��4u=�Bx�@�c��r\c� ���y�wK��G���o�9.}��76���^.F��?5��E�l�k�bO�'S�7=P/�����b�rj5�t>A����e�u�Ö2h[㆘����d��G`�%	��ǡ(�Ș���-�IL���1N�:�/*�!�7�B���#_ar�bQ��N�R7��}š�8f�9�1L����[{Z��h�[��b��,s��s����=u2E[#��bˎ��w�����4�f������Sn�nǶ�xk#�_�׾���L�||v�����[�u��fy��\F]eG|Q}"�<紑��܀�b�R�d�fZD���$9�f��f���<��.�*�V�!��*�z�Wѹ�T�R���r1�T�y4n=䧿?�Iu$nZϱ����a9<����`�*EH4r߱�U8;�b�����z��t�M�7|�9W�F�#�6��~r���KI�
0��9�2ؤ~Z'{a�MIP%>d�	��S�=h��7�ٌ����7M��)(�FL����y �E(pV�	,J�������F�#\���0GG�H��XV8G(=���9����F�2�>Ex�>t�_b_+.�t Q��q��ὠHr�Kχ(B��!6fչWؤ=�����&��T�̿`��u��L�=��o��E��3
��ޢ�`9�4WkM��X��5���c񋾎��$T(���m��M�
���j�n�*>�1�.��ݑ������0p?��(s���Ρ,GhrMU�:��	�F^�����Z"9�bY4��3뫳y^*(�r�=�+��0j�[燥)8{��\O�����CF�@,y�lB� ��=��4�j{7��B_j�p~k�<E
�>��k � `��@���-���R�f�/��t�&\�C-$��-�N=C�&VXE�naoމ+If�@������ P�y������t	Di3���]��t2tzz��4m��Z�Ju��4�W�0����|b#_��439.��}c����m�>�h��rK)
�.����W�o��	jX�]��H`������;�zQF��!�IA�y����pY�$8�@�_�hQ�$/̄��'Ǣvd���v�O�b�'�����݈,��}�l��@@��ͧ��w5���f�v�S�)�nC��S�>�b���e��CL��}~'?��zZ�t�㉉D.��6���Q94I���a���c�&�
[^�0X�F�z�R�v���h�D�V<>�g���π˶���"���S��8!�|���7A�cWex2�z�\�&��� �v��  �@,���/A+�K���*Y���]f*v1O1:�J�|��&���N[>j-.�iK>�_=�����^֤T(1��!���P^lV�!+t�����k��G�8zy�=��6`w�	k\ V��@!����O���EȮ�t*_��|�ϧ")�nq�0w��wm��r� ZM��R�l'2��A�g��/���೴or�=���ŕ� (:���\�2�`�"�B�pO�q^�Z���e�F'�w*� 8A׸�.|�b �-�CS&>wḊ�	�P�r�$/y��R��W'.4=��ò�lT�]9Tyy�[֚�FW82��X���KB��L������8��ز~- І_���Ҙ�v��%D��k1h�V���hR��T�@Ɲg�-�y�E� �:�r��l�C8k����#��#J��
wCR��'��WLK�z_�K)yc�eE-� `q?̝!���sr��%�@~�~ż�>LC#D�a�Y�Bع��Ue�*��:��Ϳ[��ЦGi`j��g	���M2+��t '���"�Y+g����:�,�6+h<��!f�����XײՍ�d;���9_�7�n��#��y�>N�L��gʍ@��w��9uB��矷�k*䥗�\*/N�E/#�*��r�(7�ub'� �>::�D�:��y�w�p��p���y�ғ�!�7�V���yN Ax|�U�]���e�^�)��v��^/�Du�["�����gvPM��&�̆kPa�d�ե�l\_9N6�1�65J��V���p�G��-t���<��O�Ѷ%kjOQӒK�7����IKθA��v�����J��č�A���O֕��U� ���^X~����S�c�\%�{Μ�o�x�̤��؈�AQ��`b@����g(7� n��[����T��wD� IA>C��E(�#y��u����ȉ�[�r�0�e(Ėޕ��jx�F��,���s���%���re;��Ia�By�49L U�E;Jh��LF�gm	󃴰y'H�6�h:��ݠv�R��A����Z ���e�Τ�d@��;83��~��'}H����<�2-*�r��	���油/<M*ū�;#���Zq��!I�ywԗ�j�����?������ޔ'���]�|ꠈC�z����w��HYK/<�7�N��X4�8�S6��&�:N[� c��
t��_�jS}[�y��?��xD�Z�SJX//ׁ>#�=mgF��0�1<&r�N�� ��v!ٜ�*�6�79:#T�ӯ�v�>�� ��ۊ�=ֺ�8_��c�'�t<�'bRw�m��Cݽ���QT�:�u*��
����$��q�wN$*�#?��:˓�ci���J<G��w�i��'��r鳝?��>��7/�١T/H�ET�������oŔ�I8�ǧ�a�}����ޣ�thn�vXX���Z)��Bvc�����k{�S)Z��P.3%��W��^�g �<������?�U|x��h�R�+B��&�i����ǬQ�5ޭA�ޘ��0�n��Dv�C�`چ+�IV�uv)�<�t:�"���.)+1����L�_#je)�|�K�]Ⱦ��Ξ�+���DR�g̨�)x����)�r�:m�/�� �������Z��^�1̭c7WO5Q�������<�N�c%Or����/�W*q���+˴�VlB��������oS�@`(�ѕ��=��]�aR4+9����B��%���F���f �7�}�kOU�eZ41|+c�2�4qj���:�V��)u⢷����J>���ܽ�<w���0��	a�Q�YZ�	�u����O���J�G>��1��Ϧ�6��/nY���sQRщ�%��灎��)-)e�?�aϣ#&���U��:G�r���K�|�T����<���I��?�t��S���mE�k�d ����<����
�3�kʥ��r�HXu!�V/�_���S��'hB�f����	�HeL�
������3��Z6|>��HL�@h8ux�b'����j�[�?�d�FD�&�� ,A���� F��X��sR��8WΩ
��Os����bSU��,���HCK��d�f�-N��_n�Z�����E����L�B���)�QV�u(jsXw�ek�N��À��$���l�*�@��ت�I�h��$��_:Y�w)��.��5b�oR��]�p�d�SS��\���؂����m�c�ew5	ӫ�A��R-�H4Ͷ��0��3R�yg�U-S�І�dE)_��?���b2w������UQ�}�V�:����9��whfƈC��/��W�l4�L�r{��$3B~M��&������h)�m�x1��"�mYа��X7��*�(�װ�E �`�k-����<4D���o�m��'\��eӘ�V3�4���>p�
Q)&���c1��F�l�q���ݢb���9J�Z�cw*~|���P���K�T��ezVb��r fMx$6t�8��ڃ�/e�'.�0�&� ��h�����s�ia���W��6�{z���q���2^����'5�+QRM,�H������<�Tq ��d-<���n.�ECP;k�!�6w�|��7XSϔ˦9 {�AN�E�����R Thβy���1��s��L�k��I�!�~��g����ؤr�	�y�T@�{!T�лR)�ˌ0$�p��s��|m jj��d�)����G�M��9t��4�bGT��5fv>u�{�����t��;МҲ�DLk`���/�j���@X��5�n��F$)4��ڇ���U��hfG[�g�H�Ck�S�-��4_���o����GC��T��1��������7v�/���E��z�&�ĳ�v��:P6ߗ����H�oX؛�L� � �L@a�k}�A�Єa�9��h�ϧ�z<��c
&�����*x�����|�N���3�zQ���.�ӯ�~����ԔELǙt=T��b�KO\Q$��i��cáE����ǿɂØ+�Y���L��1ch�4[m0��z��.iH�
�:0�<�D@��,V@C�����.H���q�z�9vŶ���W�vQ�ѴP�L*u#��!���
Z�����Otǁ%)u GÆ��un�T�ؗ����Sf�ٶ�����\u�k��l��.��'�W��NX��1�$���N\��Cp�R���E"Ք�ju\	I���ju�R�-m`(CK�t�m�Fz�A)K�97r���X�ga�qJo.� �U��v�|T�	�x�2����XÁ�.��SA����$��7�
y\m2�/��6P
��=Ro�.�9�HW࿬�`F�ģ�(ͱn.�������kq`�-�4�!9�R; |/(��2m��&�'�Å�W&g�����`ՙ4��$�'N;��M!|"i%7_�b��-�(�x�G1�8����E��-���o�_M��D&���@�,�N�y(g��ӖkU.�!�:`������$�aF�DY�dq)�Cv47ɜD>̴��*��"��;����\�����:��5R�|l{��/�ֈ�����3�l$�_=�I�t��:$	H{�]�"�_�����#�.��ɼ�2�f�73�L<kQ/�,T~Bs����ٴqtIFL�(�R��=3�?Ă����u��W�x�)R�fi�$J=��m�FG0�K��v*�h�5���3,�uo��:ăj�M�vBr+"��b|T^e����tE�ðYp\��_�_P�Ϣ�X�t}aT�us�-�Z�3���t�5�����8^�Vu+¡z��1�Z�8�&��s���F�I��\	����^��3��zm��cg����K��\����y�ʭRfTr{81�����{=L��<�<T�t �]7���w�Fw"��O�M�s3qSu؝W@<�6��:��,��e�(��9 ?������ G��IY����o�O~��R<��UAL�����e��O:�D�+E?��6Vm�&���΄WK]�<�|ͯ��#���Z�Xg��yq3�����iٍ�I�c�P���N�W��F�{�Ȁ���qoaR/\�Kp�������*Hk�$�Ď�Yf=�s�#<�K�8eKrh�z�'Ֆ[A�ƃ�#[�ܻ��f�a?��"&K�J�Pu��8�j(Y������;��� �~���fpJ��T���/�>:Ɨh��ق����ɩ�Ea��1T�JY�zVVY)]>�z���ճ`ۺ��3�|ӱ�Y��ٗ �B`����_O�nC4ڳs�����aEĵ�8х
a�t������YU�R�]�\-}�J�t�z ��~���)"yY�
��	\]jY� ���K�F��Ļ2��a�*�M��������MGvF�V}��+^\��r~��z��zC����V��ɀ��npi�U�1��z��٘ͮj�O]V/�/x
kl�9U���N�!�-�6�Yx;��lث�!���!�Q,���a�m�+��$)����"��S�J�"+ӂT�[=���u^�p�j,��ђe�yz�̥��\&�Cp/y8�5����G;S����(�`L��42��+������W�~��`���ivz�$��WfW}*��Zr'������;JR�/4�̥̊�ǁ��2���$A��*�>ٳ7�M����r������pU@x>���p�0�q��l&)�K�p��qv+g*ˢ��^��q�K~w���R�'�
ߢC]������[�Iܢ,�j=%�G���p���l� �bf8/H���_u����g��L:��~`��u�c$�k^�u�H+��2�K��<����,�xh��^5�î�˼0�MI��\S�.��f� ��E�.|>|�?�����c6�t;acu7����ӏ.KW�*!��B��3ixx���lz6���Tf�Y��uy h��&Aq����/	�A�������0c���P�['�cq!GC��m�E�	 �u=<�J��fP�-%0��L=�֬+g�l��O�|Jޟ>|5���r&�AXˎ1?YJG�z��<)��c�d`��&D��¯�j�(���t�e��r���V��~a�4\�&#t�0h�kv}l����	�-/I§gˊ���:�.��Y�"-o��،�(1�0����ʎ��v��!?/�ʋ�rt���ac����:��T2c�����{��p򚄗tGO([,��Ԧoܒ������D�����ؗ_�7����$��^�Y�9}p	s�
���l`Fb8}�~W�O�93���!�O)�����G����;�K1�s�b�2v1�b�O]����ۓ��v}��}�@��< ��V��6�J`=���a3�	�Vϣh?@J�~$�G�)NE!\5��~�@/��KU/Q�߷¿3F��^�-�q-G�B��L{6C�A��F|�� a�t	i&����gM2�U($_��n��%�]��ԉ2���Ku�8+�ej٣�0t�#R�or�"H�8�i�{JI�.�����k�N���F<E����)-�j�_��'��7����AS�g�ͥ����)�Dy>[HYnB�.�����J��б����Mr�����.Ύp��+��ρ�y�*�Yo8������ݹ:���=.zHj7�s�����H��ރ�A�	�v��$�=v��?btё���A�+�g�Fw�T���ܣ�$����V(oN�xT�3�B x�����ܱD!u���: s�������-�[��Gd'������wŇB��r�}�k���
�ŋAub���D�W�/�n�4S>�_q<
�t�(�(��?c��� �!�ΦSVQi�O\��t`{�*|�$�\[i<���D�=��~�تm���#5�&^���*	�b>eڿ,�j��W��j���q!����I#�2�wL#�7L�4�)����`b�GΤΑ�(�ב��X��Q@�\�NCs����c$�I� ���B%5�q:K�*��]����u���%6�� �C��<P��;������`YD��AkI�u�p�����mfct�n�b�5|w_����q����C��#:�A_x�=��䃸!�9�ib����׼��d�� ���� 
U�I�pR�K�Wn�Ob��Ȭ�L�Ά<�\m��!)�]wM��ƀ�Sdt`5�J��q��<z���|YWmŗF�u��}�8���y��c�fƣq��:o����X�l�U��7�uw�����[����Ĩ�o9FX0[u3���H^�k:?�}���
������� X�LL�����ߠj_~���T��y��~y��Q��N�:Ԅ �p�h���QS俒��w����Z|.����ɷ|�ѫ%������`�i��F�B*�/|���Bŏkd��XOs�c����w�g. p��`&/������h�	��ae��L��r��'�r���
'�h�k�P��;����M�E��v%TCц�3�⴮���~���T����$g�@�L�"j�_{�� �/��3��l�����B|�6�_�?�XYy�Ym����֟�~U0(TM�'Y݅BP0^�F^�!o�Y����>w$�}MA ���㛳�X�a.m
^Y�p?�Z�݋��ZK�k�lH4��}6�R���q�В���W8�/\�=���i�ht<�f�W�H�s��x9�v�XԜ�'�2_޹o��Z�qD�	��V�FJ�)M�RH��u��7�1�+T4O���5۫���f��HoN�|��& a��m��aF>bp�^I������y��{Q��X��S.p_g��2^��&���ā����g�����x���Y�7|����{E�o2�ˆ��#h��k���.ЅNȯ"�6��
������Ǩ�r3 ~Y������kh���T#(UP��V(w�J��j\d��"�q:�,a�w����i9����Yܮ����h�����z�Y_X�x4��ŧ{,� y�_ӠȐ��W���=�N�F
 ���@���&�'1?��ƶu�<��I��=Ĥ�����UR��f�`�Lg�n�_n��C�D�J��a���c}���o��Q8��r������P�x6z})�������#w	ֲ��ϕ�oʃ؅-Kޓ�r�G��ɢ<���O4?"Vs����=ϕ䯆�5��LKH�*Do�\d�r �l�DD��*)�������S�1�4T�t�L��Ix鲍q$�P�piV!u2��Ҥj�!X��c�+�p���q�$䋋���h�:����C���EBG7K�Z�� tڟ�R*"��T&���/Ji�hv6���ZBKf���WL;l��Y�6���a���)@u�3�Z��I�i�)K�k��H���*Q��]g���=�z�J!+���������m��g���3��I�A�r<"
���,�]��M����/h|Y�Hg݆/���jڼV��H�t���l�o.��V#:�1A��i��m:�4������N������̶_
�j+��>�y)���K�<T��[>I �����^�g΀[;
V����0�L,,�����	��d�^Ҫ�:y�����������]R�|�)�� �Ԯ�ܻ�犄1".���W�1����_����#W|�,D=�F�j��n���1	�2��X���M#�v�B����d���*��Uk(ߍ2��Ῡ\j�d�3�D�H�t)-_�/d^C��rk�����I���*ZU<I��i�Yܴ,
<�x0PQv��I� -R)^f����EQ�S��j��M�-ȻQ�)���)|��.��ڥ�+vt���y��F�\��{HX�`��m���A�E!��9�y�9Y.�o��n_���gǥ� c:7�#t=oI=��q�F����h4^Á(���∏�.�m���J�i���*nt<���u�ع��Rn�s.1�\��k����PZ�����ǖ�'�2��V��N5�
s��[��Eh����֮_�v��-y>g������y.ӑ�˳�@��(��b��tV�U�5���k�r�r�ݦx�e�����c��j���<��\i����.�J M���Xzz��=W���y����>e/�MD}�X��'E���w����A�7���2\�X�N~�N��7>2��9~�>V���ȓrA&j�i4��KyИ��py���;�y�K�3Nsߍ�-��u�1�@6�1�+ϝ�������&�J��-�Z��%2q�L%�*�p������R5��Z2�reQZ��9̈.�aM~
�Pï�$ -w#�;=��T�7gۛE�:��n��b����l	4����fI�l�iIB�=Y/��Lڇ����B��i�;� ��g�\u?���^�!(��J֙�t��F�Q�z�a� f�v������L��mD}(���|��]T6�krz�,�E"���К��b�̖W|����:gՙ �h�X¤{��[scqf7#�2Cy��NL/A��P����x��A��z�2��aѽ��Eb(N��
3�֑�v-��x��������*�+�Q̏���߉?bc���t�{7sP��I�p�J���QJRM�-c��������+F���a�w7ʇk8l��c�>V�h"��
�ʑ>K�{���5����KNK"涡�B�Se�+�^4Vꀍ���P���F�0��B������l��橝6E(�@�F�>Ĥ�<����!읓�<��0� ��}�%CP9���o[�>;��y�Tn��?��艛Uµ���4	��6`9�B���#%�5�]ۮ��g��
�*�s�^��NZ��o�c�S"��۸�Wr��|��x�7�R�k�Cጮ�7AK@�πcDaT�Pu�#?�dV�%�J�-r��e�����8���8�~J��� �t"��}�a�$Bs8����[�� yl��� �M�.��Ɠ�9�G ��O-��½��#H���
;��E�F�b�I�$=�0��/R͑a��^�1�s�p �7���._���0��y�G|�a�|ÍF�`�^�r�a�1�s��$���.
O	��|w8F�=0}w�+�z�h4��g�Θy6@9����ɦ��bZ
)^ox(�+��2�Cvc�]i���Ԙ�0��;���c��V�\��
�`�z���ݑ�l�Q���t�����d��_F��|b�����;���"��:��B
�M��X�F�eN�劐�o3C������u�O��q������KH�R���焥�5N�YO�x��>�}�䭴C:7�1/!�䐺̟���e�;`/�i/�-�}ě��ٿ&�Gn 8��܏��]�l@j�1	�@x
��J%�(a+W!�Sڪ�j|�O ��P�z�����o�D~�Gg��L�B�z�
��#\�N'�p�C�=��A�,R�%'1%c������N(����w�+IG����Y\$H+"2-G�Ŀ�����)�h޻)�k��A�&ʵ���3�����Լ�v�O��iA��-�6R���ү,-�� t�K36{ɠ���&_Uq5�ף8��l)�͕6)�߲+GM�z=_U$b�;b�Ξ��1{PB{�u�43�ѣ�Y�e!"�j]�шF�ٝ*Fi�^��46�.ſ����>�G>`(��,}⮜�{"��uG[�|�����������6%-�.R&��J_h^��ypJ�Sg����x6BUJ�˰-�K�'��*��,����X�=����5r��r,�T�@���X
�(��>��U0;����<��o��E뼚1�{OMpD�f�J;��x��w�~���=~�~kY����`X����Z����J��2wB�d�����q�e�T�4Y�꿕>.?�1(���oB��5���U�9�YiXG6.�7��W����:WL�Jh���J}�eo����9R�ˤ	Q�Z���C����9�]��ysx���ܪ1�,f�0��6�F�	VV)F�H���A�T�}O�p�Dn�A�BN}�������?�KT�����	��ɭ�D���;�+���+����$/��a��E�W�bjʒ;q�E(���Z�S��h�^c':6�E���i��jF��̣fJ���P�!$�p�8�[9�g�f����'㟿�	�)��q��{����#U���%�Ҏ���Z
��.�O�{��u��V-{��w�`@���\nJ'��dC٦�y��*����SR<�������U-��"�s1 �\rN)�����TMUT8��zsn��R#b���@��Q��?�u՜��!82��cXR��$�X�J$��LCb��O<`�V��J�1�a͛oU�>���T��m��J� A���{�؋�'�5�9`��@]֘%�ε�I~��x�kN�	�$���_����(�Pp���}@�e��4j���z;�ac	Y�?SH{�cn�K�*��֒�>�v�z({��)X�&�f�×�^�� ��f֧7i4g�XF�f�[�� ���t%�8p�F�F	��l���GJ�6`��Z#��U���9Εtz@�nx��y(Ox�~ֽ���]e�<z���*<���F��v�ʐLԹǀ�e_j�x5�"��P���͢��#���;�U�9���qJ���N�*�8Nɼ�d�C���*˄�i:�E��6q��W	�L#j.4�|�t�����'�G#��!}�^��Ni�F�x~�u��2��IՂ��X����/lf��)��j,y�ɐ���ȿ�!��X����	XqA�kQz'�X-�H�/�F��E��+��6�������}{��8�\�')F�j'$o����o^OF��MR�; �t�h1���3ϜL�(ʋV�v7���ƭ�fz$��ŀ�sq���ZP��
lU���$�@20A�hꐐ��tD�n�7Q�q��E�-�?J�"��_��`�H��O2gn������g�r�j����?�'�C+G�م�[�<q|vD{��gۼ��� 8G�.�-_$�KQڂet$^�N���c:�g�(DVL���LT�#��[��t��YWd�uC�<zP{�[�D&�C��[����5(��7.UI8+�^��[#�_���W��WT��H3Ɗ�$y@2FuC\��H������Έ,+�ˁ�9��%S�IS��w׋�_�f��1��n5��{y@p'��V�ْ�1�hO	,#]B�w�6
%���9�l��x)濚�(��!rL�`�R�/�qf�Z�E$��I�T��B8C��[z�sB�����m^�7��ғ'}��,9��
�ᅆ�tթ�>���Ua�����Ĥ ���4�0}0�$�iBA����%���4l���Y1�z�����N�/�A���ݠ��{��a`��ao�J�j>���6��X�:߲�v<͞�ҳkdӉ�I>n��2�*�!0?�H���$z	�zqk��\�4��n�J��侥)�~CM~J�o��h.���,k�O�N�����"%���Pa*tj�ݘ J���#�$d����k����X�r��M�>oĠ:��f��TL���z�KO���Yg�����gMZ :[�h�T���q�D��*�Z�i~�ė�f�WF���}^Ns*X��|�.��}jƿ��*{��9аƋ�ֲ�D��5��؉��iǖgR�ޛG/Lĸ�}�&@�&o��[�H�3���&���r�24�����_=��(d	Y�v������S}w�YIi9��Cs��o�f#��f5���&�NL�_]r����R`Cم�R��9��������z)6-ዒ��&�-�R�{'����;,�]?�3R(�A � �)J^;���7�M&�w�O�ƞJ{�R�s@~��$�ƿ��lDn\���=����ߔ�&�s��}�)������wᔇ8�T�.CaX�ȷr���6���,�,��$ɤ�7HPB�l�/�B�6�`�)�7����A�T B����3�!]a2?�l\����H���@ G�FI�+��J�#�#i����:\ ��������%�{ւ��6�lZX�Z��:�)�/!"�N]-������p��w�Y�q�X����d6��dΟ$���R��}	5a��"^��ض;��a�����nS��8CK6�8Wu��6Q#�N#Ե*]6�F�|?x���� ���4�P>�P!�!󚒤���?����=�;�)~�vH9�M!}�,s�O'qQ�lr�}�\�8�|��Y�l�c�@-��-��,|�y�xF'�A;X���X��xgh��G���\��HX:VOGz���_�b2N��j�g�i�E혫 ���J%oPP��?Oߪ��`H�ݜ��h��P��Bg�6B)���p{d11 �4mߘ��gg�"s�-XwlgyB���:�4I#T?:�g�Q\bMX8ԻG��F�m�ϸ�(����sٕݵ�t/"���D}�
�3>ˢ��<�s����9Ѕa;��0�:mR�0'�|Uzh�������&�˧�7ٽX��	堆��O�	}��(��e@�
����Һ:H��� ���� DB��#	��9��"�S� L'����s����b���0�����t�-2�"�׮_�̚M��7j�P�ӽ����r�@9����#��칹���������"F@Υ1'3<��<e	A?~;����D�u��yz{Q��}ځy^�;F�x*�?�
>�'+|F�{��Q>�����6�-)��}xQ�[߮�<ǰ�}�Krf�F.֦-y��]��z�<�eݝc���#e��wv��B߈Q;xA�`'���l$����&��^k��8���Ӆ���i����4���10]�L�����\��]�Y�^�-��?��eי��Q<&P��;��t��G1���BT��LV;����9$�?f!����^�^"��!�w����O���� f�b(���^f�[^1�۳ft���]o[xA=SU�⾀B4z�x�<�x0�t��HØg�N=���N�/+j��i��+��X�����Rָ���Z�
�4a����:�w�����~��3$S�E������zk��˵�w�əu��̩i8�Rz�%J��xu���J�h1lH@�lx	����T�g��9oA�e}� ���*nE�\�-���U����HܛO"����'�a�������d��2o�;F��g5ic��\-���5?_�(4�w˘�+�|�<C_�;j<��>v��Py���M0h8�Y��%Hcz}DNi��-�p�-w�1 ܦ�[�ٵ/����F�[T1ݤ��-�B �K�@�#�AY����ry������Y�7��K\~��qc��vB��2���I�K��U���o��D���D�,��,s��
6��I6#���wA����R�)
K�1�f�t�,����dn�@�a�Ö/?V�Tx�%��i�m1'��I��
�t?gp���.il*Q����� ��0f=N�R�-������v#�?[��[�G_��05�R�'�-Yu������K=��,�x�N�(��|�����#�E5�)���h���r�"2���v������`�2[���Ex;�(�.�����J*���=xT[с�5e�6;�r�B�%D}'��AxWT�\ۥ]�/�{���/�-e؉b��d򋾲>I�u�AQt}�ʑ�R���n�+�`g+�S��i���������[*=ZO}��O��e��ٝ\3�D	h�mHӕ������֛���2vKXS�Y%@��d�z9��W�	[X�	J1��_�S�B0�[�13�y#�X%��_6�ҵRC���� wJ�ԯ�$�q���m�<v��hIXE�Q�n
�W�� �
�����we�ޛN�X�u�u_FI?d��g�9w�k6i��9��C1��D7���{�p�uq�+/���˹�R��);��.���"c�FCq�C*Ś�|q��'��Q۹�K��T���`�O�N7h�����)a��]��7/O��ݙj����soT"�d�Bp;�5�F
��2�u��0��@����mv���D�� ���X�2�+_��;&���it��*=vP�OȈ�R߫	�s��p�R����D!���:.�ʣ&L�I޼|;M=be\9<��7?�G��n��/~����w��I9��>R���e�&�&�oce#�`趌���0���Nw�;���a%�h�.zExĩx��>ᕤ�ᠵ�ZPG���G0 ��n85�8T$ڱ(� dp�&����~Uʉ���ǂyĘ�Q<l���^V���RKG�����]� ���#;�TGg����ww��3�5�;Z��k@.�S��d�e�6.N?R&~�:�%k�cB\e�	�g�p'�V������3���&\�RW�hC�";CKP��&)�����Ѓ�"��?~��Ǫ�	��<���%�/Bb�� �뽝���3���V~�������J��w^}(w/u/��1g�1t%6Xd��;^|<��Q!���*Hi��0s�塌��yw��(�J+��1�~ԃil��A
g����3r�g{��H8��%��u|�s�ۭL%`�N#q�f���V�m�
�lFV���i����.�Нt"r`��%�l�@���y�%>��H4XDj��^?�ڳ�O���2#A>a�K�S�,M��6,��E�
�E�F�@�y��d���$g;}gt0��6	q5g6s���k}��IW�$��ӏ�w"��["�i�5^�����ZV�`K�M�dI��$XR�,��M��K��V��EĶS�	��.�9��_��NwZt������n������Le>�C�zx�b�����B�p�IBu�@����ֹ%�=:i��麳*�3i�[H�0��6q͚�'bv��r{�������j"Tj�A��᰼��������`���*�πI��:傐6��hbN�b�~�|TeJ��v�f��)Ҵ���F�|e�'���Rȹb"�`�Mh�����UX�=�8�m=����=���Ί�{q�s*�woxCו�L�a�0���1���桹%x�/z"S��Չj0�D	u`@����w-Ý�~�N!��f/��uOr�y��Y�W��b�))�S%:W�yz�~x�]�	�O�1wJjn���g8�ى�Q�Q�n�.�Fg���°�:j�}�$���SO��\f�bU�6ĝ3,m��GH�L�`�N��� uA�h�{0h�5��8&�ȃpĿ��ڏ����\�{狏��[֋��#n�eƏ�k���ڄ���_����M���]���)�/+��X��xF7�~r�<>�|]���M ���k�ZjCL���
� ��u���JrG~�ξ��<�H�l`���c78��n�+�,�^��*D'F�PӨ���7`�1C�����#�XZ\�Ա��_A}�)�$��j��xgɓ+TP7�j��ƅ��p��8J�Ŕ�B6�z��]ݭ�X]����Q=rnl��C#L�Ae�z����҅�'lx%���)&Z��r�X��?e�Ѣ~{��=!�G^������{ߋ^␷���}I�+u�_���	]Yr��߮��Țe�͙�������g�\��?%�w�_Mޛ�����^jC�(v@^�d'���{�{���sD)
l84�`U����n�f?�?z3��
�5�,�V���L�Ϭ�����=��@l�N]��$T���uw�O�~���~�Z����7��AKIL�I�rd�IqSO04\~�����U����(�er4�W�H�"�&e*�g� ���$Q�Z� W�Vf����y����%b�	�I���"Ț7RG߫QG� ���8a9#���''s�[[b����m��.���"��&��Wv�$�&�8�!�cz�\[kuw����r�jǁ�X��o�Wљ�s��E�I����Ī����T�4�~�S��H��ʺu��㎼��u�pzO`G�1G!@3f|�8�(㬲��h��Z�I6m��9�\[ �
�.x�Rd�5V\�z�Fn9�^/��i�3��t�����(��
a���h���V�V�k~�W������࿞J6_�4�DY�'񘊕��] �`2@�X�KN�gp���d�8 푙�.�+�-��˃���V��1NG�a .fvjA�%)$�|���6r���=��zv/6��l(V=�˟����%��2���_�a#���9���6=(W�u��гF�V*O��5� z�'-�w�m����4O��0�ju+�nY�2-pK~$~']�9���x��Ƣ�}�_/��W��m�wxF�E�kcO�_ø"��$�]��K��廯1� ExC$�g
�gU���,�����v#=q���5�_u4�]"㸦/�WA�#��T�e �x��3�.b��[5�KI�c�Zԍ2q&r�pޕ{{�"�Ie�^פ>Z{d !E��
�>h�����[�y�KE4�?��I�:�t��E��f�F{�il���ժW�ʇӏ����E[�2/��JED�7-���Y�V��HBu���B�|%��G�Q�����Ƿv��_�ݺ2p��P�	w�6	j�����r�����a�ҳ���+�k��b����o1[���|�V\ M�+�|/�x�"�:R*1��'�/�?�+d5JWr�,�x.Uk�t:R�i���$�w ��T�io3�g�!��X���ȕ�WB�f�v��*7�����v��e�)��/����R����rEj2���M��q|�;�e!_ C�w�2�,�{[3)�qKF��|��#[+|�XX'/��j(%!��eڿ����O�Rx�4+z��z��1V���>�.�.ºV(	W�Wo��
?6�j�O�`BT�p4P�]�$?�2W������&$Լ3<�F�w�F����\>�s���A�&�����$-�$Ea�a4��ݭB� m!�^���V��*����[��_ұ��a� <X� j�&�[����ne�x��#��>�îu�	G���-	�[���݋*��hz���Ľ�)),X�5�D��d�
>�p�a��-�@A�@ck7��y	<e�Ʉ�g���� ���E��Yx}-պʛ�fj��Z[0�U�}�"�g�
���7P�╢V��	���F`��/��T�*�i�e��2��4�>:l�c�>lS����"��M���.�4����L���w ��}��$��k�Sh�>���4�(h��L�yi����ss��ٶӁ��op��՝�J\�u)�_����B�d9�]���	�{�lq���GO���̯�c�8YR����/D���1o{�k���7��:L����g���.e��**�pj�|vI	�p��.��F�a�`,�یL�	���������1����ޯ5�2#"�M-�y�+��8A�3Xc{3{�}��A/d��f/Ӷ:��~�Mi��lH� p��[���b�(���E�U�3u5���P��� MG���zk+��)t���L�9iۏu�A��P�
JT&:���B!B�_�^۝?���+�[Fz�]H9�,|�bNBmO��4	���s�f����+���y�}KE�Y�YV.H�^{E���z��ғ�
���lFRes�!駏N��=��AsQ�]�T;�*�|�B�D�*q(Y�^�%�s0@s
�K������e��)롹I(�W�bsߨ��J�{��B<���[�Țn�vm�t�ʞpE7g��m	M`�T�`:wj@H��A��>#���W��}6o�,=��3�D~��F�:`�
ss㬩t0빼��4�~����z9,����D"��S��+�9f��Q4}�S@D������Zb�����e #E��c_�E�JT��H<��N��@3MU+��Qk�;��x.�2\b-�0��Qn��!�Xx�˂�����,KR���}���[L��N��Z�Q&�v0.ZjM����
NP�Ax�C�K�5}��S���'��8�2�cRŶ���;(9����2�н�g��^�4��ĸVMu
���2�'[�Dώ+u��3�dӂv��
P�!l �T��n������W[�z�u � v�����8C�:��w�{K��8��@��1#7��69Ӎ�&����*�>�S7Cn���J࠽���$�x����H��+ʆ��YbGa!��=�!o�l�ҿ�@م�?�9��aq�k�.�w_�а�*ڿ���z<t뛚"�5���
SB�-���z�]�r�1m#�YUC�GLz�E$ǆ�7׽86�D-��j䚭�|>��a���2����Z�M���2�gzH7�2xF�%��$�wS�3��KD;r7�O�1�o�HEo�,�]���~y���g:j��j���Y��,G�x���6go��"�j��ԣ�%��T�n?dw0C�}�ќ�D������BT��zC~�E��/Sq�/����Ҥ+��7��ƹ�Я�3ǆ���}P��#uy!��(N�M����63����Q �:����)��W.;���}#?�E����e(ޯAǝ�䅰�u���v/�S�}���~��/x6<2���XV�*2/!H���`frpp�����/k��C�� �Ԫ���UN��h��` ���$T�r���TU� �
$Sǳ}�	���E EߜR�� a��%.ytpL��c؎�H��vq����y�y#`eS(��m�V ON�w�6 ͪ�P�IŠWe�{	�;�\���ǖ�.�������@7/\�a �*���&~���P��A�)(�hޜP�5��d��ʴ�l�ʃ:�������슓��)Zx�`�\soL��\�X�Y ��Q��LT��g�����_�^Q�aI�j���P5RLA�]{1�{���[>�Ĕ��l��+	���!m��T�5eI��*��gh��0�gz���g�cY�a������5L�*�����l�§?M(�ڃ����G�|{����E>D�w�L���#��/���Z~FM$�w�����_
�AS䴪��T���d�1�<�-����[�^�Y	J��Wu�F���׹�|�U��Fx`-F4��J���2�_�m�~�VH��*	W͍m�)��jBK�������.��A�a9������3��	D����At��{�cw� �'�Z(�͚��}�����s���`�V9_��6P�����B�h)�`�O rm����Vpe�����DC�F�4�t��W���4�C$�_�_�<7�AG ���b��!��S��{m�JHuz!�E���U�J��DI\�#�d�߁,�E�n?�����.���*<��b���>`<�h�u6�����2A%KK��e-�����Bf��x!��0�XX��:�^j�&��c���Z=���UV7]�	|�t�zo̹��6��E�G�n]��lVq�I�=q$��;{�z��?�6��R1pX�2�J����Yț���5�g;U6k�)@ɜ��a��&44��$M���#��DE{���`g\'��>���2 s�R�˚���W�B[Mix���$��SP�VvRd�%/0�?0OK��� ���ޏ����_���;p��i��:(>�����s/�N�;������R_�܊,��5KjL�alٖ�tl D�X��x�q��]o&�q�K�dt����@�A�B2�!8$��#Y2b*Y,8}[�IP#s[�R���Wf���"4oR+5t��Ǩ�Y���nL��I��&9�؄��&�=Y̫�G3DK(�s��c�X˛jjy���2�y6��y�f(>���ɝ�%[tj4�=`�B+��3�����M@.)�����!�˼�$��J!^P(�������/��`x����O	��" �� wR钩#ou����s�c��'9�;@�݁r��&�	c���?D�o�F��E���l����c6��A�cuֲ��~�>t=_D�˓�:��\&�ݍ�6G!���;��ij��F�s6��Mq�8�s��Pd��?g�PL � �GF�y{�f�
��<�U*�Cگ����9V���Wįxo���ߝ'��tȚi��s�o3���x!�
.�C��p��*W��r
�]�D�
�s��f�{ �z{�2�|�t����u�����Ҡ
n�"Z'���X$��)�81u��(o�,�������i����ZZ���-�OwJp��NT���z�D 
[a��c�$�k����Ń��O`r�P������;� �(%�l�*�7�3�T�18��k	��I M�طк�VW�eWD�ߤ��JE�ZfuO��^�J����5��������L��͂���h�ݖ�f*��E<ȿ�Ȧ}!X���J�֪��ꐊKO���CqA��vSUT�����K��J$Y��0"��K���n�k��	�)8SJIF����[^�sG��kNJ�h�{İ9ߢ�T�b�u���m�6� a��|��,�MA��T.-���-]Ӄ8�@�;]�4S�Ip�n�I"O�6G݋uV��˶̻����nE6n��b��T.�J�r�s��0��(aW�u��)c]��z�0��o�5#gZ������Fa�!�"�_��,�i���� ��ӷR:�&cF��1Ʈ{ޠ,r�,�-L�P -�l��P���&<���z6
�ܧ���U�R�6�;[!PaoJːz���Ӣ��M���^Pi�&��a�4����HQ���z�m���D�U����R���)���7�`���#I�V���O��O���j�>u��%d�I75G�O����oH���?='W��=/�xϳ�����.�sO�hv'��Y���$"G�h�����+a���c��5%9P�>Ȅ[��x���6}�%P���/��� nu^p�rA�&v�v�;�+i�'��	��@���o�U�TP���S���Opz�(^���X%����[(XB�k�3���w�꧃e�sb-5W�2D��X�OJ�R��ve��#%NQ6\]&~�-��o3���e)�P^-�3��g��p������F�5Ba��H���Zn�Od�ה������u0�Zp�t����Ч�I;4O���J�� X���*t����N�z|~
�[��&~�+1L��tM�zS}0�"	�us�2�JMv��a�#����R��ũ��W������0K#�gk�u6>���!�|���%�F"^\o�>Z��-�"��%1�?�Gn��e���	�{����2�o��_���
�G�C��dN��\d���x?��ꂱ�b�bۂ̩U�S�R6��������7A����2+�!.A�}v���;���v��Ij�e.Q������=���F�ȥ�չ�V"pe�"W#�=��X�ꃪ>\4K�y��ʈ6A���)��m��9�b�G,��^IKo��F�.��ޡ�N��'�`�}�Z�[�U(��"�&�Gd-� �5�|��e�xP�8k��O�!l�li �f�Fe�c�8�Pl=��|��9(�$�K]M�J9c�*�w��;�%bʃ��=`	��:�MHz7^��|*�)r���23���
�B^^��������qx��&�B���;�Џ�Uz6�,�k�Q#!��y���N'�GH�t@��s"3B�U���������}�Jj�3�!�wRt1�0�"E"ncq��_�J%×X�栬\���/��b?~-XK�FRk���j,Q��z랅z��߯Q�p\m�*�$��xAH2�E翿�>��$�2v��+5���%���L�L����� �1Pz�t=ՋǱ���o��
�i�x�~��'���?�;��fz�h�Q(�q�7~ES�uR�4�A��������[
A�'���\��K���.�$?F;�q��$G"o�Hr��(KbԁMN��H"��cS�7�2�����*��)�o��Q/�S��\<���x�_��0�"�۲G�����0��*�`�Sls_�����c�� �V���-�go(�Y��h���ݪ�.�S�����1e�'h�kΦ4W�T%���38쑛�#t��w�����?9���\�a!�m�#��`V���o��6�ҵ�:����!h�@r�ψI��
�y����+/��I  9)� ۯ�	f^'9�����4��F�,C�(�Sc砷�Ա�7<ik�����W�^˰�N��8M,���'���h�M�VϹ�$��գ*��8R��e@�ÒX���n BMjR�������QΗ�r¯����p]:kF�727��k�&�Xi� ��%;�����az�� ��x5���
P�@�����U(�&��PCN#�$�-g,lk�����N�t C�����;�֨��ڛ��#[cZ���ݿ��˭q� L�
A�	J�F>\�8��#_����Eyk[�>:$����;�1Z�.t��E��O�����X#�,����mc[���f2E_;��Q�����a�]�?L�	-�j�Q٩_L��_V��$�O�Z�ù/����2�o�pI&������q�a`�r�l�3��#(T[���p�'Ѽ2�έ[��ڝ��e[��+�K?��JK[[�:����11��ߢ�r���B�UZ��[����O�����$�1ѕ�6Y��v����5ǃ8Nc]��z����F�$��Y�VC�'�4%Z���Gs.U����)g�>�3>�D�ᔞ����L���Ο����ě��;�{��|�6ĩdyl�p�L�2�2r���ATϹ,sj{�5/	cp�AOP݋���Xs�lb�:b���#���8�ܝͯ�a������NK�$<�e?@+�+���F��U�72-�}��W;�I؉�R$a&ѥ��e#{�VF��a_͝�7��T<��V.S�Cٷ�`�nz��I�E����A�o;�}��C�� ��i{~l$<�V����j���� �g$��:�=	�B^t;�n�B��gs0��V�/"����N;tT��Irk��Ĉ�Q��M���tǼ�9��8);n���1�O��5�3o���EK&��� �M�˧-c�UAxp�S�D�/hT�hcPz�c�_��:'=c��5�(t�h�K���#�OY��dxk� ���}"	��=�=��������%�{?[I�$��dTE��"�P��Y�m��j��qޢ�:��S{�S5!Z�_Wj��p�{A����).����s�ZK�7�1V��=5�6S� .I��d���T��7Ʃ�{
�ۓa�%H�-Oo� A�Z<���A�U�$$8:6ʒd2OM�wi��a��'Ǜwt�I�<�1�2L�B����
6������Vt�%��u`޷�j��(I���6of|�q%��R���AWW��������#�`�ב��soS�*��+gn-j<7i'�r�*�~3���>��H��{�=����:�K�i"�VZ�rD��Ok��?V	@9�M\ ���!0��8�~)��&:g,��>:��F^ɻt�Q.�o���V�F�Z�e��ͅy���zoKE+Ќ't���4;	�H�������w��L!!�Â��`���r�(`#�&&5BگA��!�X2Y.O���c���oP�]�9���V!"����v'<0��"RL60�x��o�[��K���E.tL8�V�
�n�f.=:���8.=O�2�Y������ac������*<�F|��&l��2}Y��j]p�t@��R�ĒN��'y�?j'ꚮ�*/;��Ѭlܴ�QG~%�B��k6}��z���z�V�6}r,яb�e�!���>[̇o=�Kb�v<A����Y�< [=�9�n�;΀��	��v9$yM�QL�� ���L��t|G��G�U�(0ۛ����GE33J��KɆ����(+�Zl�?p��)*�r�F��n�p���0\jś�� �{��\�7+hmr�p/Cy��e1�$
���s���j&��,����/� bdKV���Ǧ%qޚ:x�����f߯��3 /�e݋��4u�u`O����tjcZɵ�6m��!@=}�*��K��Х4M�0@n��i�\I�(�+�Zm<CH	�G�`-��3'�KER?Qom$Ft �7Y�ӯ-�L���2x\S�fCex�Vq��DP����|y��?P�w2�=vs ii��4����I�g~���l)���/��n)�%�y=���M2UAgS�O��FN�|?q�FT�����R��E#ܱ�}�Y��N-�4\1�s]b�8�|oȿ�D��W��W`<���)j��-�{�"�%-����k�SJ
y��(q��ɫ��a����O��۽��	��Xª
;0#�
Gip(C�e��eZu��F�,��$z�ā��t��Pt8;LӺ��4���sK�I�&���І�gw�ȧtI{���)t�$R&�P��te����ao�����yN&ԓ�w!u���$Y��H����\{z��P�G��P��c��CX�/���4�Y�n�V39��X��`��� bz�8��!l�����v=v�Ŷ�mn&�.��":z��� Z�_���S�ڃ���2f�I�*^ r��.��ŬM^ט�p���̨<|N�����>=+�Ksf���!X����T@Lj�X5���Ӈ^?��F���T���	E�ԛ��y��2��:�8犨)(��~�{{C"�"�� {B�/�t�Z�Q�r?:�yU�&ֿ�J�Dd����}��B��L �o���I�i��0�Gf���-L<�4��dY�R�X���XV�~�� < ͉ �7�����(�tgo�ҟ�t�r�� �_!bk ���tۣҧ�K~���F(��6�Oɨf9�@L��6��g�(�rՉ7x���0�|�����H���F@h��f@왻�ȀyW�r3)��S#�h3�S[x*��A�RP渖�O>V-�X}��Y�T���L�9��~�D0߳���Cc�{�$-�Xl��M���&����]�!����v���?��ɲ�=�|���"�};�t�i^�,����p��e/�h�s�h�q�Vg�ڜ���mR�Hy�F8{��=�����G9r���-���0�6Ѩ~l�R᎗���s�����H|��X���C6�@��r��;Pr�s �u#?��w��Sè�cѴ>࡫A*9N��Z��bʔ�(�B<g(�E�swҔ���J(�*�%I���V�_l��`�R�G�AYWΘو׏�oF��p�����O���MS��r �؄}�H��/�Ɏ��f����g���ɮ>:�s�cJu�ʋ�	�:6<�i��z�ee$�,��UY�g�	u�㱨�Y�T���s4"QH~H��	�|�ӌ����O����!a@��Q���' a�Ԯ'x�sxT"z�!B�J��J��ƺr��;[U�IQ�(��� �%%��?��I�̳����J4�{W������;�^<:�	ѭp�r��*r��Kv���z�#��:�.ܭ)0K���b셻۾���y��rV�[mL)�S�e!hK�M���֖W�b"�]�E�P�����5�1(Ж�����kC���|'v��٪?��W�v��z�)�n�Sɱ��N�}!��r�C4�����v���]���H��~�/�Y]8��L�?��-jS�h�Wb�R��%3C��$ď��E��vb[H� j��k_:�T�c���<�H}!MA�y-�f�+P�!v�6�O����1���"�"�OvxV�Z���ރ`�*I�2@���+%bj˧�1PYlC9L0o����W,٠�7e���#��p���zi��r��w72���=�Bd�
m.;�my0.�T��)���B�"����I��ά栱���w��<�J�:���hw{�1�#k��>�$>�(�)�`�Vg��ж���a,Hގ�<E���.Hzw	s��>^�Mܲ�n[����He#z��6ﭏ������ k|z����ʒG���=�!)��[��`�R1�W�j9��O�K���zq�~T]~�n~c����?I?����/��5!?n2����L������e1 iaru�����f�㎵�8��p���ܦ�
�$���N�nLO҄�4�u������؝���_��7���Ff�@�I��k%Ĳ�����Ѓ�Z.��%���*M
�{ȫ�ҍ����] A������9?v ��5��$���7H�Nwi�`����]�Uj)����|U�ݫ�|�Ob3��g
D;�����U�N�� ,�K {m�;�����S�6F�p���l�r�%�/Й�����_N����)�k�!�狘��l�������H��*����eM�İ��̻��|��e�r �\A������~V����Ã�`����W���i_��
��{J�L��a�^�?Zs���W�y�y5��
<湔G�q�$�}�f&�q͹��aqM>[Ig�]_��/&I	��l�����եnT�"&��2t�ɤd�v~�����N��z����4��r��i����_(/���DP^��r=��;=�1>|�����E7�;6�QڻC�aN{����âR�/�7�������Nx�m���!��?�2\liC��%�m^ʆ��~3}��}F��E�u�p3����e��i/H��" �ZnĦSh�B�N�����/��>xh�E�s���<�<ZQb�h\���]��v�Z�,_p��i��tj@L��K��Z��=����c�(.���l�U$<<V.�^@z�9�]�v���h6�㚮�u�9�fH�f.?�ڽ�M*��p��NC��!��_����a��)̒�׺��_�H1*�#_���{^U��I������;�+}�����v&��2��w���%����?��4�K+����Ts\���L��u.?z�{�}�#�4������1���kD����u?J��Y龮`&D��W|�e0�A��qrjh!���ڏ����տ^i�\�Gm��� �:��l���=�uz?Y:�҈�,�,�����}@;&i�Zbk:w��G;�c��������'�	b-����`���Pa��ɣ�L���#ǆ�} W�G�`��D('�F�l�S��ܙ�R�Be"���i�ҭ�ʃ�N[���#)����P�����8���ѹ(����(��8�Z���)�h@*t����EX��*3�ֳNR��dW�k��O�@>���ޫ�̞b� ��ʄM���NP/��	��B�y�Y sH��hކ҈���u���-�9�B�6�x��4K�_����:�|�u�G�
�X�Q�/�FM�>���=Inw��K��*Qǃ�{w�����>��M���y=�Qc�ʈ�N�!Ǿw"B�v��4ekģ��ĺv�B#��BgΒ����-����wK5��6W�ɞn�f���x�ܾS�b�`�yZ���Q�>�pܸ���2_Ǽެ�p[��Mz4r�Q����c���)��t��S����L��x�\�M�\�����V��k��k��-��c	6
�P�����L\2��v")'�>��j��$�O�_-8]�6p$�H܋���A�M������ˬ�!�AY�U�P�����z��	P�ұ��ʝZh�����o4�C�v5$�4��L�/ă��p�}4�οfܴn蜪�8��0�4�>V�e�
i���P��0�����2�@���7gX��,�ɒ4��#�a�s���۹���&���b��eh�71 ����Y�mb.���6DhO�!c���=1�C��;�����n2�.������p����O�Y]�{�dnl�/�1%��r��G�O��M��on����V=���t�3YS|�}��^=�F�������o}�&�|�Y�n���ǉ�	̔,@M���W+}�Z����g�zk��#��e����3�"T��Ҵ$Hg@N��Q]r���z=�"���׸�����Fu�����_9��r�����+䞪b�����U8J�0Y��Ƚ���d��0��`Xf~�\0�2��_�c�<gϔ����rO����\Em�_������~�6���ÎS�s��4;��h�c��/p�TR�.�I�4fh�^�V#|N5�Nn$�e� ~	q�����ij��5=����X
������ʵ�x<P}�S�e,�D��yU���/ݞ�8�8d��frI'�l��oq/5K>�\*�pD�x��4]M�`'Y#oEt'!�:K8׿29Qkt������(!��'���������~�o(���p�X5�d6�	�l�C�y�l8�l�.p%ї�Z"��B������4D;q#��ƈ�^�PTpU�/��Z�MCҼ�g����y>fcW�)`ǒh�M�+)��x牽)��ڡ�5�Z�k�":�����B�b\�s1��{������/�8��K����f	�n4S$) m��W�)��.A੮�\��>�`�Z<�Yٹ�o����<�!rNq�$"�o0d�<�
]E*��V Z�j@������O�j������2�e܅�����(�:��O��,��`��.F����^N8݂x���\i���$2a+2����/��V�z#@w�-�[|Sl)���8Ȗ\ٱ;�j#mB�Pַ1���h�@�Se3(J��	��\�*N/Fd&Q�P�����q���")���i�U"�D[R�ʮw^������.���t �G����B�|f^��g�a�<8a��� k�������ݻ<�!�lW�(Skn��ǁ����3�m�\��j�� *�x�!j���C��J�4O��ӚH6J�f�5K�hV�����w�icGR �)�фu�&�:�uN#m��c	��^#�h� �#v���;s��w]��y��&��ú� e��geˋ/-����p-��-����ͤ�D��{��#Go�����!k�B{�R.�9�O�c3|��m̱^Ǌ�k
h�KRȠٸdʓX6u�� ��O�oo�AY�J����)`L��m����O��O!��X�j�t5?�{��B�DFs�<���S�Cē W�n�Jv�5��9�N�
���nR��M�9
�3��1�Z΃Jār���$�?�Ȕ����E�]h��T��v��?����o���eZ���:)�^�k`��XEҕq �8r�}ů왫���M������`�/��M��[5E�>XL�higkZ���,�ZŉN;���/�/!�C6�,8����v2h&d����/S.A�����p�GH�j(�0Ù����}QH햠(�˟C���v1��O�G���S�;���$Y ��k.;\�ۣ����ݎ�X�0�>`������9�zz5��C�ȃ��߬��R1�@&�6:pa)O?�>��1���Qtf���|9l���j	R_�a��fm�ַ-��7��-iK �6��g�%d�X&��2#�]9`�\i��H���El�9�}�,x�����|P��I~�����e�
8vIR�����I�*R>��'n�;y��佭ْ��߬����+{�Sn�V6ǷӀ�&^*�l_Ґ�_q�D�J2խLe�F�<1�I�l-�.B�&����x�J��@��b;���[?��İTyD{��2��@<�Ir�Ɖm�γk'A����#�J�2{;d��ZE��G��vF7W�es��c}�w�fA��Ǜ�[q����i���Ep�,��D;G<I��t������9�7��g�ht����|(}�����](V�i��H�QS(x	��V���n~r�nr�6\Q�G�����:�r�x��q��O��,3V7y��~.ֻ����t�?�4�P��IkV�����ö���IsǪ"� �3�.�@�8�tj3�uh��\w2��9}��U3 2ՍH#K⛤���l��\x��CwB���s�����f�_����
W3��]��_�|�O��x{����+G���ʻ����Wj�bxtf�|U�r�c�la��qX���x��>bpBٳ�w�+-%�RLTU���7�y��+g*RSJ�;��c�ָPޅ���������J��톜���lI��c��A��9	.�_�d7^�L�<h����O��ģ�����q?�h����7z=֘��,�\ؑU�ٶ�<f�ܻ�k}M�E��w՜����G�v�۔R�}Y�h��v�PCdE)�� �ͷ�z�8#R�Ò���Fr������z�v��� �n٘��ju�q���U�o��BJ��LK7J�6���gE��l�c�%�,e����	��m��ݎ')1]�� ��٦Z��p�Ы)4��Fs�L6�`�E6Į�@�im��L�{�MA
/!���18�8��7����9iS�9�]��Y�,�Ay���B,j�qb��B�@��RP+�ЗP����V����a:UѾ;X�#�׍���d��q�g/��?F�y�@��B��/�]:}�PH�O���Zϐ�AE.6�6�FZ*�:�ʩETH���C|7{'�
������$��&-�ª���<#*��0��>�d@bJ7.�L���:��E
�Uv�~����y��c-�(�E��OÄ�Y���K��併�H7��z>=��x=/{�K��������bEQɓ_K�3W�{ޥ��A�J%�J�%܀��o{�Zm���Ž��|m$�Mg�r�y#6���3"vK���I%�XB����@ۗ���L�Dꮲ{������'��Y���x7h�+ħ����]�ד->Zj�����m�8Bs��V.����Sk�q���Z!��W_l=Y^��gw��ʺr�&�{��T/�i�LU��qI���Ii�>��?�[)�'�oٰ3�����<K�٩o�D���:G�>n�m"0&�L�S޽m��j�8ОG=CI����%)t
J�����E
?�?Ql������_{�%����xOs�b9$�p�o��+l>L�xkx��wDԙ~�<v���,��R�r# �$ ���h�,3[����zxb����OAVJ��Հ�Q��G�v	�"���-��kB��`3[9�k!���Ώ�&��.�����T�l��P���g�^�{ǏX�8�j�e��U7
��W�Qj���+�m�r��öv�:v�[_tD}���.&�ջ}�z8�]Z`�\Is9�H�HO���.���7���0]e|�}��m�@�u>�TĔ���ЫB>�;0��5�g5��T���hS���#�i���ڦiz�a�0���]3S8�T-�
�����yJ��$��]�Ux~�XR[j��|\C��
@���6��8#��h�D6�VƌVn����	��8� �\tMi@����]̙K5�p�س�H�& �hN�Y�}�+��o#���_��/m�@��kgɉ2���rӤ�� 3j:����oȐ��H��h׫�%+���ȭ�{�j0��J(\�����>��o��܏�5\��1�ѡ���6��Q�񲎗�ј� m��It�8�4x�&�i���	������!FM�0k2�C'�M1t�����ʃ�����O%�k�+����K�?�]6!��tf2Cx��/�r�-Ŀ�o��k�I�K�/��0��P��o,y��~��_r�������6\�xhV��!���@����	��k�s(SR�&4�8-�m�i�� �����8�xU������uW�Y�{!VS��;�'{b����^f:wW�ٌJ���� �V1L�[�&}VV>i׽]-kJ�&�SX�_��ذ�����%�=X�0Xm����s�B6�:��d�G��J��
�W\��ݐ�T���{�E خy��o�0O\&05q��Nf�K�^/�G�}J[�4���4���M��lCͪ>�J�*L����p�φ���0]�w�������WW�4ņ�x��Tk��.�֏Т��rh;;E��#y[���������ɡ�s��b��d�yr(i�Ѐ+�*YX"�n�Z2���WO�� .[93�H)�c���T���Ekp�����\�AS|�\�?�>G�ȁʡ���bЁ���'���S����^�.��G���a���M�H��~+<�����H����#�x]�`����+���YWr<�������uzlfh�h��j�@����M(��XO0��5��\���C��q�m�tXiu��v�~ܒ��_�A�@�����np$K��HSt3ZY��Ѣ�L�R0K&2�� +ߎh!:�Z^oS��)�CDq�g�]O���9����'s$�Z$(l�,��j̅�|ԗ�Eq_
䢦�oJm�j�^��?�����'<�� H
cG����כ��_��7�����F��b��y��K�~�h�p3A�z�2T/�'��v�.�x�o��BM�ݞP7�*D騺������A8�¤̎:&^�+�Lс-�-1텡�	2��x ���e1?ڒJG_%�*̩v�9ĕ�-�-����i8O1֝ˮ�����B\�#��vL�T���X�Ds�n�)���uk8�c(�L�7��&f-�ᱝ�;=x��U2���*�W2�|cN�M]N�Jz?�q�&���M8t�[��s�h��$��.��QS�y wQ��CWm 0+��q���� ���H~����-�}���e�L��˒���+"�{�-͔1���U�C^�z�ME	V^!����d�t��<���LW6`n%��>gp�Rh1�3ys���u/J�ok��T�$���u�M���+�P��eG�ہ_s�3�y{��A�vl�5"��S?��V�e�b���?�=D�F�gP�?�?g�	D�j\�����Sb��t:��C�G�l5B�3K4I�Os�Y�D��?�(l�(�wƇ���q�{WK<3U��9Lp?\���Zf��ܿ%y�eR�5"b�2���{�EX�@��Вy$�t��H�ؒ*�ھ������4�E�OHi9'9}UW
�߄��UDo�鲜.:�~�#��F�H$B$<��k<�TqfG�i� �6\�<$�KS�RѰ�7����\�R�hɦ���_G�>*J����0�;)z���X�n� ��@W��s��UQ��l���,�A=擷h��
��Ih�*���>ZZ�#%\�|(��F#��1���I��D��;w"J��&��m!�#��Ux?н�\��Uu�ˎ����r��b�Aa�u��B�5l�F�2�L���E|}z��
J[ޢG�Pv���ov
��Z@�赨�R������{}��:1C����5����dX��a��"~�����m��C�ȏ�Je���|O���Hy�m��`l�.�q~�]χ��Q��E}+�Lϗ��7|����PN$�+vyo�1p>yϫ �p�M_ ��Y�`���/�m��E�w$K_�7��/�:�����͎���H_�-n�������<b� �o�yĸ8�(j��΁Ò���B�˃���y;+���g�(����n���3��c����|�t"��',�R��νRA~ڎ]	��`�<�t�U���(,���+��y�VT�+���R���k�e�/��Tj��Y�Q����@�9�Շ�UDϠ�4f���ýB1l����:�O�N���oG�}��'�`V�!rRҊ=��V] ��,.�g'S�%QkGm��3*���x��1!X������N�����p�����[ˬ7N���%��4�Ɇ�ГD�Gn����be�J�dCK=R�C��MK	��-5�_dFM箩k�����pg1�>�d�s����E�L��G��.�N��[Q~�7L��i�d�tuБi��I���=�7-1�#D��ϼ����:^Mm�CuKխ�\g��a����@�u4gK�(���6O\&G���Z�s�$��3g�f)�i%#�cx%M�s���j��B%�ޛ��G�2�[�����G��z&F��֑����bs��z&8FE@����[��7x�rݵ�\s+2��9��Ԯ��ҧU�0��`�4�ь�¡D;Y���*��l-�v�ə;�Jd+����u�Pz{5��Z�Z�
H�����z,�8�#Iv�E���M�ݛGѕ��׋�>Os���P���ƅ�����L鶻'���C�kX��{6��8��S�-N�׷Y�4\�c�<�T_��c"�W>�h�df��CZ[2���Ief{�eJD�3��fX4����k�U���邸�h�2�v�S���5U�e�������?���*1�u)�:��Bt�q����<�d����(�/�w�C�iU�� �f°B]��Q���@���5U�c��Ԓ�iQ�n��̚����Z�R~��p~
mȴO�x;��gFvwh��өqw3��m��MX!o0�]��t,��==�:DCX�y�?(lu��c�j\�О[r:<8CSy7�N�dn��$/����4z��i�8D���q�W�Ġ��5u�H�T�9�0�d
G�o��!l*K�*�ّd���QN8����S���(xs�T�����O0�`��`7ρa�&>���š�tQnw
���v�c�gG�v[o��5Q�OI�w�����E���f�jB�UA��ۏ�|�ǍM}X��*�˰��̖�ݠ��S�4�3tG��Mx��~��W>̈́�]��M^�5R,�]2hH$�:�sDD�F��>�o^�� �F�{Foz�	t9�䷷�5���7�t��2�-���n���RiށbuOUla׹i�tB��r��N���N��;_kn��[�f��M�F�4�{�d���%��`�˶�k%�[n�����p��/��㸼!�1���5`|�l�yW���n��ά�p��73MT���-��1y����Ia�m�/������fz����LL@�	RT��+��\���n�c�z�@ZJ /G
���
��a��r�������+���xU�e٧8�~`-q�ox�����`7�}6�2I5rcK����2��j	G�]�\��
��6�u�˺јd��3}�]Z~��S�L�=g8����O/�_,����'������F��JE��jt4���P�N���s��-Y�eo�Ԕ@-Sx��t~�|5pJ�y�~/�j;g�A����3d#N;�˞�����e�Q邜��>6c����d��LcYl�k����K�7~^��Z�҉?��A����)2q��.M���m4l.�Ѽu�����o?m�yZ`!���!M#]���l�5wN�5���n��2�Ҝ�5Ud��L C���Ml����W[�:;	�u?=�!��%E��Y�uD{G��)n=0c�-��3i$����0C[�6��Q^=���_L�Յ/d��,����Z���l]yh��ۦ	�����Z@��,��.s3�}z�/�Ȁo�����$R�z���:��5�t�VcZRw���m伞o}6�j��"vXO�e<N���[s `�r���������Y!�s������p��0�zW���)�-�М�gA�{(̈A����Qۧs���7 �\�`� +�6H�l�E]��p05ꮰ���\��B�	e�_��*�R{��x2݁����,j�0��G".j�1�0��$�bqhf��2��5�A��k�\z�V�i�\D��d�ߺOf@�"ޣ\UV"�i�g�]��H�^5i�,�@�h���h��9ٴ���
�/����Y�-3��PECsZ^>"_"}C�&�5��� 1ϛL�O[űM��:��l"M�r�l�������:�>M-����W䫎�Els��D���
D���U�b�-���j���ːc�R�>�h�z�ҝw��5��k�a��Tl;'�ʫ��'��F����?�ਫ਼��"��n�����:�.zI�9�QB�;g��&�gU!C��g��IYj>�5���pqG��*[�V����F��u���n*z����m��;_,u�r�7�� H�<��=���9��n��Cu�x�}6:�D��A�	��U���i��r��:�ES=�^�A����l�KI�|�R�r�U$.�P/���6���l������m�w�,N���Ų�V��jPlb��6���e*�~�W�+��y��5�u��Bf��f��f��� ��_�+i��$g���H�S"�k���K=RbhX�?Z'��Q(7UO�
���a�YU�a�2~�g+����8C4H3_y�ޓA]MxB��Ѵ'�TM~�?/��g*�srH�����C�gqG��t?8	k}�GAS�fZ��D����~b���?���k}��ަ�8Q�� v�Br�2�Z��;n_<l� ��0�m�{�3j�l�)i�k�m#�˚��4�۪��.4���y����Њ0[�툐�~N�p �!�p���8���;#�y���F� WlW����`V�H*ʁ��a&�Z��GI�}�棄�f���ڟd�N�$Qm�;Ը���I�Y�R����G�7��=�q�t�	��U�����8?��@��N��2�\{�d�<�gt���HG_bҩS���,�@e�3��L�B��$��%SO)�E�;�<��ִ��3���%��̭7���jd6a���B;���D��Oj�ZV6�D����V��z���1��>z'�������r�������'=��9�a/�z8���'�U���֚cQ�K)J�L|%8E����6��������Q�)���%g/[��E��[����u����p�,�*�PC�SyH�1�����J1^�qe��XD�*)� ������E�8��XAx�-�;!6Ix[�.�L����Ԁ�H�=i����!����85�����n���]󐼡�Y��m���di��<��.��#�U�<�����i8Ҥ�bv*�eֲ����c.5�$���m��a�,�#� �f��䉧�VɹKB��P;�v,X����,��g��M>lO�+�"������=7|ߡ�HF�?[��0�����.i�g[�HQG]T��v��?�����q�h��K~�Zc�^��$���F�Q���^�3y��ɁU�ب�ȴ�jؙ���u굇�,��y�hE>S
�	�m��;5���+q@�T	%-�2����1،,��/{N#���Z��}.[��e�7g$R#P�"�N\�C__WL��y�¯�� c8�xf	����
P�]�/O!�uĆi��/����.�fP�CW�\�+�H�0?�e'��?�2�Ru�+�a(r���X#�g�1�[
!�6{�~d���O��Ĺ�ڟ����t� g;�����fh?�rE���?���f��N#��D�u���uJ�V�&T�"�Wd�D��5W����X�,<�0q~�l��$.i��V*�2Sڋ��� �����
���w��cJ�g�4��:�D��'mgoF%\�3�Zi�3�s��k�cOW��w(���`��d�P�Q�-��ֈȦF�Otߩ���e�C���?f�TW�����i�|�M������Ї�t�0S��N:��q�QŦ�ʃ��|Rq�4�E?�F`f	�����B�M?��X_���r��!o�Ac�S��D�N��RV���H�����߰���'��,�B!�6���b�2��V݄\�:m�8�`KLA��O�#��8�If�5U.T�n�b4�&�B����H�1�P�؎��J1���_Y�dš#�Nث>�I��G��X�};l�fG��9c� �/9R����]@�_����<���6�o>����� ������\�G�u��ɼ@��:/�Ѓu�}.���2��Ɲ��h�o��ȅZ	�'N[�P��8�d�br���,2��wKqf�-���V�"��0 ͎Bl Ӡ���#|���V#Ĺ���-�|��2#�����Y�ah��g�[}p����=���h�Ob��Qx�E%�c�X1���9�QM�⚮���#�G{̓��y֝�E v)�N��spj�x��9������!YI<���ߚ��$#$��t�&�v2X��	I�>´�갅�����v�z�Mu���c�,�w{n��l�gŧ,�%�$ܡD��\�D�
��r��f�?ND��e�n
��6�f�̐<���O��7���o'b0�����r��Y�"�T����� �vo�(���N�yU}�Q��k�Z��Dw2W��Qa����cz�x/�I�FG���[7t��@3���UX��3+��o(]���O�0˒Ϡ3��;s&y���88r��VC�T�5#	f짦<�ɽ�z��,�.��+�R{{p0Y��.�$x�
_�_]R>?��]ML^��dn};Uԃ{KFK��f�8�k5�_��$��>�/��-&a�1�t�Q�9��L�f˜�!�Zəʫ�h���9`k=Br��o�{)�\K3����HX����ǂ3fE�� Ad׷Ȣ+dx˅Rٵ~�3���s��ѷ>D�IP�ߩ�
���±)z��M-o&���U�kiA�Íט�e���еt�u7�/�,~v!ҵ�dX��qP:��SߦS�M��Kb��R�dH�S�'O�O'�B�c�
4�-8BX�Coʬ��o�|wY��f\o�q�8�iG�S��q�}R}|�Pǋ틹��o���Q�?>,�[&q�m��'\p��Ƣ���/;&���]ۄ_��u��Z1��7������5`���T+0y��.Ī�K��jWɾ5�H��\��|���#=�KGE!+��TE�
�
}��k۷�	Ai*2&��|�����7T	,���EpZ�����zm�:z6�m�6 ҋ�� V�>�ߍ�0����
&x��T ä�#+��>����SM�b�<�Ǥ&�m����Ļg��AP�J��ߙrxq�t��*�}�| �d��j���������T�e�w.���!au;X��8��T7<o�ש]�$���Kg�s�0^�`�)�nk��.!J�����~�+A\���W������G��u��׭28�.=0M�E���E~�QɣH���;�e��p����!&�t&�=X+Z9t�f{��V-+2��$�huy/K�8���p^.I+zn���㲐�:MYj��ܱnm�ٵ�]�� ����;Kl�e!�m�:;J獴���V��Y[���e�ż��oppէϙ1��*��
��J��'��tֺ�++K�Դ�U4�!�b�ǿx�\��O�M�㟻��8�e��k��ݍ��B>l�0�^��h�F,�^ �M�r�����e�u�"P�=����ɛ�%���¸^��{IT���lf�Y^��#�>p���%�|/��C(7s�Ɍ���)}lc�0#��k�ꋨ��<�GY�jm�̠����?ȓ7��ϖz�_c����:\ɘ�L$�3az�S9�N���i5챭]����:a<�y��e���j�7��#r��}�-���)󊝫k�?!�ʨ�{,�}.���acU<�V���K�>%S'z�D���y�>;��������P�����&�^�ɐ�BR �Y��5���h������#_i@X����YB��U..���]��R�^�B�����c�z�Ղ�$�h��L/�pnė�����ۡ(0�jW�}��g	�i��-"5H+��za�?1ZY[�]x@IjeQ���i~���
]�)��/l�-δ�4�\2Ͳ)��K C��s�w�z�U<8%,4��~����!�8brZ��uߍ�vC�����g��U����<�=�2n���hzD��H�ς���Z���	���H6�*��Uó�ڧ�3��j��ѕ��{��W��m����`�*���G\���Q����=z�ڧǅI+��?b��T��c�V\���͙e��� �+E�p�rƯ;�)i�ξ�E���*��~���[��������2׀��#�e3Y�H�2�K߻5���E�4x�U|����]y��[�:}����,��}��,����PO�&��s~��݁O*��&�싉���u�sWlI��P��'xC.�x���	�q_��� 3n���O�ʔO
��OxMw�7�N��~,���={�?,�W��ի�֝��h1�V@ӂ��jR���͉�K��e|s=�b�nh|�Ǐ�[�7B�p�l/�WV\�CL�fbo�	�`
���gV�������!9��R0�N|�Z�-��ؗ�6�J(�li����+ڶKx��]�v4ؽaa)�Z{u�Uh�Z�ȵ��'��Y-�;����������؏�dc�����ܦ�,t�tCs1B%��*�% ��^�G*>'�!�~8$