��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�8k�)9�k���J�f ۘEN�R��>�Ug:�&�1�X�,l�v�ZBΟ�%?΄�͂���z�B[O9ֈ�b1�c��a���߿����6뾽���K��bP=�?�id�q�*���z�U6N�$�Y���R�he�~r9q8���>Nk2H_l�B��x	}U�~���w�IÌt�=�u({O�lw�����޼#�D�H �(9��i����T�S��Z�0|0��K�CF�>��D���~�$�F�1^�1�5�,��Y��@��O�WY,�eU;+<�!rR�p8:�U���@.;?7J��G�z�(^��Rx��#"Z~���O�31��o:{V�K���ҘY�$T�!���8��u���lA\Ϭ�4A�p-�����8"z5F��p�k�^jX�de�O�{�|̖*��)\XL&�Doe5]���e�q��,���N0��7J\k�`�m'������T��sq�*�� ����[��ٷ�ZÔ�. ���h�M�>Y]OM8?���j�u4"� /�3{48�5��Ma��=^�91�o.�E�np��хjEh��x�.��#���檇�	El���4�Q�f�v/hd97vH�j��Qs)��o����������=y�!WɹPW�Ѥ
\��͉$Rn�>F#�'P�� �4˟���k
!��K> �̣zn��uG3Y�?�eOso@��CpH�i �VK���N�|�T�`�f<ο�����<�[���FvD�U�8<�%�K]E�],l	�rB�r����5�y�q�Á�������hݮk/UFN� �{�����?@9d����v�?H>Sä�Q*D��#i�j��9� %�A��㉭jZd�lm���COj����w�t�gTr��`�u�"M�9��۴��R��z�ݨ��]�kS=��g�"L�k��i�j�.K�1�s�J����|��F�N�ny)�I+�Z,����P��{X��
�󶁓ߢK�\�t�D����R�*øxE� }l�h�z+/VӾ�@P5�2��H�ݏTF��O��+��O56~?0�z+�TW	��4�0�K)[��!��#<�P����&f��c�H{��Y�$��`к,�`�߫w:��3L���8Ӌ�����]�t��$�	^��̲_+$�%�����F�8oM��T�(�����	�fJ�8�wW�[/�
�� �~�gDN(��o��6���
g	�#��z�����z�՘��O`�qE�����2®�\f�@��&~�(x�X�( X s��^�p�|��.{I��y;@cPM��7�S{b��ع��&���'캞JH���bI/�l��Al����:]D���]��iWbl��LZt� �����>J}Фu���A���z/HB���=S��.�8����@#<���'Gg�]?ǵ2����8*F�Er,����Ju�5 �9��S�T�楄y�@�U�hm��3�[�ɇ�3\��ޤ��+�Ǆ��]�Avqf�tZOJ��ӟK����~�!?���!٢��sB�����\ɤ�\%��}�(Py⪨�����ڡ����*]asD�3�g����6S^��r��ȜPAj�����O�)��5��f#g�OY���&n�ڈ�" �F�F�&Z�
-�_*C�7�"ӕҩ��hB�&��j��z+���(�P����/������L֡@8E��|q�y�Lֿa�f�._��\,;�=�A4�3�{�`&�>��u��F���D�A,+�P��:)}!Ku��D���v��9|��\q~M*-S7��y�rO��u��f�Z��G������k`QFO��4M��}�5�����m ��Tvk���|�$N��.��|�@ѱ3,ɢ�3���\of�
zO��8�� ����|nDMQ@/���.���R�{��)�]�9�����d��W�I(z'���u-_����(��9XY+�E��^�E58�A�W2����k�9�)�p�0>�Is���U�-��O�l���\Tɇ[ʦ��:,�Rt36�?a��ȫ؋�g}g�9���$բ|�mDP.N]���T�yk6z���^tه "��P��,�f=�l�@���[M���Y���N,��}�M	��\����$Yo����t�3��U�L��e��+9�}4�`m��veQ�K{���%tr����%X��,�.�9޽���[DL
m�w���K>�-�\��뭖C��i[�y_�K���O�RP���TQ���z�LnmG	J��v�D#P�Gs�-DC3F��M2.����ݿ���5g\ ��e�m!��	@�{ɳv���Z\g��5p-�͚��[��JKox�����p_ۀs��.������̪��cv�4�t��� ^�����n�ߩz�Z[[�0��b6��=7/Qρ3�t� �q{�\�.��J������Iȭg�|!�A����y���ɀ���z�s�T��&(5�A��Ula��¦����N��D��$~ҟ�4�/��s��]�2��9��,�Qi�s�6|C���5i�} OǠ��DX�w;E�L! nV�tA/ag�+��)8��8�N��QB�߲Χ�1�!�V�@��L#h:�1�4<4����ε��o��L��j�,˓髉i=r6�v6����3��]���C0BԷ�d���fp̍#�\���o�F�����,��O�c��
V�aHwh��'HdG���ο0�Ѝ{g$)�A�FT�R�p;,���(g�!0��YV%t�������,��Hp9Yp���yal�_�i߭����O"��"���f��0��-�Gv\�����b?�iؑ$�F�֭c��ۓ�Աp5�h�b�b֗aK�t��s�p뗦�9*ј�CH>�E���8x)�p�S-}�e6�Ҫ�Cܳٮr�����\�K�MF���H��ű9�H�G6N�%�E�P���rko��d$n��k1�]��s�?�C����e�(*�(	�ڊ��x�MG��\	�8� }nbR��wؒ�e�ʩ��/N�EK�c����������G�����I�e�Ѩx��^�Q=�w3�Q�$��'�mqC��L�G>�)b�=��R2`�T������l�%T?����$A�XHR}�=����0d�T�s2D�ܒmq���p�����?,��C�޻[�[غ�!���w����r.�����!?0��.z�4��!OlO�0F�ן�-[I���3;#7M�-�t�6�a2y�+~d���=��k'���_��TЬ�z��2luŀ$�X9�bX(��Z:Z�hk.�y�W�Ћ�,�
��b�Ip�j��6�t�Aɏ�u@�ѡ�Büp�>��"w�c��+e�Gz��n:�Jf3�`q)�װd�Gb�?�Oظ����l���}FQk������x%�f�t�Yy�k�B.���߃������d
��%34Hnya���$���ؼ|�L������|}�C�������J��,�	}r ���n�N�q@ ��ee��� �5��$*�W�ӏ�I��%�����ׅu����,�~��ތU���x�~A�;Ƙ=���C���	b�U�9����6�J�N����)q�$i�j)^��X�O ���#���1`E�k�x�����<	L���M`�z�M�T�7F���K��&���&���N�GhIwA����!'���,� ���i��7��K����H7�[� �CÕ��$��j]TޭQ{��SQF����w��d��zER�i�T��!$
��>QD
l ���8�2��Gy�ǥ]@`U��c��������S��(J�H'v���i�	�O�z~]^�P����~]���2�^��h�w�u\�����~F?)�0�V����e_b�͡�v#�� 8�����@𶗝Xa�`���)>�+3絵��T�{�ţ�����r_]f��Q�HK0_oq�
��zn�^��ۏ���:���,Q�P��$
�.����ʖ
�ǹ��C��Jm��U�Y>�k����wJ�酺�f&A�������r�1��G�_^6�ɠ�1� H�8'T;��.�M�ńt�J�@�Q�B�8�&q�T*�24~���G��O�Sg3�f�Z����,U�a�E�`�Tq�cXp0�N.^*�1�V�`^aP�߲�;�xa���vR9����"�,�[���WcKr]#�"nQ~Wb�᝻���<=TQ�N��w$?t/�������[ό��{-�Zw�V��bY����I�w��>�� 6!���QR��4���OB��9�M)+>ڹZ,R+�T&Q�!�M'R!����P�S/C�ƃ��V��+������/���w~Is�R�l�Z�uv��8�W]:t���fS�}
���B)V�كUR9B�\�ը��l;��/2��#ꐥ���U���ȏ�_�W����H΃�w��R2�G�RG�⅗��։�&Wya��Q����t;��y�d���B�?�6�,H��i,	�DF=
�L%~��uI���cƨ�z Oi+�.s�j�G5�N�)H�9�7~5���{�_#&�m����������vCY1׆t�	\��w�}�W����%}�_(p#�[\s�yxs1ɖJBYߛ��v�*qT?/�y���A;��R�X�t��ן<������\���鲉wK�f&񵊛�u�hpÍ��>z����Uj+bA�����r���:0$�#��瞅�	C����IgT�FmpInc�>�R|��'�Ne��H*HLo5u\�Eo�GJ.�-[�rP����#��-�׹�8PV	ۉ쇳jא� O�X�N��ࡲ��D�=e���������0|݁��^%�L�4.˹Ѯ�3� >�[����,�a[��=�i#Ջ�WU�8�5�r�6_>�z{�q����r�$�Zu�.w�c��֞ޟ*�p:iHl\������2	�di�߾W��f`U�ea%.�~�[t���R.t�h�ga������`j��{"CkE�7=��� 6p\֔I�ʖK�׈�IP�L�.<����\�|�ȴ�-D#A�=�����%���w���6�|�`B�8�L�fQL}�,$u�#g���+�삋��Պh����؉���i��F�p����a�����+�ENDeYk�y�$s��_�WCG���u��8�c��!�}��A�_��`p���d^�Q�	?&���{�K	�Z�Xp���[
7nQ)LX�T�y4�UP���U��f���Ms[t�`'Ķ]]ً���T��p��O<�=��_��\lV�~�$���u��s�%U �Z�1|�����q(�	n��%3�k�i��|��Z潥%�ƽ ������~����-U���N����ʗ�P"�p��!UD(W3�,�v���Z�A<;7ON*�#Ɠ��xĉ,%8���)���;�VY��Z^���#
ut�y¨���h��80i`c�t�䩌���t�.'Ƹ����Bw��[&҉�Q#��m1ߴ�֯2�	o�-ř��<�L��(KG�i&}Pn.�ב�(��38>���zV�#C�>�Lh5:<���ò��}��7��&ͨade�tM6��ᥩ�ԭpY[F��|�Q�=B��}W��8h\����sU^;p�a�Yj��WAl��r�0_�c
�#0oQg�'����+�+A�J���˵���#
�*�埸1�d�ٻ�u	�-��t�� o),5J�n>�N]S�����J	���QL�'�=��bI�O�he}yǪŤs�8\:Qt0�_T�gi�z\��y�<j��
 �0��"t}%����#9oO����W�m�s����هN�zČ�1V�U8V]��2	�Qk^7��>��jQњ)%5���C8��F(����CծC�������?��27�}�'m���ͼ���T���)e����Τɚ+�P��?���'����-#���<)����yk	r��ؒ7#�KB�dU�<�؁vh�Ue��_�-���@t�Pb!�m���QM��j�
3��;�Rw#�C4�mje��7'�l:��9n&�3R�vL﷠���3�!vP�2[��w�DJ�O����[��b��MS�T�j̿�ū.V'����@�P/ڟ�j۵�YU
�fS
,Z��C�Jzp�q���x�Agd ,�0f�0�B��]�/i�`lT�gY���;0���Q��ԝ�IR�b�4���\G�z��7��(�v��?b�Ƙ�>϶��d#/�z������W�ID鲗�0�����!�ΐ��4��v�)��ngq��pHHI�H	����_9����|�͢	*8��齳������JQ��P��f�W)q��K��u�Y-�ü�;��%h}�÷#dR�B���_�+6�=,ȿ���K8���F*��p=K��h����|e%J�(�c/�8��|�׏:0ȯ��B���0Kl��0�4l�����-a��I� 3_�i�9:#����K�x����[�ԟ&��x�EJ�Ƒ&?�?��X��T�\��'s��������s/P̣�{��b��[������h�u Mm�u���=F�Zނb��G�>�s/<-j�6ON�b}��/C��Ag��Ux\@�3��6�Z'�F�j��*ZPm��^�\@L22#�)(��C<<\_�MB���,G�W��0w  ?�c�Q*A ��2-Iɒ��"A�>�l`R�`~':e�ى7Y��JiC1,�$��3�P<�I�%����9�G:�I��l�o�p7���삞�F�8.�Vj���Vw�0�~���ÏK_��|�D$y������,�
ƈ��7"*~ّ�큭S@eb	��ƚ��G�9/��Z�*�6x��	{=��D|��u/�Z)� �<`DU+)�d�oxE�Q��LǧCQQ޲a��%V��
t�Y��g���V|d��"�}u��:j�����.o��E��p���������d�Q3^H��Jv��ѯ��^L�^.����we@���ݮ�hSo�J�\VZC��s�6��k��^��i�G��1�O}�ķ�2K�������s�P�hN4%��y�h� ��3Ž��(�פ�+�K��H]�ݒҍ,
��X���gz�O���Se���-X$?�( �}M&���-V��l.K5E>��2�����
��p]i����#f�б���O�f�k�����;�����W�P��G�#�p�}�a�'m1���-���3��E�s�9��r.!t=���xl��6emk5�6�R���z�4BO x>kP����8��ņ?s�?�V�2C�R��K_H��.��	�^�jJ�_�P��%��T�̱�i��fRc��VB`�K�� H��'� Ӄ�4�)@��8׫E��;�1���B!��k�f�:���ѐQ��O��p���}���r ���7�ˍ�}��������<��(<��'7�Q��T=��룵'���vl��
�UV�h���m�!g�V�ȕFS�Q��C�̢f`t���B�y�S�*)�*d�l��L
g�a��G������J'�H�:�V� $q���-��Jl,%�Qeux���H5��雛i������	d��Ϊ~����M���VV=Xk���Rl��s���v,�N�fzG�w��@�"��q���=p�I�:6^�(��X�˹ ��+X2��s���Y��==��[z�b�.<E��P�o�LP�&����(|��9~v�^j�#:��oY��%������`/H0���a�����{��t��	`�d$� \��%�����I���Y�,u���E���	�-�_�4�^�h}��L	nF�S'�2~3��K���ӌ��h�:Ncr�\�S"!&O�1���6���V�R2�\�a��=��<��P�as��-I����KvN��7��������ږ9�L��9\]���7���8k7|r��"E�γ��u>�1_����B�
�i���{D��=���r�y�L|��׈$�4C't+t^�JA�LX��[7#��c9ϋ���*g0|�w�()ouDw�Pض�!��1�
Qls�������z�/-8�g9TT�9&���z�r+T��oC�<Qi��)ÛJ�F��0���t6�x
�_��V��?

��l��S����Z-����kI��=T7Ь������ ���pHJfw#�˯����l��RnQ L�'�"VM��:_�����p�&d�͊��@w���pgk��M�ʻ�v��,���oA�;өK{�~XҎ��ˀ��� ^��^�X<��N.��$��b0$Z�_�09�uw������%��?N='a��g�_h��*]?�����5���7l�}ڧt�h�]�4ٌ���8?�{	��%E�Z��션��:��Ow�i����0$|���[(%�i�_����P��>K��z��c�چbY�wP�d�t�`6��kZx3�.8\t_��W\ �٥��G�Rh�%mI8�`i���5O�ut@v�z��
}4��Pr�����|s�~Ój��Vm��}Q��K�VflG��M�-	��7�ݩ���6"�/�װ=Q��#�M����zmխR
�J�ĀƣT �U�� m�����2���������É����W܏��a ��4�x��,|�H:��6�M	�e