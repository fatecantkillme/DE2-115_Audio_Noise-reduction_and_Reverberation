��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<��魁�7��ѡ<5wC��)�i�N�o(���~���R�ې��U����"k��4Y �l���r��"�;ق-����� V�O��L��o�^��C�;Y��=_���r�E�,Z�0So\��iP�I�?#�"���~�u�\[㜑��6
Q�z�T�G����}U�k՞���+Xcw�p�����!&�?��(>��� ��o���P^1�N]�e������o����H�ȉ ;�G|*�=�����Q�W��u�����/�6t��Q��2K�ψ�=;[�tz������kf�ͺtp߼��gl�N`ǚ�u�0U�͆�b�s�2ȅ���z�)7r�B���@n��ڃ�`�����<��?���I]��R�@l��Vz,�:��F0������?\q�u�͸�EcJW �9%T)�̹��(�!Kk��^��[.ށp5�[���V������Q(����R�\}���:�VR&)C��bc�a�e�����t��uڶ��K��]��K�T����K�����������+T���B��=�:=w��ɓ�p��с�Z7�0���k4����c��膱)&
T} BOwv�s��X"`����Ѹ��&�0^���W�c�`��`Y�X��3�B*��g*�K�U�J��:P�"��P����$-l~~�98����1s�*
�.L�a�P���<�S��m/�� 3xڟ��0
����-o'���o, �T��n���$F��w����D="���>����1f0pF��z�+���&���qd�1k�χ��7����~�w��&��7A�������c6�M�����,<!�/n��(G-�Ԃ�,٫Y��f��a	�w-(@��������ҥ��9�P��X)�8��o�`�+�E+FTqƵ$���|O\Z����m�E������a�����z��U�-�M�_�]��_φ��Ze,����|�K����Gi�j��I��ЮrC�y�h�U�S����D&fR����o;~��l=	�Vj�d��Bo*����g���;%�2����8�a��ɳ��懥7`����u�l>|��K���bM���� �u>��T�E$7/�� w�-p�s[@Q�d�
�d�*�j����[ʥoe� �E������7��EX�&��I�6`*��p�9X�;�E��zr���-m������K���vbO�b��;�*
�yY��;=�Y�F�8�Vw�8��To�.�7������m��$�Wz3�-E�9���%�}��a��41��;������!#=]lx��[�1Nt<�Պt���Q��ɛ�Fs��