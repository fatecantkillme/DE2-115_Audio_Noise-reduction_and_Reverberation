��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<�\5e�)��t�`P^k��!j�X'^O���w��)���^�=�G�\�ѧ���zmk��$��s|:�n\�'�K:ξW(����&��4�>r���`������	��N�A�ˡ$����t��<���Ā8>܏(xVRi�b��]9[D�,�+{a��l���S]���Ƒ�L9Zڰ��Օ�I��)���{xX�J.nc���Vl�q�X�#:��W��K��6����^�{��^;w&��o�.D�>���f("���l𮁩�|� ʡJ�䏎��)��:��M��J�ҫ2'zP�� �o�c���pK����':�T���@:}�U$��0�Dl�m���6�܏/�|���',"�R�;hR�����U�VX�VO! 7���n�mP9���D�on=�E�}��٭���֧�!���k��6j�ż�5�d�E��BN8�����B>�$�IV��.�Xs |�/����t8����e�����J۴��:����]CTQ��J�h��.�#��A^�[�6�=�N{}HA-as�Vߴ��X���l�;⛈wj0<I@Mp{�AE�XF>jN��������Y�R�z֫��q_)܀F��������H�����KW_�����!�(`7l�k�6�<�͐�֑�(���Jgy<�MI�%:n���x�Hfˏ5��f��@f�bYt3�o�WI��8�l��� =v�q���K�5?y�E+���Z�����o�qsN��"&TӨ$���qN�;��E�=����g�Ϡpl�G���R70p��9��b=�^i<o�8�����u�-��3�I��b(�c��'ejXܧ����]��pBe�����0����m�N�!�g��~L�wz��ۊ��m�XΌ**���R���i�{�'߹6ؙ�N<&������<��,p�����g8�raFO��<��9�A��+���Ù���0O��p���N�'�Fh_���t.�@���o7J�F�u�B�1'zX�1��}Xr��(7lpZ�6�7;4����y8jERl�V� @�H`�%�h`w��i<Q�]ô:������Cw6�Ԛ���l{�D�M8"�|�_��oquH� )�-��KˊR&;(`�k��N.�F 4�}�H]�4�Ҩ�i���p��i�g�Dɔ'�Ԉ�ۄ#��QJ�oR����S���3}j�����w#���ooލ;��wVpZ�W��l��z�:�y=����T�Rx���RO�Y�>-��6�i�������-�^�ԅ~��u)kO��=��H�}B�t,��<պ�2d�k����Y��v��w�Fg���Ϋ#��r6��yJ��G_������榸�e�y��h[zu���T��.b�+̰��EOR�0L%��o\���
Ĩ���lT���,�G��BE�`ĈQ�xKhtf�#f���Kѽ��P4��4~6$;��=E��|�Ҁ�BV�>8���1Bcm�o�iݒ�4d!�a�h*Zo�泚^�'spc`���lhy�d�r��R�ޞ�㙵�;'��6A��T;�ݾKUV�GPS����px��+�*'�vN^R����~���G�l>ܻ��[*싣�;Y\]���\XnlB!�W�C�c*E`9�17-
R��Q��2���f�;h�9���"+K��F�XY�K�֞�i�������ƥ}�ο�e/E���{uP�2�mf��y��> �v�U�v@Q��P37$�*��OeYz���qY����:J��0
��P$�1�?�X{b+�W.Z�t=C���ޅV+6�K�����G�1I��OaL�KL�EO���n��c�0���p��J�
� �͙B�����%��|X7� �_M&B:�j��AK�)W�NA�0�;�����6r�|5�B��Av��!l�"�0F^�����%�X��G
{q����3܊!�1꯹�S ż�I�����m'6�2�
��\��<eT|d[���9�{���R-À1I�k�~�\l[�wr١�*�G����W!Ip8N�q�9:N3���^0��ۖ�~y���:7u�Ja&P}��:�f�#��
%�<�P
�M�pT���`��J����v;��$���_�Z9/s,/�WA��0��N~C�]���B���c�<�#��	aHl�n�2{��Q�g��1x��@w�û����ӥ{��K=P~/��o�dc�2[.�@����A��D��O9�^3��
(,�Ւ@�غ��[z*����[c�eGo�蠀��,���f��q�$��7T�;�sE.b([��늴���L�ylp�x8T�Tx*�m_�&o�ˈ�4YVق�J���%ea2-Ц$|^Fd�6x�ó�)��Tf�?2�$Ja��Q�G�S��������������a���g��� �r�e,V��4KK-��<�7�]��x������~�kV��?���
�w|�~��NJ8xŋh�ϣ����`[�@N��'{�z��J�F��S<��6�:���B��:��a��Y�W�����D7��o#F��暤o�a�֔���|�.�AX7 �����P�TI�I��ۗeRȐD$�퉫3=D�Q��yU�ĸ;
<�Avn�) ��cI����r���m�PCE����Wस�{�\������v'ô�_p�#����Ӌ�_Nl�v�H��~I2A�Ce�#$��l�O��l�J}�W�Ʊ)�/��S����/�>/���H��P[�|g�E���9i3I�%T�/����B˲=w�֬�ԋq��a�ɋ�0������
�5���R8FZA����f�"OGfKA����9j�r�����m�YŴK>y���֯Q��~�F�	�
�̛,t�F�p9o,���W�z�y�4�_������� �y�m�5������*9�2$`3���*\9�kݍHW��"���-�B�-Í�~:o��ip �)���� +�T<a~s�z_Nρq�>�j��w�-0"�����B?�&4��V[L�ު*Yy��~�ZZ@:��Y���`'����IY����fE��`��)��CH�j]�
*Fd`Z��˳�hTH�?i$�_��+��jn+f3�ô��bt���ŞqSh �2.Jˉ�����XQ��؏&�N8�t_X�,�4�\���|�x�w�R��(,e북ע��PX�辊B��`�Kd򶠅�]���q�j�+I�6�r��Aɒ2v]��?Ogjƚ���6����X��� "%TW���@�"B����ٮe?nr��	�ϙCr "��L���}���2��:<8����"s��P�7?�7�p�M���Q=8��a5wa����_�d�\4I��pD�$������Iz�����=�H4	_����z���m�q�~����n
��Q8R�$��ML���7f�93�&��v%��z#睥G�>��u����42^=b���L^�jᜰ��6E({��Ů��X��3��:��C񼥈˥��X�@�@&j�@�`(<�u�P2�X[ � e}9�Q�%���Kp��'�:�� u�{ްb�;<npE�~ �+������t|kW��ˏ�O��bKU��փ��%f��	zʼ5^�C�S�n�'�6:�A�xWBh�0�4PT��]�ꥷo�*�1�--a��|il�2C]XN��ш����h{6��R�繅C'K4������߮B�cUz�D�����~��+d�ٜ�e���KMc��4�����g�?�B�קlT��^��f�Z��q;Z�1�O�(�gQ��/�刟2�������ۧ�5^�9����q=��
�Te�m%��h\	�LK5@r/i�&Ыd��#�	���	�)a������Ӈ�;0��W���s�\ʈ%���]G�f����r�]���Lr��o����X1���xy��lR;��4�*��[�����aY_M�0"[!�ؖ��w̸-T�ݢ��[������aVV�x��@��ԔX��{� �aL4-|8P���[gR%�I�z��K�^�:oCg� $߶9��ݾ������&L�*E߹���m.�.n�]mBJ�[��ݮ$3��V����Il�]�
�f���Ȋ��{��ĐN�Db�\1��u�r����j�r�a��E�)2CM��}Y����L��X)��<1��D����ir�W3�����jrU���J�/j�U�㽐���N��P��RfΌĕ�C6'��XG ��pA����l��hF��a8b���;�_;�*CT���VI����`���M��B����+E�m��CW��#�4Z���Y�F�:�w'�ww�>�Y9,֦�[q��RQ%2J�AY?��my�i����r׏k�V�~,0���Q�#i��<��F@�:g!��Uw5?�{>�;��zKo�K��b\꺿��	��*���<H||29N�0�������3U�?��O�Cm*6n�cERGE����1���^����~۶�+ha�Dd�K��5�}PGL�̰�J���-D�����z�ԫ1'�5X���ԖJH����T"�_<�u��4��M�:�f���E��=��ol�t�~���ZOF��b
I%<���&��O�?&m��~g���1ь��k#ê���H�U+?B�,�y���t�>Qz�-�6�|�@�3 ��+w�yȩ�̪�c�,�A�^���I�Y�7���R����;����M]F3�/�x�G��5������b�6�%�S�X8�o��=�b��GGKi��D�>�#mjB� iI��|�B��W�5�i��Z�S��[#u���H�b̈y�+�΍���t�l�XR�ɮ#�թ��z�7�0��zo8Jk���;�,�l@*qE�=�τN ���\j��݀Ǚ\�e�_FX�-Z��I(K��w���K��!0�#�j��TO�=X��"
'�|�ð�&�`�����!�w���_q$�̓q7�z���7�婚+�]�G��h31��D|H�k�&;�]�bś�4��Q� �E7�����WtI�����lL Q�t�W��0.�9����؅��G����	�����Z~/.���sS��`N��3�y�<n�/!U|����Ѐ�/e�6)/p��_4��ؚ�MO� ��V��	\����b��n�_�+����w'��`�;Ύ��������Joqx�g��}o�O5E��i��&ʇA}�S����\��W�]mgՂsY�#2cp�r�׬$1�3� )y���ȩ�]���+���1��@o�ô-Y�z�c��a��g=�n��Z)� {����	����h�RR&&@���u&�ǎ�v���^�q�/7���,!I*ñ̙r�������N�@ݺ.�G��gP	 �[�e��p����]Wq��i���&�8u��2�5�#[ ��R�z��:��@l�*6;"	{w~� 5#�v��"H^1�4<m��q�sVy�����X�i��5(Fb�E����h�L	�^F�گ��* �x�f,d�<�N܋�øo�`���4�t
��G\���88Qc�$�䏪�A��a����E�I$ƆO^�$z�Y�����k���~Ȼq�)�׳8U�Q���C��袯p�)"V�+f�1��KP)Á�P��zd
!�Q�C[%��M�~��<?�u����_ܻ:%�"��pN��8���&�`C�-P۟Rj_$�Ps�D0ww�h������Vcړ~�|��Y���УOBK�,�D��W&�O%��oj�� g��4���]�/}c&n��U ��@�L��"���u4�9�%��b��5M3������Ʉӥ�9�P�E�ju@�hq����ۈrC��ˣ!��z�ʳQ�w��i�3De���S�@%ܹrw����4�b�N�ll��yH7��:���B�ԊCbYz��R_�k��W�9�b#Ο>�$�B�\)�%"؛��x��1ō[�l:X;��7����9fR�WѦ�:��q��_�NmSՇ�rH�ǘ&*V�(!�L�ܕ�$��X�+��E��'85P�{3G�f=w	��w�J��5IDwv���=�:e[;�U��,���a@ݮ�,��S�M�2��h&[-��'s7�-%�כ�9o�X;G���>�dgIّhWR��Щ�����g��g�Ì����@�=n��}7�4ְ5a��f�Np�6|Ewl}�H+r2�x̂��NY�x]fgd�-���
���zB�.xd�C�Cr�+�!�?��-&��y��6'�b B⣌�ƅ��t�թ�,�|v��-��JdE�9�4�t}��U5�Ǖ�M�I��A�յ��T�Z��PA��ݶUe��qHϵb�V�G�N$���v��Ǹ�T�q�5`O߸�l�S?�O����&�j���,HuC.��4�O����5\�c���D5;��`��B:
��?#͡➎�GTu���-�sO��(�N��vTY�K�lh^�g 	N^�o��0F꽨i�Ε~@�ʒ��A���<��<�Z>��#L!E՟|r��fy��~�mĮ�>�%�"\�K��2Fz�{l����8�j�U�X��LX*@��Ŏۦ������l~��|�����������/M�������
؃ɬ�dk����-� ��"�C�,Xq�wN6���7���<Q�;�V��e����;r��6U��})qn�t/v��棚q�v�D�y��]���� v��FJ���ZP�6���w�cɧ�`����v�u~�dD��6��^��0pLHM�]�W�#�?�����&������T�J=�9�C�OV��7͐��s&F���k���JjEһ�[�͇o��Z(x�W��n� e^�W�}�0#O������Y��ʙ���z�_���Ϭ�@����u�>W�uTe-O�L��&M�7�|,�LG*!<�Ym��e�)x�����z���: ����E�T-�pC w�L���wx�oh;��^�P)����G�-��;~�ӽIo����2,�4>/��(:(L�5"m��AQJDM���X�˱����G砳"�#G�
b�D�4@w
��\�9˫j�w`���|���r��'l��|�5uo�:�1�) }j�qO�O����t(�a��>����t9�$(�����c�R��iB ����}~,�7b�刚��J.�4��f�H�=�"�}�+H�o��P�k�Z�B�D��t�^�'xIgaF���MŦ�Z�	B�jUژ#��� ��4}^-� s4�eSģ	����w{{@^�n�%�z,��X�F.��d�t
��Ĥ"5Z�![~�N�v3�3#K�?�s��;&.�g�p�#�,Izb^�C���\ {?J~�O����Ցu�[e墦`���J�̌T�ue��6V]oo�ߝo>�����_p����b2�}W�)�V��<�*Ǒ��ăt,D��c}�L=�9J/s9o@;����(A'=ٛZ�=9���!l��fHHn3���������	~��ٶ��[�.��L����9a�*�?���3\�T�W��pGM�����àA���uZz4�UGs���,%c���IP:��a\9{b(�馶�-�\�m���I�2�)�n(�\�ua.�c!��[�xEE���W)�Xĵh�����Grof�eTƜ戀~�O!x�,��(�Ul*�&��٧ʏNEg�/I�B���mE#��TP���,�זR*�k7Wf3�o��P�TmcU�[L\�zel2��◼�U]ܗd��势
��$�)��a�/V7�"֏;}	����i��G�J�Anv�0�0����-6_���>�Ԧ];Fp�����܄�zwM�X'J;_mG��^���><`l��!�G�j�j�x�z��J�B���U�ŕ��z�eE_��z��	~���cߗNl�V����S�33�Q�S��K�2�\�	�L94g=rF�� W7��C)�K�7�َAǖ���k���6Q�Q���&�u�b��v�d
�}�ͬ���cj�ڗ�V?����>��O��5��W �;o-�+��,
IH	Tw������%2.e{�O�%n�'p���VBk/|Ϯԃ"�+ �P�N����|�����Cth_]j��T���Q  ����xmRa:�&�����V�����m�>�`M��V�jek�+�o�;u����Y7���xQ?x��TD����O�޾D�!j���c��;S�Z�Q�%X��)!դ�I������$�����?�Is�b	������f��ꮷ�~(��L"��Qt�!g)kq4T�g��jܤ�X�K	���z����_�O���5n�%a����W��5�,6;��_i�G�SG��ŷ��5��Q7M��Λ��%����<��o�H��oV[��R'>��Y-<�h�����i��(a� ����h��qN�bꄘھ�����6�P�9'����:���:��#x^iM�a�ѳn?�jl���=/�z���ч�Z�( ��AC�s��C�ޒf�G7��j��4Jȷ6��.0�Y�xuok>�(��g�ዂD������J���*a�#zs��D�!� q�.�	����h�LJ}�ğ��a����3
-�s�"�k@ө�̯�k���dܹ3i۠�Hf%8=:hͯz4Լ��������/�F"z�����U��%Z�9���{�Y�ʺ���I�@�Jl�7�����^���70I��/E�d�m�@mϔו�KP����s�fs�uSHV� !׃ny�-�<X>��<�*#���YT�&'�����:���F�T�+j;�S�H���,�u�#j{h(f�CM�c=J_֤���R晉�jI�؍Wɝނ�NM1?��afl댝ʻP�p����ʹ��_js�t�*Mj�P8�t�GR��e\%�#85�/��aN77
a��,G/lm	:�l��l�D��˲b���Fݔ�u"��ݻc��X�s��d[�?���%gʾT���FҎt�uWb�ϙ���>*�t���p��-;�Z$$=��Q� ��&F�C,0����t�wR�2`�R�aW(&b�廴��~hȦH�Ώ��J8�n�U�E���֯Q�R�)��7r�f�	k&x���H+亁39A1h�y��Z���Ĵ�ݘ]e���K��I@ҡ��p�&��ј���*Cxs�S�g�+�*�)z<�A$ZK֣y��,
�Gb�g88�u4�
��*������t��]�|*����8u�\����bv?6��$ir�,�UJ�q]�J�/�g�~aANlN���q٘�s%�������w؄4\�o��Ј]4� ��mqH��#T���N�>���.�k'��`��d���4��k����n��[��텓Y�V��OY�7C�[��Y�7�k��R��2�]#��xUv�$���C*����c���.4����`����͕0؛HO�Zox�.ؕ���%�]�JZ����0u�Xe9j�%�['
�-^���f��}���nB^jw�ma��WkݷbB<uK<�_=��9�����/u�}m�|�S�v[33mL`a�h�X�|3�i��~��p	����@�Q4 ��]NR��#B��E���&�����*X���%��mo_�w����ւ�� Wn���i ���3�E6�:'����A���9%�����?܀(pܧ���d��U��F�0�i�<������� ���U��"��]u(�=Md��fD3�_'p?G�Ӱ�{!Ry�D��c����g�l�`s!�
mn3��`���Y�v��ʕC����]��߿$�tC%랂<�:歓�����?q��Gͷ��)@��&�;Rk���H�0�Er��0���>v��/ѝV��Pz/�՜Gv-w�\s���q������=^��/��(�Y�6���~75�\���O��)��!Չ�e�5Dcx���䧕f e�����;�*�iLs��3!9�����<�
��*{���@�e���כqL�'}�e�*�[�����N��uA���������C.ެ賭LF��@\Ӥl�<y��G�]�:w�%�?��ؤV)uAN���3��^q?���|1¨�v�6���W{2�W[u��D�eɓ~<и")9�2g~��\���Yz%;�˕	�܃?G��UN�l�?�3���)�%�Jk�=t{���<,��+�-s���~�q�Q�>����s���:��d��]gpO�	�������L2�B()ؘ�2�B�y6'�y����2�nww���/"�$�ܮZr4�Y����� ?�� 2�آ<q�2��7�����*��)��^�h3xd�<e��͔������"�F���9� o�����r�FCD��/�hb�Q�c��*�\�;)95C�c����#.��!�"�n�h�]��n��)�S̆%��d��{pu����:[�Ӛ>vFF�[p3��l��z����DTK_ �[�n�Y�G���՝ c/��F;0q]��p/����M���|��|2F�`X��-��NY�أ�#�7�?��x�~E2B�[ya�E��	g�l�o���b����f�`��b�����|M�U�򯀅�My��z�)��o?y�5�t� ���:��#2���j�Z$>� �_�@�%p5o��/į��x<�ɣ�ىc���D�N����{b�
8�8-�+��T�ibj�I�����;���{��I��Z��9�C��U�j�U�<22�M��]L)�����1:��w��4Q N�g׷��A�8g 3n��ʤ��Љ�W�������k����`�%	Oh��p^Gg~��x٪:A 
�_�h٭*9X�SÍ�tOa�$(�#��(^�����8Q��Is%�XȻj��Ղ���pH��x����vmS(�'��]��|=֤,#��(h�)�6�`�z X��i�����JV���F�jNl���K,�������o���G3(�Sr�3��$�R�������+彼ɿ���/ ۋ��2K7�qN�3]�LV>�����&Z���a�/�c�Ww�/5`Uu*��3��+����(e��!i/.��UZ$��4!��� �C�pB��䏏�A%,M��($��i�/h��3L����vi�l|�o��E��Q�piJ���B�O��̂R���{�V#��y˧ .D�m�����u���9u��1�cG	H�L��MS5��1��a�å%�]�cp��*��\g�o�ɚ7G���[�|&�gH�kV������1�އ��U�\�h^�%����X�O������Ʃ�9\m��٘�_�$1!�^��}6������վct��?|vL��|Zvr�s�����9��M��|϶�W��Y1���D���o+0(C�7x�X�~��� xCL��fv��ǆ`ی��!� t�h�r�j��Ej�`'hR�1����$��];l&�7���<��������aX�-e��G7�ӥ������%*�y�dt�����c�2�e��T�u��Z ��ɗ�6)��ND��&�ܾ�%��ڬ�,���f2�)?���%�sW��T|�+Qs1�<���h�)�5��m��.h��^�~G3��U\��vr���~�pZ�2�Q"3�'A��*����l 0��#o柍�¤�?��T$�akB���z�� Oe��8V�|_�E��z}��9���M��̦B>�b-$pU�����^W�Nk���S�0�ݗ������wG�W���'2�
>��T8��~?��sA^Y����rZ���!�J�3�a�0��/pŜ�\��M*KIe~b������ҥ����1DD�Y+?t�"G�j���D��;�r��y���t'8zH.�Apb��`3��&�y�po�ZtO�R�������[���N�ZnWrL1�qV���Վ��1�:+��U�L� `�AX��jP��c-�*oӣ9��7_���E���U��)ŠMW���z�������7���O|*�����è�=с�8p8��9����M���2b�j.~�m�5V���$�̪��g���m�S^��\����M�� c�.�zbM�ךP��=^v�����LϏ	6|g+�t��;<'��D��P�&_�t��9۱�5�$�SvXE� �4��A�E�]�������s����z���r=\�Uħ/�BE��?�Ù��R�m5�S��E�y�c�vRE9?K)x��ĳɴ#j�S�I.Z�kIXKo��y�-.���R�����ZԼ(��!Ad(��2J~�#(c��!��W�W'��uߏ�Ʈ���Ӆ��5�۫�b�!窤S��*���>M��X�����q�5�]��b���aC�'��ڽ[���H� 7�F��h���hlK�����ť��Ilgw��m�Ӗ����i�'ʛ�g�Et���!it�;K�=_3V��-}���y�Ko�F{�޼z�^7�WU�)4��	o�hMM�W�S23�P���)^����NA��e��8�m.����`�v�%XQ���q���N	��$�s*:������ǒ)�!&q��C�����Z�,O9�<����o��8��J�e��e�suh��#]mD��+��/"9�@_�Z��EQR�s�#�뙞Pn�{��h_'�_8��;�}�曼ME�іRv��~�4
��%�;��,�v]K���Ψ�����
�?9c�,H�H�$�[S�ni�D�`�p	A�"��fYu�I�h-J�I�X��du���.�߉�o���r���2��j�@ "�	9B�o���J��ԋeϠ��L�|�s0SA?����Q2:J�[��hN�pi��)��A���0�oi�.�����4���72%�|����cKm���Rs��85�ؑXǴ��������_B7�����t��Ʌذ��r#��ٙ�b��L��D����l�r.���o�J�n:�7�P��>
��O�:J��J�H׷^�t������ۋ�O�z͓ܚ ��b��$<��&rJ:L�F��n��q^qz���� a��V�ضB�XЬ麟C������ȷ���riz~Qozf8� �<]U��/�K�N�?�g�-iO�$�	<z�����s��Lz���Q��Wfo�L�Ͳ=�ymu(p�q�����R���@����*����ʝ[;V��dh�P(u��[��� ���v��#g����M|xIh���M���/���R�]P�q��ɑj�v]�&#�e�<�wz����Q�2�w�u�B</N�h,��[�p/���Έ����6�~9P	X!�r��Be&)�������4]B��Yê�g&#f�����rX���ˉ��H�X�I��K�;ZUTuOe*����i��1��6�Y���s��'W�=���}X8u?Y8I����[�a��X��������0g�U�Ǘ�yN {�\b+�dӦ���J����n�;��3L+�rq�yj[6�{�g��=ȸHU?�W�<��Q����dE��Ϗ���hJR�MXg������og3@=Q� ����?��5p(|��TD~�t+V�h�W� 9g�V���&#<��f܏4��&g�QU�ֺ98h
���F7����E��X"���}4�=0Q�Ʒk�uXaj�~NY`07!��)�PO�O��\ClB�\8�N�q�9񓗑I�r���'�X�aÊ����|cy�k���
�ɉ~���H_ߓ�� ejݳ�+Έ�O$��F|H�fy�4>\eeе��5� ��tjRV���=�I ^�O�-&2��A�S����	A�dK7�t]af5�pț��������=�����a:��hG��O�r�@U��^�A������!�:�{�=���y�A~óBA�QD��,8������ƿ62<�BpcY����V�� d�m	,7n��U.�M�T�Eiw�D�N&/R��Eod%�.�Ts�'ྈ�x�N^�P9�Ï�����V�6��6�<U��������g�����aШ٦�Ke��"�;u���q��0MA�����p���Ho��;|��}���.��C�s�W����3�r0	ݨ�uxX˱�v8��y��_vqOf�F��[��4)R�������ñ�T-TĚ{iܥp�
>K�б��.��rN?i���y�B,�-���[�����	J��Q�£�z!����D���Y���X}j�_�9F�(dc��?�-���ڕ�zZ�n�h*��F1d���46�Y,26;��-&Q��zE��e�	iX+H@�w��3`h�f���g����P��dO�E���-����*~"��}���\K��}�ќۼ#/�@�S�C�:՝�����͸�e���S�aB�� =;��7m�N�=,��W�LQ#�7&	�3/���f����xF����n��~U䑠;��gDGy�w��J��0	���L���gf^R���7vq� Jp0�m[7�ٯ@� Z�XD�z�2:�4z�o�.-�up�#�����JJ�{�6�]�@]^*F�Q�]�s�ƯkǣR>����{��)���w��XA�G]Ѳ���tz۪��cw�}&�l��Al�oM��U��������%�l�\�O�!�UKiIA33s�P��W��"w�}}���2�.g�L��z�'{@Wv��	�^=�A��X�^����d��>��}0>�^���%���ږ���p��|�'�^����׌G~VRܻ��������#��Kw,+ڼnG�x���тx�XY.�x5�������F�����w�z���K1����숖��zkL�Lk��J�}�a��
^wj�+�H�|~p�,"���yF��4�W�/b��>�Oz�G_Q���*�� S���~����ֳHa��Po� ������_y�湮4"y\��Q<r�@R�I=���S�2�@����I7��Co�k����Ę��������q�f�o^��UC�K��z���*G�1�Z_/�C�m��G	���<�91��@Tּ?'�j<Aa�ҸM��J* F�h�(�[�٘�S�:�� ���}���sɌ�iגOĠKg�,�}�w|Ż�%��8�2��T���Uf4avA����t�����c�&��|�]�>�N�ዠ�p�������_�9��Y�յy�Q���;¯ˆ���9�.�7E����:>P�>�U�9h?��칩1������WԿI��w�<�`ˮ�^W�V�v��3+���^�7hHj���k�#�Q�3fhId�Ƒ�dV�y*�IoHU�bA�|=ռ�D?�ܚ���x���#�%���b&#�w�i���,����S�{�OҎ��O���O1�=��5�r��o���n>fY���Av��o���o��,h�25���Oα�6'5�6�	�t���� ��$�Gh�_[��D�b��an�U�1�(1��>`�;ӳ֝C���d9ʽY����W���A?/��%)-�Uw��qt��*��=�K�V�	PD˿���#�I0���������4$0�o
��U�'E^�~��y��=�F�!�jI*zNV�mqj�,�\�C�&0z�)'}�sy�\���׌3;��a�BZ2B�c�s�L��b�7���z��$�۹�gk�8�67��C�2��������X�uP6�7����Б-�f
�.�2���{k�H����ZVp9���^/{�}."Ҟic�@G�N~�M:��i���p����[�\2��U��	HOb;g�y6���/�;r�7��4��=8�uR�35�'ٚiR����g,�6�j�V}^���U����&$W@�0�+{�!������
��62j���9�
pZ?�l�T�CBoM��?���6������	FJA`{7�/-l[�{�~�|�{�8���͸��m����}r�C1��[7�;������ɮ4����7�
L���}'jSb���"�Qo�\5�q"J�dqu/z��^�����H
��/�
�0kT79`�I*H�y85<:��B� ����W���0xݭ�$�Q�l���W7�i��ʘ;m0K����mhPl&��hy�V$�Խ�WLMp�"E�*,�-������,.�_NE��K���pkQd����Ƅ��i��_��=��!6�u)�Ӹ����r~�-���,���ز`x�,y�Y9^�'i��/|��8@T�K�]�|��FN`>95p�Y��x�M��ef�%=U`��B��rS�|{���(�9?�k�
�A�K�*Vc��2%����LHh��-S�SW^_�He�"���Y+ɳt��S֎4��'H���������8���
� E�]��aJ�c����X�������ZAo��ENs�n��6�3�]���%��Kd:f��u�����ll�HE���u�hxG�ݕ#)�m��G��v��Kk����'q'Cx-�zE*yE���[�ҝ�?�@,_�Yf�����-�S��u�)�ݴ(9go��x��+<<�,_*��X&��7FX��k�>�a�&�������{M^��G�������B��_���%��&ν��Ş�ד鄂/"LoX��2D~�i�p墠� hY$�,�����p�M�ju^�i~L�P�Gk��QEUȕ��)@�_�m�<Ŕ���Y�����qb��/hk�h�Y�A6ő?�Y[M)-���,_�z��՟���/��w��ү�M��c���C��u�UK3�b!`�ɩ��'�P`�C�v�9]�@q�{�똒���D��,�^ú�il�@^4�#+�u?+��r~��eO��.��Ae[~�n)	��)*�0���`)��tm�U��MW�j�9pDÔD;�`Lx��'��Kw��(U|=�tz�h��m�(��/mb��]�����^�df�Q�oU�0&q]_�b�����~*�ktC�:�*
��&S���/��u��]v7i^��/^�~L����0�-�8��}�8����=/p,n���{�PTFK�Ho��L�D�̩�.�6�%�1)t-Ч�t��z�_���5���m6Ov/��VԼ�b��J!M�ʓ�e�����`��twY*�?�H�� 1f�ne���m��yPD:�!��i��8��&���}n5)e)q�^�)?���M@���G��b��R4$�:m����̉Ч�]Ͷ�gr~A�0\Fm-��̑w���x����
T|���9Y�T��f'�Ӕ��9_������LML�f��֔[����J���I�W��-l[�±�!S���������:4X�/�2M�cj�*-?Hg/+6M�5d[�I��5\�o�` �,�G���q��꣮r@�ǽ;b�I�U���0ܗ+8��<���e����m+�~�����&�԰��ͭ>�+�9���e+.�?[�K�/& �IK�Q�N�<��|���tI4� UPA���~f�܉��@�Fܴ���,�8��Ѐ~�8Q"g���x1��I0&�PIb�w�[��n��0���2s,�K{�`�͢�,Z��oeXL$��eE	G�|� WsC�g�M=8���	�/��A�_x���ho���lw� ��{)�G8�/o1�2p�9�VU��Z_)!��&�[P�Xc���B�<Ɨ%�eKެ�`����f	VmÏ@l�N~�QS\G�=.��޳����-�s�����_��T���=L�a��e�Mz�c�6�7>k��Ǟ� �V`��&��Z�_���[�A��ڱ��z��A��8�al��W�|���э��u��0hV�I�U�ml�*8�5�U8x�r[w�p�ݙ���~�Đ��P�hY�l�]�0����칰�x��<舮(�uL|�/hx<�dCL�/�� �yiϚF2N�P��lҐ�y^��D�
-�S5�d�%�Á���8`P��������͚ͣ?��==�rt�na��V�nN��f4���*%0#��`�Q��;�2��N�<"۷�Z��DHd�-��h� M�@�}���q�v9�%Pv7�%]��^\E��� �}n��M=fg$��9#��AER�?`C�2,9F�}�^ݴ$tΓM<Њ��� Ke1��r�C��~�(%˘�`>��T����2��۸Q�w������.�j��G�ʎ ���A���������5&0���x�St
�WG/Ct�t W��Am*϶�n���(��T�-^��&� �ǥȘ����`�ٵ�'�I�cP���q5��T�W��D��>)-��6�=�ʶȎ�;+qw�YY�^�$^�ki� co#h������E�<EEW2k>&'���cx�"W�}��lz�����5�����yzPa�m�w��J�k[f�b�}(6�gZ���d?kVK����/e�׹C��`��y�0�����T)�>v�v��d���jR	��E�l�rto��B���T`�o��̗͚"^�B�+���Hao�h>���|��Z.��60�Flt�h��G�W�Յ��,�H�I�{rg���o,���#�������!N�x��v5�J�z"�w�������j]�� q�Ѭ�oQ�C�mge�y
�*-wF�����"�Ds����j�ܽt=/�O����gk�����L	�n��˕��k�Z]�	�������������m�и���T��qUAQ1d����C��ֳ��B����Fј���(�P1�Q��5 �"W���6X�R�+V�`@I�	�c+	3̚T���?ʽ3!��}�9�J=��k2�;!�(�*��~�����$����
��:f��>��U焳P��u���n���q�N 	��L~R�E��l7?%|��z�g��_�rSV�����"�Z�E��h�٨�4���)P��X߾ŏ|��	G��#��lcz�f�_��4�CEv݈���X�㦆�*tǸ�s�9W��'���{��.T8�|Y%�_D��<�h����"�v/�u<��*o�ɀ��"zEa�	gl��|X��!��ˬ��X�PX2��v<�)����p�;%i_g�w݆G���W��V�#��uϺgb	8p~r1��"݃��u�N�$�H'�)���4裎�5�$��)�'i������LӚ'���8"v��Qp���*dH?����I1	�M�񹂠Q���G���2���3@@r������[����q��=�r}W��㼘q&|��fڤ�������챛ᰥ4�޶gi,56���>0jT<	�6��;u�&�h�L�J4Έ��Ud�Њ �rp�����Y&t��Z�H�b�Y%��4��`�:@�Ȩ�X�n�}f向�\����Ԓ'��ZG�ʰ �ǞNYC��U���8�n��]���w�������:86��w�a�������a�x ѦD&9��G@(&�����d&7�`۝�nLN��0��u��!z�����ko�2�n !��t�!���5�h��U�Qc�}����L ��$���>r�\G'D"�����0�)T�9E:~���m�Wp�d(��|�������O!��]��9z Bw�츤�-2�-ViOԅ	Չͷ��5�
���1G�mCr1ɯ^@֒b�	���ن-@�'À���B@�N�uo��(3���(4�չ&9��jlS���N۷}�[B{)P�E��G����tO0 1c;�S5�>$�r�-hI�G�}��`��~�$��%�.��g�y���Nʲ�U�coGe3� /���������{O�~��.E�h4 �lB(4���⢩��6t�ʐn��+��M�䕎}:���gvE�_@��%%E޸���]�	�$�f{�WK�"T�����n7�� ߵd0�M	���B�g}Ć67�������!�|����@y�2���a�����g&� ��yk��!��9nFBI �%jF4H����r�����7�R����U�[@���Y�n,����~��tkXZ��ʠ%H�cK���Bk��@�rO��gꗂ�J,#C��m�"���q˖=?�wˀ���N�$U�`?�7o�R����}^E��s.ZU���\�e�o��F��k�e�ˊ.HA+>	��١$X:s�n?���:�o��C���89�!z�C0��U{Ѧ
��kVݸa����� `x�?_o�J<��@��|I o4x�|�TL�*Oژ��c�);&+���Z�d9v�ݴ���������R[����׿�H��������z�sۨ�eƙu_�l~d�b����%k��t��L��C������L__25��0q�kz�⸢�
��x�xӠ}�o�Ǥ.���;[lrz��W� &rt��p;� ���|�DY��ɛ�����}fw��
'հ��G(���߰3ky��MW*��$�尾6��r6�2�$ws���Kи��`_QwG�6����kC��%*�U�骺D?`9���.0���=aZ��6Փ7�������gƧE����jE������J����LI�=T�V����3�]��=5E���0���	Ey�,�j��4�شe������p�����oݦ�q�4�R��B2�5eB�# ҲqM9�܁v��b�6�H�s�D�C���F����h6c�QL��m���� ]es�e.0�lTq�����QxR�O�~����^��e�W��1Ա�P�A��Y*\}ozj������X�k}C���u"T&��~�'<����9j.�}�$Qс�l�6�8��4V�DHG��yR�9<|���L�B-Ѱ*��E�����_m�0M�ڽU6.�N!���:Y%	 :�Dbdv{��	�s(p�V=9�`>��|�vh���_���55���E�y�������?|�~�NI�n��4�ƛĔƚ�3(��!Y�a���DN�pJ]���oD8�7�p��2�4�	6��-n���Dt�&�^6�%W����b���mṢ�Aպ#�~fmS迃"��H���q2��{V�����s'G�n�������@=%�pY/����1e-c{����s#�[����}�(b�0�3�F�+���� \ (��I��sZ�#jB�pp�Z�f�4����j�W����|���=��H/K�����ݛ��9s`�>����b�Nr.Ӊ~7q�}4	�H�ޫ�6�V�ym{`b�}m^F �,C��=����F��sK�a&q�o�B���+����Oc.�(��2�wᣫoƈ��ح���L�bBD��y]L�x͒�"q��t��ye	�����M��9@�|��`e���Pgʨ��U��i�*E1b\E���j^�Y\(A��K���ؠȳo?�W���-�h����itl���k�+�GB��6����S!�$�qV���n�(�2OY>9����ja���m�#U
�(�/2�����_T �p6�^ܭ׃�GA=U�u�����"�ε���+��@+u�+�ec	6�R��5Uf������d�4Q��S����:���ݸ-"�MXl����mAܣ*�|�a�L��SC�ı���G*z�ab�8N�F��е�m��=}����6}�2&��"I���x�Q��>����z��+�����G�q<�`b��r��������#�YM�� 9���	x�K�&z��a��f��N�{�N+V9�s��ߴ$,�iB��A�,�7h�+�9#���<8zcXu���q3�
1�[I���9#�\w-��4���tB<i��H�<�{o��){e�@��o��M�yN�0s3�:ٸv0���� 6+�p6�>3ʉ�6s��a9D`�1B�c����&̃y�������n�e�h�ٺsf�f�_�\X&�MP�1�k��d�?�
�ȟS���Ӵ����5���5��o��ĸq���"��8���]�}��~�wR��D�����TY@T"��_j�n\�KR&�|լ�ݞ��'��1f�B��������:^���p��E|k�YP����	�������a��T�?�	�\��� �� ��8 �p��*x��!�:0\�����g���\�5�9��0�=���aL7Kc�a�����jH;�	����v�k��5@B�.���5�յ���d��ҘI�|���nJ3/�V�L�4��t���C
�L��O�]�p-�ԧS�thY�vt��[�^ t��OQM�w�k�@��L� ��jk�Ї�z���M�!�L�)Z�v�r���2)�Y�[}6�L<�ZE����&�w5�n��]\`*�:��L�-�M�(A���9�V.g�iF�zw4�W̓ МQ6@�������7w��d�<��!�9���"��O��}o�H�2(���H9咓
���)rƴz�<o�֖�0�sjY��wF���v?l-(�q�^�Z��}65�0�.�n�A� ��"T������l7Mvq{9�4��A��.�b�J�Hn������3�t���q�!��_���vH�g�>�!ǖ�2���	R��I��U@磱�%;��$ �n��a.�4(�4@w#� g͂�2o�_]�nL��_�6D��P���5��{�C�Gm� :o�Yf�K(*����{�v�;�*Dc%�� w&]
�,<�Yœ�)cQ�lW#�z�(������
ԟ����a0�>)�������i]$p#�E�"p������~�*�k�b�6���t�'�d�G0��ƌl��t���^?�@QjW$"#�\	����V��2�D��{\���m�~8�Y�IaE-��0~;%�9��zT�@��?Xn� R�xʕ��s���aj��<�L���m9~���'�E��D+�����V3r�k��_K��3������D�w�3�+�ZC�wZak���fw�փ򳉵JV}���Qo	���9fA#��޴���h5�O�tj�����[tK�� AZ��$P���u
�z���v��C5ԧ��������?r.�,ۋ|ѻ,�������8�;��	�&����.Y�N�	#���l*HM,�;	���oo �FSa.���!�XD}��xN�B~�5�t�Oc���w��L����E�K`�-8�2jXe��4�A��w�4�� ������Ѳ�kT�dw@3��s,�C.��������������vZ˅��.��6�⼅�7�%Iv9獲�A�^7��H��F���s�� ��87��ch ��Ft��pz��I�d�:İia���$��>#������[M/^*L`����໲��0�X8�cG����:�����H-H��a�j8�_�Ԉ�3*��/��	񸺳���`�"��3���hO�N߮�6��|��:��C�Qc���l���}�@ӝ�@�;��}���dݵ��KuXD��w�O��!���͝�y%x##К/q�jyȬ���C���s����6�e0Ā�3IRbJU����'q�D��� v"��x�}� 57�F+��ԌTg1�@�j�Vt�p0'x��4���ׂO�0�yݳ˴�{P�u��n*s+�]�A>���_�yBMp�1C�8�]@o٫�m��V�� z{i�I�����
K���<�d�����!vBbڪ^"����4��
����.�BF5���<��1n)3e$cP�Q��\��-�T6f���J��e�G��΢v������ȫ�g¾���f��hkD�R?2��!�� �:��kQ�)=�=)����d���(r�B���k6S_H�59��T���l6�lȥ@�g )o0	��mKW�����������鎁��C{-n7+����r9|Chpbbje��Sї8�S0j5z�`�P8�l�L���j�V�:��#a�xS��=�+�{�q�Q��ݧ4�d=��&�>KZ��Z]�iC��̤� ��Z۞��]�C�p�)�-\���f�V���)�DA�_�'B.�d#*���2;j�/�磂�o�Sζͅ_i�#Y�Bk�T�])�.%������X�˫;�~Q��@Q�hN�c$�f�����`3�J�x~?���F�38z鎕#.Í�:��Po�
�N�P	�O@(d��X9�����b:��K���7~�Ԇ�q���
��7��˰l����K��[H����m��$�|����A��g��8���$��j;u�|v�_����=���!�'�Z�����v���'�K��ñ_����n�3�$��"+Z��LM�wk='�^p����&tJ�ţEokk�u�<V�K$������?g��y�2U�=��&i|��eF����yO�dD��ն޳G4�*�Fz������ē9E�7�oDf]�xD��
��K�8Ô��N�&xpOZ��Ar���N���z��R��oGP��/��EL��1I�c�����HTh��B� �x�>���E궏♑��ײ�N��D@��Z���S�X��'n��!���%n�N��ܣ9��Ӆ����Ƣ�p<;铢�*���"ͨH� ��⁞�'���(N�S�ݼv�k"̟y�>(@7!Y]H��v��Cƻ�nN�q]��#�U�BTxV����ߡ%ӡ��LO�(�ԝYv�J݃����LI<�,ɨ��ԉ�@]��P����Oq�f�
ku�6H���9�D^�mA��&�+���}N�����i�H���.�?b{�����i�lK�c#��M�����)�m��|�Լx��Q�de��E�b74��J�Þ�c:�*��B����IR&���zML�Y��F�PO�T��C��[B���?�&{=�{��:�v�h���$!�y��]v�QF�4�_��h�ģ�6�
���M�
ql���O;����?.Lۀ���	��|�>)e^��*w�/k8i�ޙ�B��ǽ+�k���~'�,���I> ���$�X2��Sis�m���p>��s&\�I����(&� 	��ap�c�(s ;5�f�4e �R�mJXg X��]o��ۖ�Y�����Rq�Q�$�qʥ���![ *29"�̎<�2lh�b6���������\j��?��ٔ���zN�?)�g�\����oʗF��,�<@����.��c��N4���@\/p�`����>W����ߦ}3��$��Ƅ��D�k��Z�E���Ch�f��ݔ����j.���N��a,ܜ��h��g��!Ͻ��@�k9D[靃��D|�~K9�9�5C�gF��v}א�)mF���u�G��s~1�4 W ����0�G{� ��WC[�﬘�$0\˔� 
p(�����b"d��B�$�A�G�X�� Q�ż�N���]w�r4�p��~ 6V�o�!�����DV��<>f��2�|�'"���f�a����T��i`
DZKim>��ϾAQ�I��(�Hݡ)���S,�>�֛��+;N��
�0��;�=sPU%W,!�~��-����*ب�����(�����Q�~���	�ҺXZ�8ۄw)6(��j��63i�PG��]��sD�[̠��@�F�P`�H�j�;,���b����|]��9�+���bo^V��5�cU0�K����PƏ�h@���Z&VU�m2��	�F����g��i6U� �rdv͢ ��l���9N��K�����C�mR�l����b�iA񁠛��{�;�M��#��A��n5J�)�6zҦ���JDZ�8���x�ǈU3�.&�ZL�"�^4-G��0�q��a�<�����}�VH���[�Yii���r{�b?q�N�y"�6u�@4��~���C�j�3�+�<Y���L,#��o^�"�{���f.K���gM= gQڦ�S�X�:/��Q����+��䕄�� `��b�u+Z��t���)c쥋�i{?�<u��qa2MR��_$5��A�x���!��W��3�������+6sg��k�v�i��1������ù�Պ�[^2�b?�>�݊�<Y��@}|y��(<Exv�'� ��=VC��'�J����3�vOD��So1).C�>#�)zS�|iB-�E,�nŞj��~��W���dªרJq��ﯬ���~<�\�pI?y�X(�6=hߙ����?*̜jP��e|,�)ט?; �ץD�'��.�W��T}�)^!PB>��i �w6�^`vtF�O�7�f����I��e��v���o��2g�=������}S�ľzw}����$%���k�˲m�3J ��!�z�hS�R�
-e]�$_�l
B5ا�ˎ$�N���#�4&�|�.��u`�� ӝY�ns��p�
mGý��WJV�S�x��/] )qB��ø2���V��lAp^UT���A�*`�ߜ�/�4y�I#K	�����o�Պ�t�q���^���,�G]�l~�h�K M蛌A��̝ٓ�FϽ�IAM��h\zLz�בQ�A0XV���ӎ���8m���1�P"�m�w�w����S�����6D�B���Jc=r�奒͵BBk��x� �d�z=	�mSI��G�%�o���
#²7��婜8E����6Ԉ~��00;rU�w�<n}�D�-L���w���>�� ���f�w4/}q��)v�ב5�C��G��A�9��3��nO�O�G��U��_�>&}<�
d�����W���@���8	�F��D��"@����u�"��8�Ma%��Ak�q�l�|^��t��-_���8��u�1'6��Ku��oq���?J*��rvP�q��)�s�b��JY�����%�D:����8zTX���O��[����� �nG�����	�B��%hb/�k�7w/�G|y�	�58����T�l��X<���v�1�h���C�� ��֒r~� _ʱ��z�(n��3�.9�ϙK�!�A�>u�imn�X�\_��%�e!^����r��T[�	#ǐ�P�賎��0}�]�pA5�[{b�3�Tmj�;�P	(�e����c�������k��\�F�w��[S_A�uo�Ͷ���Ϛn)�=�ei�1�e7��N]������Cr��~m�8cQ������q�}����=�K�O���WtU�X[uO
2\u�ȗjj$�v
���X���}g?b����v�N��]���K�*��M����"��g�����N�j<���/9gn�z~Q�^	�r^�pС`4a�?��L�o_�Ĺۿ?L�RrŒ��p����{�Z�]�οN6=M[Aw�ҁ�ƶ`ō/���$�ZO7Rs���0,,a1-�a(m��|��cYb�<l��#�B��-&�nf�ă�S�����eɧU<����ѰaX#F���j_������f���Y*%{Ʃ@�R3)ho⹄� D�u}�⥡R��uT��{���R�	�*C�w�GV��&F8���s�ec3��U\�	��cY��+���"�~5#����������`��+_^�c��?�w�O.��������[�Ä����4��fY!bB(̙���8n�	��r5A.�'N�5�P���'��0D�4�;T�i���S��"6�)�����Ѽ�E�](��H��F_��LpMO�?�B��%��G�j��
D�=��=�e�&�B1�OG�������U��-`�y#��:����+�V�C��@O�Ae^�m%E��]KR���A4$�I��oC��o`s�[{R�