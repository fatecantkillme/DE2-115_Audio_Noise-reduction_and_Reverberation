��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<�\5e�)��������O��2y"}����_��$A*��e�r��M1��WBy�T��N���|�å'�u�Miz��c�v�5�;3�@76+پFګ[[�e�)�ƽ��-� �%+��7��4s,��J�MOHbJ��]&j�٫gkG��$.3�FM3�*[>��A�5p��Ӈw,|���i�'f�����f?��7��L� %2Oa�
�1%��Ą�)אD��)����}����~�4�s�&Z[��^;j�i�9s�$�0��R ���l�Kи�vdYxw�l�����5 �C��ֱ�S�U}���U9�}�\�얤�g���Z��fu|�q�h��˳ͭ��D�l�����F��XT��4�5q�A�M#�:b�9�n�z�Ǵݠ��@/h��hw6�һ�0Xɥx�y�U��t��<�ނs���)2n��Ԥ���R�T�*c}��?�#��[HtW�}|�d�7w���8)��\q$;nu�d>|;���J[�&��U}Ƣ�i�SY�_�,�;�RU	@$ŤC3�n�I��0���6X!H>�Ouz:���dB(�V8m���_gNǨ(ȃXM͟��݄�/�a^��W��>�0��d �¸�*�q��e`�s������q$E���Tvb���މ咤|��ķ�p���a���"Hq�����/�a�=�x�?KauZ�_V#� �]���0�P���ja�o�LB��������%�c�n�r1�j*8zE-636���V��xX
v�B\�kL���?�y~*N���i$���ļW�`9�a�g(x�,.�Z�3'�Ø�1m���ӍJ�ul�O�d���MK��lL��W�H��s��sN-���rJ���
=�ӟ�R�ʄ'`JxW����t<U��N�~�Y���}�͌�a;aQ��ƗP�n�D�:�1��W���	��Ƣ{��	r� �*�@�d����������|y�H� �,�X�:C$�����C�����Xk��e{a	�@p�Y�Eש���0�N�Im��W<��BZJ��_I�v%����g�Զ�Wi;�b�6=p'U>�m�^˼vY�(V�7���T�@3�r>'6�/�b��9J���_(�~�����l�o���f=��r;�T���̥�0Lo�Tr���^�c�};n/�+ &�����!�]�$��7���-�q���N�fؽo1)�s���h�3L[�1�iL ��W�h|���66�B���U��/%�&)>N�4�����y��|7�֪';���ۓ�dU��*"LY��V��J���5��t5n���r]���TRp^��{���{[��2�7�>p�@[ς���;��e�d���}&U#�0ʁ�@n4��� �T�&kܵ�j)/l^d���u��yHB��*Y�/�M�[sH��
�)�&>s.����埍���v%���&'9"�X����MP�N6X˰;_�V��nJu��������@HY�h�����c�����Uz��og+�(S�B���.�^݊��$�N�=�C/����s�=�j��If�:V�`ƿ���+����|����^�_�U58���TՒO�����[)���_��n>�nw�����N�4<�1�x�,��n��i�����4����5'l���}_9n�79P�#��l��|h0bGh���ٝш�ܝ��4�C"��|��Cms��f��$sq'�������+�y@V����X Ů�G����.��i���Z�'�S�U�6��W��
�i9W�|�����^��: ��gGz�w�(h���H�D8�tI��.v{ă�f[A�ik`@��0���J��ZN��L=�E�e�=)���+�T-O�[�?�Bߕ4(_`�$\��!T�j�#8	���o��"Rq1���o�%����YGt57��ꖔG�(�~�^\�ͨ�d�%\��Y�nbş@�,������N}�L�:��� B��F:���t�U�0e(������k.���;�~�ɟ�=y��Ƽ�j͠ ����z9�MW��^�T-˃܁z8&ZCK�t�����D�����N�����⬅ҡwT&r���Z�++O�n���^
X�<�&���j�l����@j�	�cm�%�Bk�S��i�w��o��}؆C��m$w��������B
c�zÓ��o�h�	��rmfF��0l�;�]��h+����v���( �'�	�I����*j�R��c�GX�8x���e����4LW'e�;�`��N�&�Yd:�f/���m��	�l���6��

�2����%��XB���ݠ��E�u�G ��s�X��TɊ��0b5��w���8�0�ב��	�OSr��&���┹����t�{�#~���~���$Tz�B�3��\�ZhTg�1I�����p�C�~u��CN�_B��2M��R��vlmnBٞ�5Ǐdݩ���*�4<�Gś�p��=��Γ݊�K}��Jd�Ǧkk[N����7~C̓r��~���}��s~���:t##�DU�=뿔F�!�_����Zi�&n��)�0<՘n������h|��Z�}��u3�ο?v^�g�,c�V�����r����6N���0���[0�6Gd�0�s3�br��/�-��8��:��)�S��%��$�wѿ�E��3�YP�)I��~��J�Fsr	e�G�F�h>�
�	����!�$��H�N[�yY���+ڙSr�ҜX�So�|C^�wh� �����tK��FY_*2vN'��_L�����e�lp���JQ����(=r�đk�V��M(`*��q�3�G˞/G�pV2Y���pkm*%�c0�'Hi����܂)�����N����eA4�wVQ�� �C���7�1�H'�E�����>O�f�&��A9=�#yh�j�"����\��� AY�A�s�֮]U���/s�c2�@���bq�w	��|�i1��I�,�-n.
6����@�!L�j�H{$R�G�,�y�\� ۉw�2�=�Y�!!�)��/KF�X�t�=��aT��9e�4f9�� /�K"�=�Ct(�LH'���_H�_�����WP8=\���3�{_rVzlqz"eAca}l(�m�07��ڊ�����1��4�%+�����{r�b��~UQ| �Ȑ���8q�zꄣ�ޘk����!�e���7j��t!�_�|D��%��˨D�3�]�S�i���TS{bZ�W�%����t�]�H�I+��>��GV�jE���]x_�!���D���M\�����n�q����	��{�0M���bb��|� �p;�k\��w�Ad�"�?�Lj��>kB��Y���46�_��������O�r�m�����Y��ѝ�<6�"��� ���l'�'�㲒�t�"ZC-Z>_@��i��Ɂ�?>�&l �CPj�$JH���i8Ub�d�4�ٺ�ö~'9s��jـ�Pt|�'����u{�)�[(��V�3��1�_μ�}m���'q��+�E�B&_	ڒ��@ߎ�M.��CE��UeX���h�bRG���.�DNً��/Ak�����@�;}��~��D]����3�Z��,�.�R��w-0;` N��2К�(�rد�u��0U��S�|��'IM���@n��Pk��	/ ��&�;�SH��Yqt��ӡQ�Ê�c^�������J_:3�h�E6t����[�{�����?���eޅ�z�}���x#N�xY3*�u�iL�m6�x&�,�H�z���j� �f͌��cDC���_������60�A�ܩ-C��'<n��$�N=�c{���7���I�M�تoc����s�rf5s������2��R���Pu�Yq���s�[�A�pmMZ���đp��r� u���D��0�V�HMW�f��-��1Ik���j� nNc� Za�����<H�G�x�A��;2����M,S����o:>_a� �(�ɸ�~3r^��Z�q���YKi[4�]�w���K:��q�G�62nَb2��e�ݟT��P�CMp�E6k�r��^�[��=��{n&�ba��'�@:��U����c�L��=�٫'$�X��&艡hz�����Pm����]ʃ�MtNm�������(5j���Y�eV0�[����JN9�	l|oT�.l�`� �A�E&A�v�T�&�	�wtB����z�j�����"���
Сp)�ֺ���$�F��^Ј�/�D!&e ��N��}P�q��Rj���=�s���&.�����T �%�7����
7�b�x���GJ�in\��[��H��1�G|d;��/_�E�p:�r�"�_ܢ�GF۠f*1���q�ו?�;POK�3�5�Կ]�����B���do��K���UC%�A��O��bT�ˇ�K�h��cq}���u�<%���
"�|�%�n�c5]��oz���#����F�<^�?
O#��Y������CG�ڶG�Ri���O���bc1t�2���jW/�^�/�$�켛^u��Z�iG������	]iKv5w��W5��ec�M������J��{+�Ѝ)�]��m�H���[��:p�n�@E�t�7�����;l�E+~<���:�l4i�վϨ���~qk��|��p����ɬ___N�^��k�r��aid`�Z(c���F�惑q֯��p%C��R�kX�+�ܔ	��a2nO�Ϭ�L2~N�'Յtqۖ/��Ŕ�3�a��r�<�taO�S#��}_h�)�;�O5H���5Q���0���{I�"�p����$��]�#m��i�˫�X!]�w�3���%g�8cnL�j`-c5�L=������8����5��Ͷ�4%l�2�% �U���
��i�)jlON��x ���� lw��J\��x�sk^#��ݟ��k�=҆y�ҫ�%EpX��cM��B9��szMC5�Al�6����* ��rǭ��{���ϴ��Z����.���{�M�J*�#0�k)n8� �6Ȓ!�n>��N�� Nԩ+2�J��#x��>x:�{o�?�S���摝�6Xb�:�H��F�]�wr>�Mx�%]�<�x����!V{Ǝ?k��F�k�\��-�3Yϔ��������]6���Ɵ�� ç`��oI�'ػ����w��L�HF��?F�e���C���Ȍ����h՛ʽ�ˈ�~ u*4B���-F�<�O��������^DZ$�`�p��~x�Kk98q:�dH);�[���Ċ�.�]��{�F�W%&��[�=�K�˴� 3�*�i{~�\�)[9ż�'��r���W���}��?X�*�	�s�J=���Q�QwK�� �D�3����������%?{7�pM�- m{���Þ�)͠p�l5?���rk�U=�1�!L�3!��K��6������F��+�X�0�����?a�9t�(mw|m-�a G�-���"5c���R��VGc�r�\՞�\k0���i���N�!3����-'R�HY4!�$��}�g?h�d]�[���Fk��<���c�����l���K�L8t�΋����������]�1���pr�h:�.i{���u���B���!���T�v��q����1[\Hw�M�Q��2��ys��u@hf-ve_r�>DҌ([;Ԓ���6�܆ۊ51H�q1RY!�@�2�t�����}�L.��b�8�h�C�ǰ�e�����5J0U�~F:l	nt�Ƥn�����D�E���g��x�kLd33<��~-�_�-���2��,%�6�eaF��j�#�s�l4���:��Nﱚ��"����^kV7������F������dY����\��)(}��5U[�&Yغ�ĝ[�\2�	�qv�܋p�ޘ�1Ǟ�ڵI��D7���VV�rX�;�)�W@�x1����ü57I0y����K��b��%�O���H��靨�2��ܬ��C�@��N���&�	M<U�0��zÔ�������xC����づ�heʺ����q	�
�}�Ag�$%;��ু�Hv���r�M�˳8 I�z��ο�"��5���;AQ��/*����{.H��e��L5I�G$l�T��D�8�@a����)�t��H\C�4�"u��C<ݶ��`B���Ӽ��@d���P�����m`5Mz6.8Č�_��f���(�w�����.M�<{���1J��ľ�Qw����ߦڤ2Jv����T�#���\���J�X���Q�[Q�[�&Z��nh��]�_y���~���'�����]�:,s�;��j�����%���M!�޸cJ@�v��vĳ�uk�e�KT�f[K����C����vp ���+����Z@G4��z�tku"x�YU&��?9�%t��Ē������޷
1���-+� *�:�MRp���@�;v�ڎ�b䭛��!�=���wH���Գ��1;�,txƁ^lXȼ���l2-����`���N!�r@sf���t
Oz(�!������i�a��� CW>qp�<
���j:���V��-͍[�ԂkQ	��lZ~H�QKJ,G�n�..������6��?��@K[p���B5M�s�yh#z�+�O�ؾ��c������:��;D�緐=f$�E��n����.6>�V�=�G\wDĩ&m�y{_э�������	�����4c1��э�ah�f�4"k�֠e���<��.�s����*�UQC��v��G�qW�W0W�O@�s��tT�����B�n���W%�U�OŸ#,�f��,�j/�[�Z��3gIou�W�;j�%�q��#S����8ډ�B/�œ�둦��z�a���6��� n����K��Oȥ�Y0���,~���H��|�lK��������gl_>x���l蝕�l隉���q���*��'���;Ђ�lT�U4�X���	^p�B7t�I@��ϖpҎ��r��
C�հ���%�����وήw�i����s6L�b�s�
(W��:�c0Gwl�p����ֿ�4�b Q�1w�ߙ�}9��Lb'�� �^��
��K�=)Dy�R���X�Ա#��)i�7�ox��D`�oSI=H/�s~�\�����\l^K�LշN��4`/�[9�'?��A��*��,����I��/s��pR�YOP�OU#���<7�u���Dz���~LlZ��j�k/�Ep��4D����{���k�49��ek���2�U�݌�ٶ%���G�{�c���d��I;E�v��JqG�
��U�6:
����,�s�'Gȏ��A���7@���CUE`Sn���A�^�YO5P`ڟ�=1�;S�BJ����\�f�Ra ��6�~�ȬL���k�����������?�_�U��8�*a�wi�	Aiy4+��ar@E��r6���lXS��c�Y  ��p����A��f�y	� ń��x!��	�	��c�o�9e���c}1��p��Ƅ���ɘ����%�ؙ8���b�GB����\�ӯ��uϡ��נ���y�Rg\�d�M,n�Z�'w<Ң��5�e��4�#����DՂ���� ��\��a�E��Le�qKm�:�X������;j+�ƹwh�t�q��d"��_eaxK�����y����Q�/���!�GV�{.��Zwj~v�ߝ&xKlD���n�5���Ĺ��7W�iJmLj��C�B�ā]��F��ap��������F�˞���u�7 �dE�m&���(�z 26�<i��WT�Z�s7�TeW��.}���~��D��8�&�!���<lT�ȕ�ei;��n��Bo�_��j/�j��>��*������ф2�^Wd�N́�(�i�I�W�7�A��0O�&v��]��9{�,����,W�$�S��Tg�Z�S)�|;F-�F"�ġq��|��ا�B��e8�$WQ*���h���n�d��a �_�VT_�@����͢g������k��$L�k�x��q5����:���!�=�� pB���~�j�(�l���rGk�4����[k}���ƷEc�r�����<���u`�S6O��{�t�l���R����Ѵ�X�0����`�*��d�}j��Y?���PVd$^c�����<�����x���L�AF� m������"��w���%m�~F�P�66�-CrfH��@���)҅��]���K���j�F��j8��)ο�ߗ�,�Zaʗ=4:f�� (������!�;<�;��`!�p���|�}���a������u�yLd� �t��Sp�;�U�Gs��Kɇ�ȑح��+�v�U܏'�˄�*Ɠ�����Q�߲�
��UW�T%Q���P��~[�]��� �6�����y:��!/p�d�u�-��\�έ�L���N� 1�SX�2���5��C��$�;D�1�yH@d���=�� :�]�F{nZ��T|��&�,��\�� ��R������F��ٸ��楎P#	�p?nX9@ʡ.e��T'�m���R�hpxvOKAӒ�����e��������;�q�����#\�3h�|�8�RP�
�������~7@=�]$�m��˲?��6c���B��:߭U�l������qc&�0&�!	�NC1>@�Nշ�"SD��PS��DPe{1���F�N^%g����r��;O<atxY]h~rhh���f�y�����2$K����h�gސ���{�`�̖jk9o�=}M�ٽ��Kq��Y#O��	����L�5�����K�%��5�n�6�T7�W�$=7���b�wQ~��ڋ�ʕ`��xخ�����q>ec�s�ɳ7ƽqʺب�8�I,^�� y����[[�\�|��,aZ��!QL�_a$��B��Sf�5KT� �֗���
E��&����W�j�@��emy��aWɯ�Rw:T�(����	�<|�ʨ{-���t��5$|��W6��ʊ���n��5mk���owl�6�'}��%�Dc�1�kK�U���I�.#��v�^!�kq�03A�ȭ�V�Y��^���Ɉ-|�0ĉ���}`�D�� �6�j�ڷnde�h�>���������j_��t_��Rl��+Pt�wvI� ����'Z�r�';"�Z�p AKR�Q�.W]�Xk��}�)�����?H]�175��^|�'��:�.뱒���tJMV�]
$�_j���Y���LٱNd��r$nӢr���y��N��e8<��`�7ЪK�=i�� ��_&��'#Ӕlw�^M�	&��������JS�xEQ�O����b��O����c�I��7�miZnS-�G׍(�ˊTo(~Ǵ��.K��L'9Qn�^��Y�i�;��a��ɵ'q%n��z�/y�g��4��a�m5M�L=C�[�L ����:�[�
'�g��c�.�j����)�>�=���7/R���DvD��j¿��qfv��3/j{��8�t�e}�:.��/�t~lhE�s�SY�Ҝ�����0.U�~xN*�xo�t_�J��?9��A����j�H�\GJ}�~;�ů��H��J[Hв1��h����P0��"	�7Uh�*_{P'_�\t�_�V��
�P�:�m�����Ss0JYy�H396A��� �w�_��l[\��S>��V�ONI��M�mM�"b��ӽI� ���.�,�핣r�[�f����b�[:� R�R0H�=З6a��H٭d����Xy�rm�O�)�<���$ɼ�$��s�Ӛ��e��}�P�rs}�2�tb�5}FZ�N�o�p'���(͋��)mI&s�wѠ�&4w�FKE�7mD+|�
��^9�å[a�
B�ݸO�򎭜�;N��*i�Y�J$��b
a�?m)Ϸ��f��\g��%��<�4��^�\�����������y����)D�䟆�pN
&k	��CC :��c.\*���%I+�A!����3ԝ%�����D���Ղ&�|�8�Tv�QrO�-�3���I���3��,5c��_w��}֛�I*#"�q�Ԝ�W�R���y�����4TZD�v\Fhbv�k�8�N�f����O�緸�JxQ \p� 07�X�+! ��9�P����/�A�	=4�JE�̳�[��wr��ڝ��B�ķz*^!�����p��=X"�ЪmpR6���N6d�I���k�K_a,�������;�P��:�9L��Ҿ�1]��r�"�;�x\N�%�]�H��2'a�۔��I��Nr�8�=~4�N�l�}�6/]�ƥR��X����S���P��
�;rguUu�[(���8�}/���s��@��0 RsC;���z��{�������"�	��6��y��d�8�+7��˿�?;�*�J'�D�6�aX��M�N*�M�eQ�2)��!H�c#�H���a�Op^ b�i�����HR���1��ק���Z2�W��q� ��Lt�ϫQ&���3.J��f�l��nO����z�B�����w���!���q<�%��-���R)�!� �W��{�{pcUv⛎+I�>�! ��zJ�A�ߋ� ���ǶR%s��ݱ��)�+N�,��b�ƴ�8��%Q�_�q�L�_h
uϱ����+ȘKD{����q �xZ�.��K!3�e".l�*8H�(�Ho�:��}~g���D /QT��	4Џz�)�Rt�]qv�Ԗ*(ಬQo[P��c�x�	X�EL.Yw�����r*V�[��Kͼ�X�;��++��~��X��Vz%+C�_��l��-�P'�+ߗ�p���Ϣ����.���:W��]�w��!�q��%��7��toƸ������*��qi˃̼�mV��"N&��$�|xȟD��	��`Ms�)l�u���O)���*���q�EDle������h?�����˼h	���>�-�����֡�!��f�y�-���t��:�{�!�{��Ju�UI�y܆1l�3�Ι�:�ba[�s�_D;��\�b��S�ȣ+��Uw��{8��`��7.�7 x�Y�Ө�i��2 �^8=]���yo�vH�1�s�r �Y