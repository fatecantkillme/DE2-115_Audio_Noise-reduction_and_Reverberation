��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�8k�)9�k���J�f ۘEN�R��>�Ug:�&�1vB�dK�N߇0�dO�~g�2<YN��Yq�h�A2�2�K��Dȏ�p����F��Y����<Q�#�����ӝ�1Î�-\�����GJ�v�� !)əCdJֺ��"g@YQ����@�%x˕*%B��3�R|�X�븮��4�<+,�_䛶GP����9`���@��G����ay<�FP�G?�箪���"!>l=�p8�_,a���D	)#�!�BS<1�o��}��M��0��-5�߈	��>q��_���,�ϋN�|ϼY>��4]&/��Bn�#)^˖ݮ
���7kNH�o�Om�O=�jl3���]��2xu���*"%��7���ԪP�.�n@^����ϋ�U*��lf���Nʨю�P�
_�֒�2��1�u6����H�1�ǃ��|3I7�4�ŖR���zF�Y�vksX#$ڳ|4_���R�S����c{��_�j�Wy����<���B�!��da+>����ns���I]��a|ɹ�1�B'K���ӌ�C�F�����U�~3��E&��(W��!IȾ�OA��%��C�!���W�E�?uϷ2��8/�a��������;�T���9��H�p�Ajx �wU�;R���'bu;�?x�Q��)g
W`i%/�Pֲ��
�����V�\T���@$��p�]���vԋ��+�r�r�pY���V�ݒٖ[t� ��񱉃e�\���t�<�
= ���X�+ϝK��}�D��|E��uI#�s3K��Z0�O�y����@H�����w���l����_��Mݺ%(1�Z�W���϶�LgBe,�dو)>���o�9�0�\�����F݊'���f?�$�w�D��\^s¡���H=f�e���j�����8�UM��zK�����U4Pe.�9�Fb�2�.�����s�(+h��r�����ܼ����A�#w�wrX��[��+��n�I�z���Gm�D^���AJ�t��QK��7�*�p��p6���0��A2�x<�y��~a����/=�do�xc� [9�h:�Ӝ���p��p��"��Z�ƻZ�Y.ђq�E)�`��4��IX���ޣ6�"����`{�+(�hU@�Q��w,��-���Q�(�����()^��<c\C�I�x}u>A��U�,�i/�ޜ�Y����,>݌YT�slΜ�B�G~�%A34��[0a2#o�r:L������ay�K9�����,�����E�W	��<�v�n�C�I{���R3�Gv���B�y/Ŧ��H�L�$E��L�Z)ܴmM�ҳ�y�Wmo���$��O����i��[����{^�-��a"e�@����E6�S�T���: �StT�q?�ƾ$fN���Rx�)�?[��Ƹ���N;6�����J��_~|C�(B�2!��	�0�ꍌ�Ӟ7>+i�T�7��Z�64�O�?-�tV��Rns"�s���f�ݿ�=�u��c�􂍅���/��r�71�U�]����h�Z �_g�!�d��\�l0�Yl�t�V�1�_%o[�C*P�Pk�I DLQ�onGB�������;K3˕��M��� Ɇk�:+�_��f�V[����e$3��W�n�u��p����`)���
�"�uW.�)�x��L�%�l� �)�h�Q��#7���ӱ��HIE=b�
��t��J(��1r�UVO��w���--�F��.JL_�z�Ӄ����F3N]-}(�#������**�^c�LV��'�Ư�;�� �;�pՠ��/Y��`g�A>rz��}V,��C T��qvC�
͍�9:�}1K@8���[�N�����|�VQ�Y8��$`^EՁ���+"�����.p����?��n���"�	BT�D��͸��d�_#'�i�B:tj���r��>)�Bv�o�d:|�j�E��s�OG�Ԑz�|(
Z�d�~Ӧ��sԏ
*=fG/F��<���6�ym����[F:8�OvR��6�'����C��f�5eb\��4?B�9꺄�m��s���Sl��H�χ$A>&Md�1^�SY� ��kO�ټ�w���iaQ%��É� (f��d
��}l��C+Q��#��#��WO���J>WzO�vn/7�b���*���s�m�d��Y��c���	�N{���B;���&�-6�»� A;��KُR�*}/���V�����^��(�e5�P'�o�7Qe�cH�X�!	�
tj8�qpJkv�[��h-X΅!?���'���)u����o�td@G>r2[E_�`�Ie�%<������k\D�j샋�l��(M�Tr�W�7o���O���{��G8���(9@�\���L��'!��G����_�<T[�`��y�e�gHl����<�\����|]7���6+�P9�o���{���Sq0�@ο�I��l��f킻�'��̺�'�!td\e�X�/���Re��Wȏ���r�sJ��'�	��`�)�,���y�����&Ff���9��NR(���c�w;Ӯ���{ʁ<��T֡���U��t�%���?��i�r쬆6W�ytxJc�r[���MRNT�����p����9wIES~Ur�A�;c���	C��=��bP��3>�G�C�T�ww�"���/>��6#�뢪3OX���r!�����ܥ]@�7�.�)n�K9��X�bH�F���@C�C�L�n����~���]wDA�A	'���y���Onk�4��uw�^ac8j2q��r%��Q���"<�����Fƨw[)����ﮩԽ�MҐ*�{
W	��~x����k�;4�3.�3�a��@h"���C[xJJ`��[�*�2r�K�޹�\�%���0�J.?Q���͞4(̴z�(�{�����RMP99������b|�0)�]w��?*N��Ԕ���]���n�8ݏ�/�\L�����) ��H\V�6���o���H�P+v��+0�ϧc�;z���W���ٴ1�Ā&ƃ%a?���`���>2T�{ ��
�.��q"��,���n���<��އLZMMI�m���J¢1��!�C�,r~����b\�=5��ɀ풑i&��.���XՔ*������ ��)�_��pβW0o�>�L��+ֶ����I�;�	�9�=[#���t:<���ϕ}���;�M��~���I͡�n5b��E䙠�$���%�s���q�;E0$��9/MG��������XI��q�T����^B��87��2}����Q�t7 &'7�[�s*��ϲ5&l������]2�=¶�⣕�n��N/];����~�-�W�[?��9��O�ꗯN�Z]K�Ӳf��o#��+@���(��GZ$�:ZsF�'��)�N8��HڝF�����^��_��a�WN8�z�F��,���L���V5F��-{(.�T�(���ա�����W��!��TM��im������\i^2�F�O�ؠ;��H|�&��+r�C��"Y�����#!:pw�\Z6���0$4�2�p�x���$@�Gs	�w5��W;1�(w�k�i��opQ'5�~�j<������T����
;@���CѯJ]��	.��g�l)%�-�1>�:��Tf[�^*�;��x�;�w��H2�^�T8h"��&G=���R`���-&��)a�Zv��xK�Պ� V�:Ē��U#Qԭ��A1��L.ss���{9�Sd�
~��N�ט�#Ipl1/�t,�+g�\Qc}a>����Svց��H;ǈ�S��g��åR�>T.(V�a�]<�EY)�oV&#C(��
Bj#��]����\U��:i�uL���;�"r���Rl�2��8Unś�O��[�Yq�x	z�P�ab)���?F��Sm���v���R�Uc���hEh⛗�!$;�gڻ����>�A l�+�>H(�eH�F��Y��rQ��z��^R��?�7��.1�I�r�s��Z�P�H��f[ OSg����6Cw�`�O��U��I��J�Rf�Kҳ���\����x���ۂ�4���H�5���ajʩѩ�Е�:�����"�u����4U_�)k5q��uX�)F��\���N�!,���V@�ԁ���\�_dKK��c!���	�"��+pˡ���~��8��%2ց�E��~�a�S���:��667�rn��\u[�eJ.Ch�F��l&�ݤ��+��re�����늸�KbaփN�7s�=",Ҟ��vW;'�������Ȭ0�f�e���76x�bv��^�)�t��'��^r=YVZ)���Ǜ�UN�X�ן�D�"��vO�jF��ʿ0>j���*�Ke
�����o����z
�@���ܒ{�|���=�J;��a����`���@Pw^DN��ⓧ�>U>��U�<|��7u(Ì��'�E(C��*�{&��_�L6f��ϲ����8���R�Ph��Y�l��ɡ~�,��_���3��~���.3G�,�0�F"���!7S�ԇ9�����3�$��Q#��8���	��O�{l����_�0�_�ط%%��8�C�W���NR������� �ԋ�`-I�S��v��w�@q��X����W|�&	�M�f��pV�$}L�B�y��c�+A�v6
�����|ᨐ��7�J�<��=;KA�%\3X݇��0yϻ8�h��K3�������� ��mTACBy���1j�lF����`�j�(ѕ�0�Sq丛��	��}��!�:�_�u��w,�U�<�f>jw~�z_������E�Z�	��{DL��#k����:LVJ.e��@�������س:��`������2 2W�[��,<��?�Ol2�m����~PYY	L�s>@�}�`�n�	���RZ9��k[`h:�Dt�Re�Xlb@���Y�����T
��!"1���h<q;)A<�x�]e	lX�gݤ�O���b"]r|z�����c�'�Ò ڈ��T1�p�W���sa���tڜBp`A��T��OV��Ϸ,-||��DJ���2��������A��Y
!3�'VC[��L���Ğ!y��5~R�Z�p�����l�:�>.4 ��F�Į��iJ���+Zӄ�N�N��Zw���HS�G�a���Ҏ�Y��]>��,�8���OM�����`=���p��������������S~�Hc���)+S�%�_���-x�0��K5\^V��R�%�ZϜt/��W.���YMb~t���n�<yc/��Bu�)�{b��@��%ꗄ��/����!..^J��L^����$�?͈�"f���5kwS?�l�2�����h�/I�`���b��S���6�Y�G0���Ml���sG��l9�t"��_O�
��Q\Z�XVCe�鋲]�0��\�_{��0�J}�r��[u���V	ȕ;k8[f��.bW� Vw��*�d������fg6C�p�OX��(���M��®RH��A�y� ��`:E,Ay�՞[��V5
�0�C��î*��'x!#�D{�@�XZJ��0��8m���)������l��-�U�F3`Jv8�"m��wmЍ�9&L��L�Ӝge�c�9q_P����g��0�..�b�~�B�����z �*>l�q���oo���q�1�r�����{ L!�Y_�@z��ûÆ<���F�(H�֐�\�͡�˼;��%^�ͺ*5�6C����$5�t��'�l|aUR~XFSH.5G�y
��2�>�7ւw���u|�w���:�KЯ�ѱ#�����t���6Q�0�{��l�9���r:� 'νx��+��O�0�?�]�&|��y�������߸I>$?�C ⥃��wM���Y�p=hK�z���p$_�
��j�/�ăR�r\�����U���9�6�7�J	��ʁb���[A�oR�x/����%̆ӵ<�~3Lˎ�;�-�E����JLIDD�VhP�//��!z�UG�bdiT��A�wc##��J'z/�*�K�%������3�5��I�~�r���1[�0B�e�8@��n��`��|]Z��+�DYZ�2������BZ��ܿ����dh.�>F�n�ߞ�c���J V@*�E�v�P�� Dc���E�U/�Y$��y�rq��r��'6X!�"���Й>l�������p��;�7�m²�H�����6e�f�V~Z;!]��项/1��!�?�+>��ᘴD�J�MW�&�|�5��s��/��ٟ������H���a���r�Om�ud�7+��]���k��	)}�>�h�6�2n�Bdcr�9����R{�{4�F���3�u�0�F�zr�Q3��z��[:�t�ޭ��E�^|������:�����SF���a�_�ދZL�up��Ϋ�Im�Jm�p�����W�����%=F��E��0O}iiW��ȼ#�)}c]������廳�^�C��U�F��ǳ�l�%��s��WJ�� ��{�F-ۄ�EY��e��V���:�1��VO�yd����t���H�s��S�/ٯ���K_������,!2�,}m���-�-Fz�n�ؔ�?ǡ%���r�R���i��ߔZWD	OX�g
v�4Dn)���j%��#A
���6��b����o�����P<��׮�o��*�_̫�&�������Ζ��5i�-�c��(`8!^`d�'���,��	�#
[�>��L�6L<���~^�6X�'k�Oe�V"E?Q��P(�	�`b+i�!z�y�hC�Н���x��	��d�˶G��*B�\) �[�[�l�]�p4���W����F�;���LǓV�;�+��`2Q�=�p���9�t�igv��Ʋ�1nH4��<t�YRȼU�}J��!�,R�`�/(������aϟZݠ���}���mV?��d�ťI-Y�72ԣC�����
-��0���ϝ9/�E'ߍ=��j�VG�d���X6�Z�X�H�u{3��7t�z��p�F�s���1�˥L�Yv�,���e%�#�q�t�i�#��L!K���7}\PO�Ո�� _l3�����7��@��"S�Ssz	y���a9��`���y	��-��L���@P2��.�]�uH����3���f�}�z�S�7�II��iϢU��׻C�1L�nGӕu�t�a¾��r���s8�'�L_a���"�ĩ}"�����
��057�8*ÒA�L�m ���U��)�L���"?Z��RD��*��1N�~���P�g���ȝX&eM�ߡ�*rc`"�D]�R3\������0$o�p�I�ؽ� ���)��&�1��S����8�#�4P3��EN����
2������F�9h�C���O�R�Q-_w�ުWU��LE.����5Ķ<AQXV�\�:�Q����~�"�%��)$�ӹ��d(�W�{x�����崘����� E�h�.�3�E-ָ}�ouV�Z���U:�٪W�^g5>��9�q��;���u,=��tڈ�>Wx��Kc���Iu�ߨ�am+��k�
��I�Mb�^<������'aU��͞�h�<���9�e$C	%w_��f�Q`͢XS�T���]@�JD�j0�#����vhn��(��@E=��,����j����Q_��&���F_��{+�����Wf^i�a�t4�l��<���R����Y�%�`���=���2��������Ѷz��]O����p�?��ʩ3�k;X�����ԡ6E���_*ڠ�A��y9ۼX�<X���gjF�d���g�Qq0�U��7�Y��H~"�����Rٟ!�T��_p���5��)�Ķ�J�r�a�zKө����l�ã���/���Л��Ϗ��j���Z���?X����}G���H��D����SzR�LQa��
�;�*��r�&SQN��&�q^'�Ѐ����~�|炃�U��'~�a*'�<�\�ת��3qF6��mQ��mIO�-焭����"İ�,�W�-`�2�j�WH����L�F�e4�_VB9ģS�!�ӆ_�6no�DY�Ṿ����W�ק��ed8*�i5�GԽ�Pg.�`H��'�)v���c�GSZ���1{`�a&��;ٳ��ď���ӵ�_��,�����Ϧ���a�m�M՝<��&xm&��uc�.��}��(�v�6�45g�h����X�@���Ō5�،���ߨ6�#���ݡ� �����>�|5S?���d�!��Q�"���tӊdG��SUnAf�	��5�@k�����x�H���=�)T��՚#�[	��/���n�
;yo)O[9�G�;�R�A�;����}��з!�*;ƚr�U���r�#�J?�M�>ʟN<�Z����\���b9P������Q�ހ�S7��A1�C��c[8aJ~_В���C})�ٍ-��;���<<6Er�cƝӪ��yЭZ��8���Q��d3FD��$�Uʳ��A�o߅���*����L����e�_M豘�*Xȧ-kQF`@$��P>D$m��L�22b �$>m�?��RG�fD�Y񽙄�
�q�Ο�F��L#&\����An��O�'�Df������v��\,�p�8Z4��z�>����9%/��>�i�Ȧ]c0r��61,�zF�[�[~M�US�[�i鬳���&�2p��M6�f��,z���ݯH�z�$ٜ��ƴ�~z��H}��MsK�ES�v�� it���/e��h«�1�L��o��|��H���+0��Ֆ���6��$8��sA%����v�F1G�I)�!(�C��h��u0@C��ؾ�Ry�����f
������������E�2y��B���Au�E��xE�Sd�h�Hå1��I�	 FV��L��p��Q���ݤo�Q���F�ؘI%Ըc4o^{��?q\V�9SϺr������g��M�o�)���O���v����S'2@���0`�"�H���s���Y�J���2�� b��T��$��9��pAH���'��]������l8�{�y���>��í�m�������yA�d'�0���Ob�J�^>Ś X�w#wORnf��C�'�:����{1�jk(@��(^[m��U��J{������(���.n�gi�o��g1�FlLN�)yT�R�z&�W.���;y�>%�P?{�凙!��E��y����^q)@��!����d�/�;<G���U(��*&���Fs�-�B%�Ύz�+���19��ˎ�NX�P�Se�/��m�Ι�Ft�8�*D�1���l�&m5,���:ҳ�#�֣�d�+=m�p�Qޮ��h<X�w����`9��V���a���"�D�9�P K�[�c���e&�q�.d@cgrm��)��U�+��EԻ�8��^e�[�9����OE���Rjv	�SYֺ1�K���(	���8~X2�GF��fx�8o�}�<. fR�����?/a	��(��4�0��0� ��X~=����VQ�
j�q>�J�f�.Ζ�+�Ð5_�cX6�!���}��ա� ���d#�9y3B��󶹐)�;�p��y���6��C����{�P��RS�ͺ.��@V�O���x�o��=l��u/�hp
���$�E���%��N����#��9�҉�kpJJ�wG>ͶG?��a/ T��4�݈r��f�?�W"E<�� 0��k�aHI(Ul^����]�:
�l�U¦ɾ�GF<��ږ�@�u��D;��E6$��,���+�I�S�y�ڱ�_�^��[�DD�6t��1��OS��Z�׃�Md�^�<�.-]�(�}w(?���U�K^d�z4��:;��T�+���z{�������ā���mA$�'V(��� E�ϰ���F,�5-��v��x<����)��
�ܗ{��ۗ���V��}XU|�\=��5���7�W��A�笈�̜���>G@W@���h.�d+iLs��B?��m~'�#M;���Dec���7�@J+t�ڰ�C��E�Y�E�8���7c�0��rR��m1v݉h�"�Kv�<A�0��������uE�*�V(�l`u�}�d�u9�Ll���CoT賆���?���ٟ�D8�8.>M�|^LQ1x_��`Ͷ4M�׋��m����^{t�G=�W�e;7�+I��x<W�j�9�_��B��l���w'����p���D�!����Թȕ����'�-�9W,bidh�v��N�/:����4�2a��Ћ谀1ʹ�EYp���b��c��.Q<w���v��M�V����,"��%,+��{3�����ڦ*�n�\}r����ʹ��^�z�1���gb��*���О�Sm�+��!��Q�Y���_�U��V���!��U�@o�d�{�9�5��5�ܧ���t�n3ڒ��.�b������ �6@(����X�xq�|��j�z�4]2�X��6�½��kIƋ32��	�S�"�ȩ����)���EzHg�{0��"�Z�����,W��5}��P*�Y_?�/�<�"����^D_��@*_I�	�[3�
-hմ�Rٹ�~/��k�����^�ifǹ��x��$BC���4�L�!5����$���m#���3�~,�JE~��kxc�{"U��Vl����pc����,0M݀��3L'u7b�v��*7����1���^�Ɨ�r%Y~�l�8�q�D�eiޅ���3_�M|�{�Z1-f ��r����9�,��(wb�B�L�@@CĦe:7�N��E���M}��%|�8�w�I;�bDrF�a)4�$;WJ�IY�Y��"Ő��ꎖe9Fd�� ��I�Y�+�0A�Y\A����j�`.�M���\��L�����~��'�cIun�B�Lwe�U�>,��RA�z��~�6���QW�m)�r�v�M�ΛS1@]�g�I�Kr�J�����:�M��϶*��<�M�lP�v������Ai�A��Ӎ��IGh�
��H�eX����4�!��IJ'�5�����U����ܵ ���T�=0l��fT�<��蠆��bF�=�,/ˈ�c&��b2�#6�����鮵2��%:S�C8����.��|���A�X�@���˦�'1�K�Q�<�U#�[�7� ��LS���B�vy��1�����\D'4,�5�ޟ�u�X��Y{�ԫ����	Y�:|޽z�؃��(���N���=oq�	wmP��l^�+�����mszN?I��#�VD\t�`�w �&�g5��͙Y��O����d�_1�
��)m�@�"�� �-��Y0F���V�XOin�rv��]�^#���eG�@7D{�
E��v~�1�q���5�:�"@�*5H\�{C�)��l�M�H���^��bDo,]��u���7����e���3�݅:�-mԂ7��w�{��F���<�XK�R��;���^�jTd,��x�4�=ػ+þ�:���^߅]]U� ��y����b������6(ˊ�}�B�&`U�ᨶ[��r�����-�W�x������'K3�m�{]f^00�!���ӱs�y�O7�@0E��{��楤'_�M�����X�"9Y�$��{��;3E��0��!y﯁��]uGJ!���|B�]�\�]�n�
>f\ϓJ{I��s���<�;�7�.[�3��cx���zGp)ߑ"�'qB�~C�L���0��,_����~ٹ�|>���c���dz����_f��k�{�|Y:	&�Y�4�40ݦDgu���B�1��z{$�t$N;��-۞tf�Bՙj+2��I9���ήזU��V���j��wPxX�������d}�$w��X��~z9g���e$ÿ���ϣz�>� ��ʵ�x�ZgP���"�Sy��n���%�K߲�J �u��X(E<��R�oh�t$���>��U��'� ._K;�qۅ�Ё).`,Jǹ�T�l�xE�E���C-n���n��~��a�DfOlۥA0s��&����TzN#:�m$��Y?Vv�Y��a��?p-+��D~�C��u)�@��~��U� *� �����w������1��7�	�t�xA�w�&�R���l��E�3<Uk@�����U@�
�/�*#J��)u]�G�}�Ů@����@��@�L�(Qs�cb����&^,#�	R��k�ޥ� �A�0��eQ���6���If�hgc���[��G���\�a\`�XLj=["��[i9�jsB���$���.�U��&_�P����FJ
��Q�����T�N�0M�>���sT����d�+~�](��0�Q%o�/��O�쓂b�W��֚&.\r9X�Z��QՅԣ{j�L���)�%7�W�v(ÁD�v>��Q�x�Q�gg��_��^�3�ï;]�pܹ��G��}͗/�>�`���'�gR��6l�o��ʏN����.�۱(�a��|��އ�
R?ڶiF43~5���]=��f2�(����9v�
���{'}�1_�ٳ�3U���Xb�vն�ڭ�?�r��~M�T�
T@(�/�2��W%@�_(p�;��s�+t����I ����ks�Zq���;��<�&�dT�i�ދ�Ѵ��]��Z�V��6UGXp']@`i�Ntc�y��T�^e�3���<�������a[1@��N��5MWr�'G�K�D��������V��`����w@�T�K���{N� D��q�.�~N���%�N���C�~J��Y�겸H��I������:��5�=�Yʷ�Ot���+��`Y�fg���k5�!�o��`d��mN�H ژaٚ�;�Nޜ5STrHq�bэ��{�R�E�O�߂�6]�,e� nD��9^�Jz��o��:��#��� ���nR�~��L��6���j���r���0����!�c6_��q�j�u�e;,���3�|m�
h�$"��5M��8#��7��,y�d�*#U�(�`[�[�"�.��%��M�|��ϩ4���<�2qka{Gn�^~�85�G-��z�2��Ԁ>U�r��;����;�
?�p�N�5hbO�mEڟl{��T[���� p*�å�)瓤5��K��L���/S����1����{+`�L�3�+�ā��Q}Njؒ�uS��X#v�>`�W��e�C1�a��T�V�FG��լ�?��d,���26&XQ�>��~H	\g�9���*:k��(c�sQ�������#�����Y$��I���P{e<6�r�avw�B��l�2_�eA�t�\o�c>M2w�����iG5|�J?����*�\C'D��?�TN[C�{+�!�&�p{
�O������ϡ~a .K�l��~w�Z1Ȭ�[��С��I�"Ϊ������Y�B4P0A�y�9���Q��<�<��f7s�\/�����N|T�<���R�`K���%q�L�+Z~2F[�Ť�
�KCҴ��ݬ���v`;�z�Wd(~ɖ�a��>�:�� ��b5�Q�68�g�N�<\ݒ����,Z05�fz>�,G�j�^�ǝ��TH{L�23}�n��p:�Kb������%�x�h���I��Y;��$V]�P�l�����"��8����r��D�F��#�F��!x��X2��jQ6��(s읙��l̷��o�=db)�9�s����?t��Q���f�pY����\��n5w���4��i i 1̋�dC�a�]̯�̂1D�2NPl��k�J�%gh� �-�}������x��L�7�lO�̍A��\>A3|+�,�NnG�n�@��������?)��D9�>�|���dfHW�����& ��ڤE ��nJ�d#���2d��I��l@z��L>͌( +� ��~��+�z�&UD�,K�_.	g�c��!�;p�t��5>�T������"��Z� ��N9P2�<�a� �Z+�hz.v3�G���ͦ'��e<ßE3�v��r�ƈ������N���f#I��j��z��!< s�Nm����ԝ,s��.�>E�AI�c��@��ٜ)����a���;��>����@����JW�K��ב�p~����zW�
B!�!ԣ����?�	�A�d�����v����e��q�(z/'$�'6����f3��M��2�W�L��!R+D��^_k&Dԫy���-8eXʼ��j`���#�ߙ��t�Ђ��f/�X���*� U��Kp �vub��R��V���MK�EUV|i��fZ�����)p}��P�9y�q�8��M�|O�>.w�`!����,�a��x��] � �M/�I�J�^����Thz�^�}�6[�L����,j�t+z�k�˗v�PA6�$�c9p%YAW~�֩z7���.tn��{�r}��q�q��xK
:7���U�j%�*�)-��/�	Ye�>m��hd9�~�Zz�y����%�	�?Ak�d�:�/Xn�y�� D�wR�����y�k����.�R�
���� �K\W�ʷ��˧��:�9X����U���Mwܘ�3��s��wr��
�`��������:9 �|��u���5j`ƘԊ$�<1o��Ie�H�$B(�^Nm�,'��ϡ8Tתe��9ެƊ�P	��U�P뇎��u���dƫ��۰�͓@'s�*w�z�m���]�-ϴH�o�G�{��-U�_�[ }iB���8+�,Wi��?��l��T�=�pr=�5uYoEQ��D���e�&�'�����+�mH�1Z��X�uU��K�4�IR�&m����ɦ@g���C��������HDIa�`��[�W��i�dO+�G��N^N��Iqҥ0d�a�>��{^�>�|�X%�P��s#ܭ�!9NMs06� ���H�g�����1��F��IIɦ�
�u�x3�)³8M{����lup.�y������YBP�bn11���vOe��8Y����d�q�� ӸA�ۀT�B͔���2�ŋ>��`겺���WQ�=�
�v}��X�rv`�ԭ]н
�'Ӡ%B��\0�UD� ��M��9�@�5C�����C�'�2�S/�̰���$���k���G�+ηI�C�Ѭ97�p�'2J�5&���xKK����q|��V7��B��[�7R*��ꓵF��P���7ȣ�At7������@:�N������c�-T�fE�2.뻖}1��)�F�� �PM����/ ��O�!"�.��ۓ�Ov;m��%6��/�$��Y�{�7n��`��������WZ���G����N)�4�S{@�={ߣ%���4k6FrJhK�#�]Rc~�O F��e���)p��jTB���M��S#b*��_@a�#_�� �ή�9��ܾ�Wv-hW��Ҕ�'�������MNrp�0����4��.=��zC:���j��L�[k�S>�qA�:�ÿ�7{���ԳԤ!}]�����l�*|S�����D�cvB�XN��`AhJ��b�^*?duh��Ԙ`�ٶR����B�����l���P�̳�����y�KdJ����_���ֱme	��M_�ʪI~�c�)n�S�*��H�,�G�sȸ�G1 ��fD�F����� B�ͺ���B�7�+Իe�K8Tq+�[:�#�6�V'�ȅ��@j��;�0Z"��8���'���0�����g0�<i"�P�ݱ��T�����-�\kW���1~��08�#�d}�.���^M��a� ��2)(z*�Y�#�/+[:g�������ց�V�����p�lqƐ)`B��������\@�[�i��M�����1�?l����ي���9=���D)>�v�m��a��U���|.\���Fx�_~i5:;E����F�7!��d,f�Ԕ�怕�l�>�W�p �C��>�������UT3��O����2xY�L?�{��Z�L��iI��4�8(�[�����sZΨ�x�Z{I�?����m��&�qdF��[�����y�YD?D��=�?�D6P/g�+#~]�Hǘ���e6��ZG���22�1�_g�}����]|b�j�����C��5*�"a�"���xJ��v�[?P ��E���:��q�CFr��N��]k�F_�=R"
 �'�HNDmY5E�H$(�-v7WM�I��"2L�b���y�����0O���E���\"��*�z!eSO8�~w�����.B�0�W �5ypHvL�C&2Z�r"9�ʛ�O� �y����!��ˮ�$DB\�V`�a�3��L���yN@o�'s���-Y��wƈS��XfG�v�s�Ȧу�I����� o3Ԉ�"�+�-�����*�1�EfI���S��2�%h�[;����iɇYs����:��6���\���7�=��VC׽=�ªjQq�p���6QQIc{�4�s�MI�g�Ҙ���{<�;-�W���ލs�=�R��ۋîp��'�5	6��%��f�Wo��r3A�7JӋ�,�P.cq@%�E�J�t�C;4$F{������
�R�C>Â}�y5� =�>�~��Z��,s�ӿ��J]+��kIT�ŀW��d�Q��XU�T����D�D.{��EE�����M�}X>M�K��k9N�0�Ub�L���.�i�g'��l�l5��u{"�l�Pk���u.�;Sڂc>����u��x��~�����I�Rc������@��=
F-��N���+a�1� /kT�!C
��	�5f_=�{����������}6��A�2��
�'9%�Gx�����>�i��Ī���14�=�s�� �rUt�-l���n���ʢ�GO#/j�R�qR�.�e�O�g��w8�Bw{ �r�N՝�}D��
�B	lZ���Ѿj��pB'ؕն� zu#��X��Sm���`^�y��3�������ۘ|i�!����+�T��,[m��.Z�����m��$[	��`1.�������@[�}�W��^a􊫸ڴ ��Rሱ��R�v[�D�mM�i����鑬w����ó��'����Oy!u]�$�r��	M0b;ח�E��b��'�,�*F+W�P��_Is��ď�.���p���jM�R\��e�R��j!%���$�E\�̲��wq��po�Y1&�	l��d��o������k��q��$xV����X3��P�I+ϝ_1�k*����Zh ��Yl��Wz>�����]�����)��a���D��r�e��WǐVF�,Xӑ�E�d����M��z��C��7���4'�0j�}��Wߦ��lr|,uS��O�Y��Ӛ�� H�>&��x[��(�o�STک�_1;����2A��Q�&v~΢�}BmF.��()�ɓ:Z����Σ(��ݯ�a��C����]?^�-қN�d#���s{۽����/��=��Z!��#�Ytn�F��W��s:�=��5?�s�W�����)iE�P�I�$��g�Z���"��������K�6JWH/�+޻x�|��Ό�k�\@���O\�U�qN�Aa�{sj��8<\RFP�EBw���t�׌��!�#���&);�����e�2�l����@��`���GM�v�e#FQ6M|���gkz?��� 
�;�]; F��dU�E�o��ɤ Ε`h�⫈�=�^B�e��e�y�~��&�%b���$�t�{?ts
��;��(GzF��d�������P}��"
Fq�2CN��!b�Q��+K��p� �d4���������Y�����NA۴"��D�34y~dD���q.��xam.��Ȟ����1��o�9c�	E����v�����Hؗ�xe��V*��,�n�Jqm\�N��,�.����ю���w=�T�4p�oԎ,\g�R�M4Q�a-���u�n��9`��xv���	���J���)`|��M�A���i	2��Ӹ�q�Ǥ'r�W�G���&Pb��V&P����	��;���F�� ��6��縢cph����H�Z,�06�]߳%S�ȣj���U������[�C�r\�O/K�B�dvߜ�6Q ڤ^N��?�P?`>�թ�k�C��mǵ����Úʺ�?�A�۶ܐ0O�<T���ڞ�1�RS��c����O���L�/�2�o�����C��ݜƠ�{Țq�<y�����zJ�\�P�t�:-/A&e��". ���'��M,QZ
L�ʯ9��ؓy�7�2��������9"
m��_�#0<�_Z�È�U��7��x��z����_<p`���pmD	Q{ ��<�ߺ���7�����b��Lo���W�ك���w�)	���}���e���>dr����`�K�Ÿ}�Ќ�rD�١N�'�k�Z	�����UAq���Q�1��&U^��E\󿱲��M�S�!n����T�6�V�����lߨ4W�,�1W:��".I�X��7@���X��
����`�بD�����w�c;��Ϯ�.�zI-��i�����a�%��r��p�����qX���,$7�h詞��d�ma �btL}99����=�f��V��#e�)�V�9��]o�QR_��Uڪ
�Q �T9�yW�̥]�)��t'L0�;�����3g:�zA����r��m�$���zoK���C2j��#����^}�b��a�N/r���c�M�PB���R�5�[9�E�<��)�釉?�s�X��L!V�[��~�x!m�ykc}�<}���ˊ^�� ����R8]�dE"c!�$I��j'ە#u�ى��G�s��f���V�0��Yq܅V�]b�\��6��J�,����<i����ʾ�&�ρ2�?Z��4a?^��&q���T`�������~:8Nl���Nm�_�\�1K�lٯiO�)�?L��̲�>�Q�V(h��-�J
��"����oob�,�-C�Nh��hp!2M�2A����}��SN!*���H�6Q4$	Bz�?cQ��P?����9ctܛ�%E%{���c� @�3���u�<���E":�qiϵ`v)�Ό��В����FKٕ�};�%��s�ۊ�H3��V��X�}E�{��a'�Q�X%���oT����
X �Ⱥ�i�<�B���U��<mׁ�«���ܐ��j�J,�O�9$�����=8��� D[K�/�ܘ�P�#ǈ�A��^F��y��%U�<-|Vy׍r�͌�Ls!�|
��l�&�LU�R�}(����
�|Ui۝R�U��[O^i$���vY�ӊ*9[<��;tCѽ�H�HLF<`���8�5}�`�]��<�N��h�����@"QU�T�^ƚ̄>߽�$\y��/��.�t�滂�?�F�3]���Ɔ��ܵu�a�!̦a�����}�m䔠T`4�Qr�M��L�<�/2X�!'�	3&T�n:2�fr���5�,4d��n�<z&�C.b���d���]�e�&C"ᨶr�h)�]dBD�\�iH�H�I��Ķ)Kx��n�}ܬ��x��&�#��5<�r���P�@՞�Y	P'j5&�Y1��9�8�=������x�$xl8M��^]�+�K5tp� �^5��������~B$*�H��ZG��Z������hQ8W�+����p��Gϧ7�5��z�j��,*��j/�ء/��7���5���s�Z�^�xw`���#� g�lFwƹoՍ���a`@9�J�wo������`*����@�?9��|8l�Rf<�߂v=|&�_n�T��R�B��»°���*����Y�M��{\6#����8^ǩJ??ʛ��Ng�zť��wh���[�}?�f$	�0����N�/kS;S-��7e�6=�)٫����;J�eTC|	�&1(��l�I/��2���]yRl�]��-�{��1*=�ߓHI�l�{�#z�T��lz�^u��ڬkt����dFu��T���X��<�x��~,؃�vx#{��0�h��8�'��'�����,c�啽� �&�#)FlP6Y�HN[b�zb*��ß��7"��n� .�c/���� �Rә~���t��*Agე[:lrJ@�����j���XG������j���"�Hx����t���C�;�)�~�p<�ܜ�q����o&Đ���%�x�e���Б����C�eM�V��*�<��}v�J릝u���ZmÞ�5C�����Ի�!��?��$"@11H+���3~���mfϙ�zM_�A�	xr�q'��'VǮ�L���K;���܋.�j[]�ᐡ]!kN�Z�#�r%4���	!'k�uWȐ�����ծ�S��[c.4tcR}���@�5����d�1ՠ���(7Eo���.��g���ٚTby��(<`�U$كQ}︣!�x۶�i��X�kg2%a�?����J�&�ul����U#��!�i�b�"Hz�����Ǻm�a�2�D�q�F�60.l
�`���ˮϊS�ȅ[ٗ��.�=�+6]i��EFF�����:y��i�\���ɧq^#�5m�q��u������J���J}�`W�tX�T��m5+�����\_�L�f�l-Ӱ�T�J���'Aj�h�l�3A��t����j���u�\]|�B���_���� ����/��'5�J� �h��Z�Ն̞o�st�Z�(1n�k�6ܵۖf��Y��ڔ�%�P(�$(-��f8-f�C��+}te �;*�16�$�NԎg�r�a Qk��m���$��4{FTIv�Q���_&�z|܅7��$ls�%��iևèGޅ��a�6�q��<�-u��0��V�����ZZ�(�t�G��4���`%U��r6����3���$��$���Î1HO[�,'�a0z8$9�h�B<Y�rB����ҮK �~�0��6Ǉ���8��p�6
�{;�b�jj��N`������)�ҶhL�~>�[tLON��ˬ'7K㶩'PʀiC첂�0H�s�˙NԼ�!&9�b�./��bݶw�:I܁P�-K�iC�b�lب�+�T$Ae���րF����?�H�v�򑹐Qclv��ط�����=�Ȭ���x��޷s&��ob��&��h�a#�����yP3Ic����멡p=����*�.Lq�h%��ޡ��ـYXN��U(�
���.�ϺP*�~wC�_�s�J/�aP;Zv�#����~��*hX9��N@���;���%� �W�Μ��%�X!�j����'��1`�o��ťU
�:��+�~t�'j�P��?<�Ҏ�*��X^�_��QE�J<�.�U;.KZ�O�o�",K�\m@��ob\/8V�sm��p�t�ڊ�
0M�`��l1Z������5���ξ-���\>ܵl�A��]��I�j�ZNgFÜW�¤���V��jߤ��)���V�vy3��E���<a岅�z��b����c�� ����U\�_�S�����z����(`���EIဳ��<�o%;6����l5�Ş�e;����M��I$�v����7�^�	���~��L`�7��4���w�4�s�l�}�fZ�c;]'�7Z���g�P���2ʽ�Jn��}n��=�԰fp����O_���"��
�@mL7�mPr&�,��I���ʮ�` ��;�()�ؓ��O�]����[�W�*�p�P�o�����dh�'��<?�������}���_��>�:����W�Vt�qw'��'�F��fZ�1 j�a�P�S�5{,������N�$�Sz������$���݄����΀7����Dh}Q[�˼ZT���T-=����WAֻQ����,>����9�
r���?s�>pK�b��8�VM�2��'G.>Y�u���o4�?2��Ò��-V�>l�U߂���r��s[���yr�m�wM��RӋ(߁|܍XE>�Zw�B�V����"�7�S-�L���/�8Q�b�x�,�u:����VE;�������5Z�Y�6���'���e,�Z�<T���{�|0ir�Ea5���]��n�͞on���4N�Yd�'|Tw��;�ad]6���#[�%����HN.:��c�F]�&q"�BDǘr�O	4m"�ׂ	�t�K6��)��p5�A>�4�3�h/�ᖛL�j�J���L�n�q�./GS��w�� 1Ĵ��ir��
Wc��$3j�s(P]�\����ʓ�M�vr��G֞�gm?�5N�����E��O`��-�,�6)�.Wa��V^���nz����;�������J�ۤ��m��Y
sde�'D��%��0�{��K^e��+N���я,R��㮶��m�^���􂒸���}�<�Z���߼���nJ�����h����3�c�~���g����wB_t�����ڥ�畊�����|��$�6��Ȁ,��+fA����.�t��C] �|ߔ��U��}I���{K��-���~��;Ug�hІ���q^����-֌�W7����ȇ\//��r'��������ؠ����3s�%�֝���3L�V�
�Qm}fɊ����LK�[L檑��|O��)���A�)��� /��������CÅ(������A�����[�(�n>���������D�G0����,`���d��*�zX}�-?+�����Iםr�J��SO��g��;6 Xg�!ߕ9���o�7to[�lk
���=K.\)L��i�݁_�M���b���"��7q���L�=1�g�'Y�|���~��ߦEA}G�ܾ��=��K���=o}"#�h�:�=ȔzW��R�܀�i�A��T�˥tb��O�N
a��0�ly�E!�:l��O���d�D6���uX�N0��I�m1b�G#�4�w�+oi��]
<�bin���rbՇ��N�(�Ə��Lo�CZ�nԴ����1ևM��*S��=
�H0�h_7��l1���Ȧ��P���"�doh���ש.Ol��̑2����*�о��&����_ԉ���?YQ<U�`��s�A����H���	\�b� �k������3qc��xiX��"�_?��y6�������?C��"&�M�{�0���(��џ��u�G^���$g��;�^T����thu?�_/^�E� �?�?N�k��!����CI�I�uq���C�F�{Ȏ�bj�B��̝Piߌ4!�KRϒ!�S���ܡ}wFU�������Λ�e锆�Jw��ONӲNA�����ז��GyN	��7c�ި�&��ԗ�(�N���1�Z��0"�4u�`��.k2�$�FçX'���7(ǣm��H��a���9ճ��޴p�i<;O@�u�:�čfpU�	P^��9���z�|�J^UgEG?�����i��ͥC�}�\E"SC`X����/[{#�*a�K�� y�>��an>��f7���J-)�'T���K$c��d��O�E��$�1m�0��Z�s/�;G� �3;���%��A���6p���)���a�W�.�]�E��9I8�#�Qޙ)����{�X&l�4��j�
����ib��/u�1
z���V�ì���Mqi�D�t�V�^��ē��'���՝��q�%ǳ��FW�7:�a�В�t<N�y�6Udy���v� ����X�F�SjX�Rk��w���]���p�8�����\��橍�J!�0�XQ⡁�-��hA"����{g���%	yjX�7��DoG�˽����׬�׌�Z�J�`2گS�f]��W4LY��+ʄJf[�둭aH������}%�:�(L0�q\��j��d]�?RsB�E�U.IT��\�����H���墤18D(���Grn�=�j� >��5`.�EH:��
���0�%��B�Q��ޛ+��SgfX1ɾ�� 3[-<������|���>��(Ҳ�	-�5��e�9�`SM'#�C�b�d��%vk� ��8�hps�e�o�+y�2��Y�w�� ݄�Ѧ4����(�6��ؗ����|�t�Y�s�v�a m� ���B�W�-0�Qn;j�g.�� WmUo���+���ZM�����i�G}!�+��n�+nk냑o�2�J����X��s��n
_IY�{�M��Y���Q �V�1��z�7�f�^�������%��<O"����0�B�:�g2�+��X��`P��%�������u���H���h��#ڦ�:&�=Rۃ�M�M�A����� � �A��Y[�u�O��w� �.]Y��얟�����<��ށ�s?��.��?��phP2c����io���q�V�CH�,��o��0 ��QO-�ϝ�U�հ����
��N��1���ol�ra*�ZaK��;�I�&8(]#KwKd��=}K)UH"O�\�'����uT�&f����F�])X��	�D�F��u=;j���n��;��L�v���Ę%BE�^Vo�G��;������i�a���1~ţ﹑�^ӊ��(R��?�,U�v�8\������E�~���>��2�jyฉc�����#��0�W����ɔ����?�/*7mY��6�Ց���1�[�x����a���C�^��n���Ќ`kij���z�K`N?�HD6�tEB'����Hn�� 6�Ҵ��Z.>q�7��	�%=��1�a�Iw(�ר�Y�pF-���*G]Q~"FW������Y�nn�DYh�vqʍ�O�]A�@&iȲ}Q��c<� �*��]�n�Lib��Fۉ�+�m>+ޏ�\�"Q���͟�LV(/�˫B� 	8�a�i� �ڊfOJ.�"��(6l�|g~Y�q�T����8Lx`uA��B֓�v(�	$y���Us����%FЗ"eˊ>{%���J���P�H\��R$�Sb�)lHf0:z�S�,&�N��a�cT�8Z4�.�h�hN�?�N/��UĨ�� �S�XqS�buP(n�`�&%O���<!1u�����`��\�X�<�Z�çHg�����w�vw��m�+t�3Ŕ��"7���l�������glueN��$T9l]��T1�:��.��+5T�(x�2����ni���֮:�J��x¤�#�l�0�F�V-��*�9,�oa溗�r��C��
S�����[�W�
Hj�8�.=��u���^����ҿV�E��m��_hn�!v,�HC<��G#,�2�rJB�0�eL�px��L��X7���g=tp�c+�I���o���J �ˢ�w�/���d��7gPOb��"W/� v+r�m����3��e�Dx�h-��	�)���h�e
�Nb𧄭�I�@)hϵ&hC�}��P��4s��ܞ8311��P��A�2B��(m�]d֠�fS�X�Qb�O{��C���&�qTB���+ߪ�k����b�W������@b�����i� "�5-!%-h�hg"8�u����ȢS�"�	�Y������a�R�K���MB3���.��ѵ}���?R���u<J!Z���z�Z���j�`L��F2�6	�Ik���=[���Dc��!wٱ�A0�_M��ӱbλ��n[k�_�(����������=��<0c�sr�J��ԗ��Y�_h��Z�� -o�����i^IP�(4{�|��9Ek�ܚ�w�%"+���~�)_��w������#�|p��D�i�&�c����+c��Nq�\�ϞZU��\^!���k��^����D[8�a�t8�z���"E
k��D3��� �	�f{يS�Ir���'�����l2�b�4.�{�@-g^��y����c���g��A�듷��D�(ٳ-iQ�l���+l��KA)�wJ�W�[S3��ఛ����'v�Fd=T[wC��qo ��MZ�ri��󍨤׳�>��4�8lp�A��b�6\b)�7��y��S�\q��5$�����+zFC{j�C�����D��4����|Hyf�C��6U�E�p���=��2���H���>�R��i�����m���{=HWŁ�֨��Ë��	B����!U^;m�6�t �����n�()�g��0:��;�<�=���g�X�SB�S0p�U����Rи�n�V�0q&n���ԇ�LӪ�idguOC�!��}��%��/B@�7}�ƔݐLu(��M�����;���U#��Ț�
Q<�=X9.��E��Ij� ��՟lԺ�)!�({ҽ�� ���
ZP��;X~��"�Y�ȖY�������_g@�L�H�8�r�L{Ge�yUԀ�$�t�et�O���P+~���H`V� ��Dc�'m��Q��t���~�L��M�m@���Oŵ�YJ�J��[�`l>$�x*<:�+V\EĔ�:i�F�f9'� ���*p�@��C|F���&��f+Fo��J*��������m�5�j��P���Yn.��V!�s4 ����iZ	�9ĝ��t�c��w�꜀n��V�$�������RYMx���,���^��!�D�1Bg��"%�mʁ/�a��A[Y.�{�xJp-��\� �6P@��N�|\���ޱ�]�|��\�o|jOd��o$����P!��,�2w�%�B�/}(g!�@�Ry��&���8���G3�G���#�P,�녖�}��������.�Lr���'���|�m�q��:"޸���s�s�IϺxs.l��>�C@a?	����������
���=!��-�3r+N<$^��U�7l�$a�9��P���*۹fnYbKT%��H.�t9f9yI鱊�\nP�F�٢I�t�>��'�/Y�(t���Y�T�����X�J��d�!�y�Z�C�x�8�v���5B;��?�=jK����'�� ��ڔ��<R۲C��
`�J�~�"�^]|{`�)�.=��y�s[҉01�&���}��������[�q����&�}�en��(�z�1�����ڼ,z����s�9�h�A3G�m'� ������%-r��8K�凥��k�aq��@��)�V!�Aq3s�%Ħ��J��Qc�'�R �h��5>J�Y(S��9~����~��V^�:��kv,�����_����������I �Y�X!���ݐ�T���p#��f�Iu[�DxB�N�</wd/��ԏ}��F���؎�p��.<f������8oV4��T���,p��|�`�D[ǁb^l%h���zA�2��n���X�]�����O�ڞZ�;��2ȭ��X��f�ZS����f��eLw�ZET�$��df�ά��j���j-]�?m��2� #��ۤ��/�/1ւl�R��x��˦��3N&���-C�g�%H��q��Z�נ�����ܭ���A�Q1�k�������i����3����8
�m�B��ShG�ժt)����;t����a#,��E9�Z�֫�l�e �2����	 ���"�j��}�߿����x�@��r;w��#4Ǒ̼��RŤ���g�R�"�~�iY�p����u1�{��:)�G9���������=�^���*����"�j����K	�P(�x���C� �x��e�}@F�z�&~�y�lm��ؘ����Cŵ�˰�޹���G�w���;�}�^%���9��:&�ǈ\��tb/����[FdE����DLN��go��2T!!U((@}]��ĦI��'��e��T���&�|�Ҏ��pU�T�&<u�s�Ҫ#ǖ�z�A�I(��n��6)��J_CjlK��J������mv`�J,������\��8$h���vO���D�=�\�6��lh�L#��C.N��qi٤�n扬ҟ�$�"�{�K%�4N�������Mk�	h]X{%x�~��>4�Y�^��V�������wU&�����s�s'f^e��뤃��o ���:"g$�B.��܄�	t����{m[���⊰�RG�-��Q��\�w�,]�e������Q)��Ɍ�"]oa�O(����k�p���	�e\z�OV4}���\Я%�W��+;��õH
��$�S;�x�#������^Wg�T�ӡ����N��m��]��Ȭ�IW���I�Oif����"����`ճ�d���#�m��1D�It���
�pZ�X-�2+6�ʗ��M�,'��{�Wť���M
��e����L0NAR�)�� �����VDٹj��X���M�E�N�="iF��uf�@��\�('gp�":|8ܼ�:�}�6���!�z�)�m��O���<�g�-�{��3�EL��A��AS�<wY��a��Be�C��]����焋SgE��zp�Z�Р���e��2��z똆��s	�e�n��1�"Ng�?s����:�ꉇRd׋��%�B�l�-�\�M*V�5G������%����r��1��UvK�Wp�N��x��9�Ǿ:�J��,���-F:ذ�x��>�b��ok쯊�Bi�C���3��ꡱ����&��(*4��A5���<�⬽Q=��M~$��)��忰�(�R��Tͫ4G� ��3v
��h'ʂ*H�Ҟ4\�3�EQc��JD�VС%�5yw�e�@��֗��g�OL�=�»�F�%a?9aanaW��m�.x�'�_~ |�R;��m�q;��Z�{U2��'��Ѫ�j1�Z�b�D���4�{C0FR�DC�+�*����G�kZRg��'^����~�[@���j��X� s�6<Q�֠��",�2��L�gGy�������V�y>T@��Ϊ�b�jE�R(d0
��!8�UV���s`�I�!����MHw6#���&�aƌ��:Zoij�sc��f��;b�%)N����-!+��QG���77%X[=\׶7���cbb�����¸;�����6�8r.�Xp�q @w4��!)�� !�ݖ!��S�~�.��p���_yװ�=��נ�8�5�����lt���9k���py���W�S:����%x�R1|�@�ΰ1ӺW�>P\�/ "Rc��r��d���c�����RgK�{.��kM��$~o�����Wrt��N����ؒk�� H����W\?�����
��������l�ϕY(��+>�� ����U9�)27�Wоg3�1����Ẹ����pkKQ�2���c�m�[�<?�	f��T�a���'��@`��$C���!Ï�4�����{�郙	�pzOټ��)����rgԩ��w��g�H�PH8����˝R]X��9$���(l(��zě�8�KWzô0(�W^b�e�����>C����LC��9N��@����r��U��>!�Ǐ����@�MA�)5GJ���6:i���+��ɬ��`o� a�Cl��//P	ڥ8���t�Hb�[@�U�L���4(�*����-bN����y%�YW���S�+ϋ���{|h��Lpqճ���T�`����?F��3�k[��ю�&j:,~��; ���oyQQ -�S�^�>H<>�G�4��W�e��d�F�./ Rx�r���v3M�<���D	�(8c��W�Ҥ��ʱP����s�S�Zz����eS)�H4��n��ݴ?���ɱ���ة���Lu�_|5��&=��ϛXB�$�X��^�������vA����u��Lۨ#׈8��3��2���ϑ����o��#|%��og����L<��]��P��v�:�K=R
��92P��q7�(�Z���>���2GSj!��Ϭ8����ܢ. 绩er���rj��S~0����xڳ�͉�n.�E�c�Q��Ml���� &����װ������`�6pl0���,��P}e>mq�#i3�ce獕���ޓ��Y��ӳ�.Gr+[���[�n����G�<����<q/��_:&���܎��#�4�z�h�sL��ћ_�l��'S�%�����k4��M���$�����Nsc5�ES����O��h��=��]�f��{ͪ�R���H�߳p�W��^Ĝ�H��Gr*^�&'�׹.j����|i>p+Q_��CR�t�����K�T?�Sk[�ƥ���u�8��Ms6��I"��֢L�U[vS	5�'� =��m]$��i�W�U�z9�M�j+�[𝇐�*E��ZB�3Q�F��9�/Yj�ϑ>՟��DQ�?��U@��3�@�2�a����o�l��(���l����2�"�|�9�M��U����M6�1ɫ����8�8�Ŷ����ߣaN��8
Ab�[J9��붢�Q0'zDL��,m���Sw�=�¡!�3O?u[QY޽�Irh{�^qPUK�S֮�D�]�nX�Qt��B��CLF��O`�B��c��n�f�U\���k�[��ѳ����p=�i��~N$����M�(Ս	�tso��D'����o����_&���*A�۽��6�g.��v�AxC�龛��K�ɤAj�ԍ0�	�j��Đ��	z�A�68�k{Z�Ɇ�� ����'`��h��3U��'���*nx���y�Íe�����KI=��X��U�����m�ZH:{��}~�o!�	��|b���ꢖ+f�L])z������y������i]�m��	�c�LqJ�X]g����I�*0���e�lh3�@�jM�ā��Zm�R6)Y����f�?�	؄�u}��w���pKQEM�hJ���<�I�#|�����m]�^i+t9��D���`����-+�O�.Qn�E��ha/����>��;�hl�D��n���3���5�t��N)�.�_�8��!2��!/\J�����y�>����i�zG{3)���I������Bŧ���-��t�"�8&cc��O��b,"0Ӑ��X(�mw�+f������O0����s� ��Ί�QCdiyȾ���2gR)�
}�+���{u��5�5o���b��ae�ꓧ#��D8���ަMI��5�R������MeZ6�z�]K����R;,-yTja�����y/+Zj�/��
.e���k����%fb?��H#\~��#\���2~����Ӡ�)y=� ����ӺE��&���E���ah�9	��	*e˩��vn��=$J �c�E����E�j-�K錾��T�y��0�e��yh���~�����w))�?�z�����1��W!pxl�V�[�r�8LsP"�et����r�'�9w�(���}he�tpT�L�/������-�H��{��9dַ�8i���<��T0z�_�D�ObJ��w����R���1�� �z����H҉w��/�0�Q�ĕ?�氍H5�Pw���h\��_v�0dn��\~W�g]�"Ԓ\h��
�0���y�(	�3����h�yt������و1��Z`*��O�'".��梛w�����/˟"���2�Znm˓�o�7��ί׏L���a|����Q"۶���m�#�8p~X~Ucr����R�@}���Ͽ4hY��͑�d�+�����/�	�^�_�r5��?�1͐kDI$QT.k�>ݿ쯦-�?6��'����d��.+�� 35���܉��zl{��¥b�fI8t(ʛ)�(�寺v�Rդu\���O�o�~����:�Q��u�9�b��O=IyR�LR/F�q��V��L&�{�.O�.e�:?�q�(ERT6����x�q�2�gߤp9+;��w��D��to�V�~͢S�񹮶s_T�o!�N��Ѕ0B�"��3#k�"��E����3���$��H�(Hp�\(���`ܔ��#��P.�&����b:�>��<(��ֲ�Z�w1n��M~c�����NHWJL�=A=��&��L���#`7�7��R8�_<_|Tˣ<��3�b�� ��d��	�^�aM�3H>���
j��:� ���L�U�$���*��)�d�&x�dZ��7EO�c�(K��֩���Ǎ�ѿtbJ��%p0Ҍ���,���6w[�a����}5�����g�A����3'+RV�̐	bo@,޸t4��i�߭��m�3@����;��ކ¥�a���
�f�æ���`��I��b}j�5���VG��0�_��16���|�l����Q� ���wB,���7b��=J��}�E��!�.��(�$EVcJ�������x,�BbȆ ����ʮ��3]��C�x��k~[ـxV(�\��4����Qd��h�Q�N-�/L^y�l{u�� ����z�ԑb��v�E�0938{x�P�'�r	�������X�
u
4f��������ټM=;��d���_˗s6��OOL:��+��3f뭷�l�ޤ�C4f᳢�"�4�C�/�T�#H�'(���S�:|�?=.J3�e�sƯ1�K��^�aW�hq��}��^zO|2%���!]�cc�J��qʯ��څ��%��}�����
T�[}R"	L�mF�a�$����}���D�py�А9���B�F�x�m���i�I��� ���!�8H[�:-!�v��δu��6΍I ?4��T���ǅg�\q�kLJ'��'=����9��!=�dR�Iǵǋ�/�<U��C��L�_ ���H�	<v��f���:��y��k������wk��2ݹ��::���Aޖ�`7����$������7/�����~���*�Y8�!�G�B�*����IV4O�_1����4�:���T��8˒�Y+SgW&�07�-}�P��1���u��,ɓ�o�ب�������F��~�)xze�,�7 eͩEk�y���C�r�aѓm
Kz��#��"�֠��I��V�o�=��B�gs��;�������42c��1�e/�Q���3��~E�YF��n�6±.�w`
Q3�/�a2p�y�I����9��9�qr*%|��W�e��,9����x� Ŋ%�]r/(Qh�r�Y��pA���o��7~:�"��f��qB�޾H�Z�O����h�o�M= �MZ�I��Ҵ�6S<��*��R'���u��<�Z��5���+1�ztx	�ŻU�Mm�����������US΋V���0P���G9ȩ�$���1�A]�x�
�%�#Z�&�lp�4�gpNAx����-�&mяh���f]��%'m�ֆ�:����c�}��t���,`���x�<�<���; tX����*�/Oq�h��&C�;�q J�K�4�k�@@ ��h�����!qVB�N���u5�!t�2�[k��%
��p!�M�M�F��j5�����j��F��:|Z�E2x����#}#�99Y?}�_�輅hi�h_h��k�8bX�5�t��s�q�G8-.o!7�Z��1��W[B��W��`���E��K7=�`��R8
����ʿŎv�f�MH��=跱)��\-V�s�<+9-$D��@Mnp�|�8�.܃{��!�L�!�_��$����)ݹ�S���FڨEr�t�[����N��OZ[d`�T�'߶�暉߯��wf 'R��H	�w��<�� ��\4�l0jb��#�(�e��	�5>	4r=�3�a	s�e�9�+ھ;v�ї�&j�f���K�;�����K!�q�4�xn���Pֻz��ġ���n�{Q�\�SA�e��σ��+������^[�"a���mRN�'|ʵ�
_~�*c�b�
�邟���DVtOd�;��œWs�$��+_��ǏZ�/���ᕼo]q1�@�F�:�P��#�T�W �@���I����50�h�k�����^��b0��;3�9'�.��P���N�����/o�>e@/'��|���t�o��B/C]�q�vj�`�P�$$���	|]nC�4�<����Y�����j}zp�KTD�7�/+�)ƕUR^��2\� m�~|�D�;��3׷�}���yp���@RtrK@��s���:��R�[j��iMBM�bb4*y��TDU2�(E]�ˍ�%����#7�X���5&�5���1���@��#]�2myyh�(�������*>�n�Bj_\�B�����ު�Y�2'���*���O�,Y���ȩ��V�bkSn�Ǆ����ܨ�iD}#��Zy������ζ(���P=KV��B����S��)���r ��.�0-y��<�o�O-��j7���L�b4����G`�U������}~%�o��@Ȩ��������u[E�v���ؚFI����$�T4W�d`�����E����`�v�"������`����m���4/E�R@C61)ǄN���+Gh_d��!��Y�YǴ��<�Ǣ�N&!>t?��+-^$����ܗ�� s9*�.�n-(�q9!rn���S$_XXme�����*{��/{���4�fth��UX�NG�/�ڦ����A�o���$ʋ:!߶���<�ĕp�G�Z��@^��"��N�<�Y����w���LM�y�:ٵ�}���	�h�3;�q�������ZM�N4����'��1�x�� f�kX��FM���nϋ��{/�R��e�>�����Jۇ���!�1����I!�?yv'�RÞ��Rk]7��s�����  �5�U!���4؛挅��ʽ�11޾�@�_�����i�vA��w▔�|�Z ��n�m2�śM����^3Pl��׮U��p�3k9C�L��� ,�g|ZS%%���o����Q�
\D�o��~��c���,���v�-Zo��>�eȢ����+�3a��S�0�خ�'9k�f.!*������:D?��u�j�f���q�} �3wӫ�,�T%E,O�ܶ�M֖r(&�z�ZH1ٹ-B�FB"��A񒍜p���j`fɺW	���x���R�Qӫ퀨A/k��l�#T�@���6�J���*�:s���4�n��8��n���_ ,yTgdF��@;e��BG�K��F��H�	�Ƃ���V	��y�[�����z5��h�����a}m0k���c1bf�k@WG���3��r��21j���9�,�u�k�N��iE�����a����2_����T8���ِf����O(W�V�)_.��@��T��$*.;�q�
z3�~q}z��b�d&�gܠ�Q��K}��}���xq �y��4$��;�?�VM�J����-7!��JVh�e�k�TmL,�HhR�_�V�;��LW�Ʌ��6�s����o��Σ�9�NG�y)�zx���Ԋ@�*�5�R٢����.���U�I]���c ���{���QB�~���!�k�w��ZY�o3�΋��C��1��}�l$(�ާ����!k2�#�f�9�(�iW�/ɏ+�;��-�y�ْLMWj�)�uWʯ� G ���X�2�[�l���%Aa����@!��!����D;(~���#)fG��6+�B�T��!���o҈D��z�p*.P�G)2tpY����<̞6�j?KӊZ+	���;�3p$7D֕��#{�t^ނM`8,� ��o}�[�Ϟ0��k��qq�3u�"�_�X�^���.J��9x��1p*b&J*����J�-:>op��=��p�������	������	
Z�ܭ�ܶ�#��A��-����R�L"�m4���O�5Z���=3��=�)t��R_�.C��+��|N�:+>�'ΐql�U�]�3��0��"mW��=��&7����@���+��f���1���7����'p�HlQ%���!'#��۷9�L���k`�eDyZ�8
�ɥ����ݒ�Ok��t��*��<�懡���ם_���3n7s�0 U����U���r���P��
�\b+�#��ޝ�jds��.�Bj�0*~2=���b�~æ~δn}�դ��G}��	�U����-Ƚ�b?b�M�j64�Ȉ�� �y��^VFG���
��׆`x��D^RjM���TJi�	N�=@N�͐p��)W������P�\�CAy�S婖w��[�#���,�5��g�T�B*5��?�/|~��Nz����q�c�J��|H�Z*��,�2�*?j�P�5���u��-������k�P�NM!Q��яQɛ��`�\��a�C;�J���0����8{��̐��8'#Jo}�+S�wu��X%
e$��m��S�EtS����ݗI���������*���Fb���iH:L�2斸�������m$��$״�X�y��SI�|
�ѵ��9w����A^t{g�k�O�Q��-�}7N�"�@�2;W��6�Ɯ�z���iI�Z<Ʀ�t=Ŷ)�P,i�����j�3�c�N�!֫>N��2*��z|��j��X�ֲ���0YN�A�AȒ��� !�&_�,��/0�٧��ɗe��1�20Ò9,�%4B}���pug>2ؤ��7����}Q�,�F@�F�
W���I��h˽�@���"���t�3������X�SӂI  ��4A,p�h�$�����eHs Q��WҦʛ}	ġ���ȵ�W8����OM�Rv�`0�v����D���t,��B2���⩡פ:�Y�} Xۚ�S��2U�T7�O�z��p %�[���A��ˬ��pX�u�*���&����}H��B�IC�^��)���GR�V�g�����^��[��6Ԣ��-��" [+ �py���8&�TR��Z>�(�!R�1C-i�Bۣw�p�SU�eUaO1���� (J����X��ƧG��X��\�b��b-G��'�_֔%��d0#�I��~�wo�F�=�'�9��ʠ2�)�*;�GW�%�U9�c��g<16�Әp�/�b�(O�p�LP1����T��Mz5p�p	�]�ʼ��] 1L�Z������klɆ����6ī�pQ-�[������0����n�P�25h�2�|���D��o���{Y�FtL�k�ͱ�r���=�`�o6_�٠2��$��a���R��S�/��e?Cѷ߿�DZkT���ؕ7OV��7����M�e+Jo�ì}9N��3Q^���2��(��7�𬣯��|��1p`��vSǟI[��UT~��E���f�|�v�?�v��ϏE��O옮����+�ؐ��v.������{s�0��Xy�B��QH�|�aJ5v�t�c���O��?�o�G��#�_	�c� #}u5�>9�Vy@���^���%j[��SUؚ��FZO���iH`���Q��?������JY�+�P�E���cZR:�Z<Y(�����!�Q���E��	֖=ȑ'Iz�����Zn�Y�=��;C�F¿�1����pqa�`���bu[�����E���(@I�<�&��@�Uag9�F5�O�$1n`�m������h#��C�WW0�쀗��9�����&5qD��o%"�fT����l/�5�LF��ޞ�9rw����B�'�䮺%@����A[�E��		�f1EbIp��7E"�� �#7��%�*�$���pr��M,�.�4!#��wf���0�!�"�|G�4ÃI1=�J���_Ւ�jkk'������1����|Ha��V�9�����E[�U��+�����RIv20y�޵X�)q�m2l!��N3&-`��:�`g[>�D�2��^�\���6ꕑ�(cs�*T��o�g�=��M�����;��s���fũ�3;��J�a�*��l����&�N��ʫ���8��  �����/�k���WF�$��ڐ��)�o8�t�p�Ii*��d�S��`a�m�3`{���f*�C���7��D?�M�]�����px� �2l53����j��P骽�x���x����(Z��2:28~S�ZB����i���c7}�z���^��[�W���	�>��rא"�a�&�y��5NbJ�ԍ!���cG�ʉ���Q��t���?�S0�om���9���@mn$�x��]�.�$��I�6N����6�t$��l,�
t��t�ƭ���ɘD���!�:���QM��-˴R��˶�*���A �r���'}��z��x��EZ0��2x�s��qiwro:YK���:c ��V,k�^I?t0�H4ŵ)~QF֏B��Q���Z�O����W�ἊJ�\�̽��U�9G��~P���Bu��V��K��(d-	�Ξhr��ntY�����I<�2h�X
��[���B��a�M�[��mP�v�^H�}+b����~U��~�[B�H��,¹��o��Ve����OL���/qvc�K�X�]�Oײ���Q��f2�Y�8���<߫�k���x5i��!àU�?8ySK��T��Z���}�~τ6���s�t�8�U;�A�ޫ��~���%��) �I�/3O���lֳ:�TSᰞqh>���w|S��ّ�0����� :b��c3��RaH��E_�>����<���
;g'�&�&q��.˺u��H���؍.w1:���xg�L��h�Q���<���6���9-}��_���|`�� 0H,�Y�`���c�R}?5Z�.�ID�j�ɷ�%X�����e�t=�i���F��Cw �H��z�m�ެ�q�����I�e���!������8����d8y���z��o�Q���Z��R�B?�*��.���g�7�*���¶�[�s-�ЯO[V�,��omh�[�4q�*4��-[F�hjb��ح�&�!K�HR<��@�u�=��@?
6(a� �n_���(�.�S�{�y���r������M�F�v����+Jԟ�a!�r����鯌�C�n�$�Fl�씋ko��YY�4m;��	�{�s]e���E�"�����˔�ᇱ<.[ݎuBk @O(Dɮ�ji$�6?����d���w2dH}<R@P;$D3`}��V�)�Ч#c��12�x��52I�8�K�Ɍ���)���<҆�z�����m��޻���H=��((������܊!)�z`���~o���B.��ᘜ$C���;�nG�a�����w�Ʌ]]�tR~)�ŭH�`X k����w���ԣΏ�Ae��tZ6g�Tw}�)e�شx��[ʣ��*$|�jy�l��Q��x%��r��Z���ctm}���S���Z�����⟞fG�)�`�K�Ֆu�A��ؒ����w��e�V¢^d��bG�\�>��t���5I�l��Bt���z�%����j��ш��o��ew���"��pߖ#eR'O����)F�"���"���%_}��G7�w#���ǐ
W���p����Rp�%jJ!%=�ʃ:���ג��t_��M)��I].�0ɰAx6� ������c��>ZEf�hB(��׼��z�8ø�a
Wc�g���������Q�k[�f�t嫱���VW�t'�H�Y����%����~��p��R�H�ͧ�J���ּ�)�k�����f��� "��F�[q^�$�swV�6j1�*��!�E91���W�w-���n���兪?x��G�b�/�	��e�W��m�egu�~"��x���μ�1�Z���dqx����Nq�L���K����;��c"�)�_��ו�����Z鬘���l�A����8����T?�\, �k���n��7m-�I��YY�)�8.xf�+?g���~�E��)b�<p��E{��%a	<j փ�a�F���Z�?P��ךRŘ�?���*;
��	Ø�G{Q�M-��P[ˣ�x�U4��wLqܱ��u�$�L���
��M� e��*d�ܝ�6���6���g��(|\��J�_"C��������yİk{�=��.ߔ��i�/��R���k�����3 ��)��??��4��B&2r�_aM����Y�[/R��"m,v� �������ϭ*3�M+�x�y�&��j�j��l)fNf��߬�֫x�H<���+�յ	� �s�4���l��rp̿"�C��h���
*�u?bo`��ˑ��O�I� e�.S�(d��(i��y�B|�x�����O`��h��5���Od��I��r���8����&`&&]�LK����䕽��������4�\R�?��r�(Q𮢟q�G ۢ��_�	_�N+��tIck���s�/�� �`Y��g��<O���z�_���Q�R��8^����>�(=$��{p^N�tV�KD��RLN=i7:K��2]5���V�?;ќ�iƷ-Ie�]����-�*�>e�0r|�7������i��b�7�ë.]~�p�PĿ�f�B�O�͵	0�Ҍm�RJX�kVK�o��MQ����Qn��G2T���M�����GU�n�r4ʦ�<3��7F>;
�n궮����HV�@vn���ãF�0��>ޜ.F�)��W9O!ܗ��'�p�VB>�� �}�Р p��cS�ܨHm���X>��&hw��|*���x�R�_
a��ۭ[�c��y��r��-�)G���#��?{[��H�SYqc���]���I����:�l�O���&R�L�A��߹:�+s=x�MW{� Ko�]p�C���U�&�H��':[�o~�<Q2ṽS$���3�a��l��t��l�tm��je�$"XÎ|	Q�	���%$*LJ���-��ht�9;&Y����р���O/W�9x�J���Z����E�i�/��иzlb!V$O��)�ƙ?�+r�$?�#�ߕ�fX��V90�h�v�tp�$Ō9����(����Ɓ���1�������-�R7���6�"8��uAd��]���+mu�V�	�;�W�dn�nTQLM����
vQ���k�_j,j��(ƿ��oe�?@�Pk,��?��OY�,�������nd&��춍�|$g@E���?�q
�x��eQan��� �H�������%����{k��r*Zh�(o��69�{w�M���*`���0�Ϭ��N���3c��8��t��K}g%qM�^ ����T����=��;A�9yp}]���g��`�P�U%ώT��k`���n���_!e�uf(��¡���%Ò���H��4
r�o�ϫxD��+�"��+Y����]I����s2���W�;2�"f��{ζ�4f����w�)r~4����J�D�~W�Gy7x:]~�VhEVoH�T�-�hz �#dp���k��ὲ=%��~AM�/U#���Us����na��NB�E��pG�C��`+%���@�l���ؘ��;g+s1�wu 3/��K,?� %���Hm��dM
��σ�©2�E�E�I"���fY��Q��GY�r/]��?Nwz?0�S�h.��I���xCB���a2�3�`�HS����q�)i��}�����ڙʆ�F/e���%Ӻ�w�p�nL*����s��?X/�N�;JF��
��4��@�d�zy��Tߝ�����)Z2��r�^X|�y}6+����T��NF���V�n[�I��>댳����j�zL��lt�7�� �$"!L�ƚ�a�[��7+QRw��}�!�6}��D7(kBE�6ጓ�۠���������YĒ�n�I�~����$r$�f�az�s�"R�S�ga(�:����)�y���O���>�QHe�Xj���p�W���2S�״4Ľ�}�a�˚�~|�T߄�Pۤ��rX����9�{�bŅ]N�����g�0xn�f7:����lRj�� �O����@,l��feF��>I[�IV�C��_�h��;W���w��w�s�50�a�(G�rK�g8IB+
�;�
��_�a#,v�F���u`?�j�����0j}e�SJ���b��4|)����Z¾?���nQk.HN2��+�!���MY��ݜ��������6����FѢi7_�00�NE��ʕF+�/ITx��j��A����*�-�s�K@W������Lz�h���Kh����Z�$��cG��<W�;�Q�̸7|p��E|��ȕ@!Kѓ�"�f@j�v<�	M�I�/�0�6��_R�ĭXΑ��@��2���N��U8��G�lh.���Ǿ�7��-�X]�������f��<�\IXq1�3�sb/�po�0��!|�e��7%�o&���ի��I��R����/�� ��A0��z���I t@*�`�ݐ��պf_'����Q����4��]0.S ��T����Fe��ȴJ��Ek�10�'�h����]!�ظ�)�*���'������͚&U�eѷv��:����%k!��Զc�#���m��[�١8\�2��V<"��,�_�<#��Ԝ<O���P{�X��>m�g��C�2ix�fO`~C�0�BLj�qccT�.�o��N���K������d���odi��m�a�:����-��Ma��g4���B���NNKXh�l!���� e=�^�p��ם5��<FJ*���A�8��<��b�	��Ƅ���B
�E�?J���!O�h�H��b�u+��֜��יY#�����rQ�;�Q�6��Ia7�
l�_�F�W�*W�R��UW�
e�U��q>���p�i�t��9)..�4�EK&��mbgMQ�z$"�r�Q8T���a�d�	�HD��缴X57�oe����Nv��̡�<q�4i��a	��i�f��B'���⌏9�%lV�nvct�5$���PQv�y�9a�a3�����6H�e��7,�AFL����=���fls� 2/�l{��;�����O[�w� @�Yj"0��<}�[�K��O,G���)��,���J��4����,F"��ď����E9H+�����Y�X{�m/���Y�6������!e�ƹ!:�νx/C�i�@@!�{�1"�T<"�^���ӑ�����ou,!㿫Z.(Ry��v�yf?�k�y0M���0���q8����r�uQK����Q3�Ge�D.�b��!�.��ќ���ᎅ�h6�]��yI��u���� ���]	�ue(�O*�}s���F�$:󢙤���p�,�.�GD~�"��sS�F��`V��x\�����V�n������v
z3��0���(9���l��H����u/�+�ό�kX�R`�o����.`�/����E�Y��}�����I�,�
R&C����0�_
w���<&����q���ߪ]4ݲ�Ѵ�i�|������x�-���A����G����R41ʱ~���I�5����:��L��~jC��r��?
����k�h�FU۳� H(����=���֔SŤ�Y���@���&~�{N;�H
�3�(�P�Gm�q�e�(C:G����4.�d���<��o�~��kÝj���/�%�+͠���)�9��Vkl|���'��;�WO����{*�;��Snb�""��Ύ˿愐����C�V���[j��w5��FI%C�A���q��E�F V"Y3b�F�v��`�|߅�%J�j�F�b�0d�38����]��Pn�W���4�-�K����c���=__5 ?r�6d�Z�b���7�����M�j�<�ר:03��%���A��Tp���k$�ٰ|\���|K��X$��&�R=�y���JY�S��i�P�2��&/Q���F��j����% �m���:s������8���-��`��U��Ղ���T����;�V�u˪n.~�I��so4�X�t �o������p|��
vGg@��v��loN$v>B˛_� �m��wi�I$=:�����b^ʽMa8�y?M*��zK���C�e~�[R޺�7�T�[E[��֞{��:�9?,z5#�E^*ԑ��Wq�=k���庳��y�1VQʶ��(��3��oL ���W��K"A	���q�^y�VW,D�#,\D<l������ ���ֲҞ��8���K{�f�>���=j��hG�VJ�3v_L�A�=)dfS�gy/��l�Ԉ���s*]1�<��4IV�!���.�l>���jS��;��Pw[CF��6b+v��u��G�ܽ8Q;�Q��{H@�(!������I� �UP��u`AN��{~�'Nl��+�{DH�.)�2�Z)&���vY3���C�׬�|5��v�C�q�ç1����N]@g�셷�ʔ��޸"i̬R���^������G9�A�M�pUTIe��D4��]�(��gHr��m}%A-[��b̽i�Sg�� K�Ŷn1���kI��������0��b�D�0����#mxR��4���%�
�^���e�'=E���,��ߗ����;�Mg�X�6�oF�Y؜d�R���i��ē卆��4�R�5��ͫC�!�|xZd��V�/�	Ue+���d�N9}~�go�*n&#X(�L��ӵ��пUmƽ�˕��Dk�~o���K���G����=�Yt�T?�ך/�v��0<��ym)��)m /oEX��Y��iϬ��n����p�_��QP�Ck3��b�T�,hũ�T h��ps�zž6�����
�5��F�E~^�j!���t��1�csh0����Ѣ���R���N�/B��'>g}� �o�%����!)}l����җx"sgܧn8� �N���M`Ui���E�+\� м+��Ot���I�K� �4��Xk�p�2X�0k��y�!��Z.8�Ä�TW�i�����.�\�+ǆ� ʽZ�����H��ΚR&h]��#����Xd �t��wy����0Ļ�#��t������kr^�ie�O�+3����oP��ud�_P;	J�	t_�:�����ӯw�q��'}w�@g���������e�ɐ���Hl,Xd��������~g����
t��B�&�ƿ�Dļ����%�dͬe����q�^�L5.I�#�c�;���;�WU����ڄm�v�PU��q��?�[�c'}�|$ �ѵ+��R�n���`����E��7j�Li����ʩi��D
?��(��\�D.��7����I���MfN�G�R�Y�7b��0k(PC��T9��wR���q���r�j�{�����M.���s�<�.���K�
haD����ː������f���yy�Q��R����J�^�P��/{�e�؁\K% �ue�Q��V��L`8�f���͛]�v�<J�\�^]�[�
�����AZ��$ �:���tuԌ���#䒔x04Q�6U{���?�סQ�����m� �L/Z�3�,�͌=�."��ג^���M.����w����di��hӒt��4�s#���j�$Ƅ9�]�!�µ�;�8;��$��xRdn_7<�Kf3V��_g_i��Ug~�����@.���a{!,��J��U /;���U��6��Ӷ���[KLtYtgW�=NXX����`J�껞�h�Y^����Gn���N�>n�]�����E`��T_-"����%��_�a�/[BM�[Z��;�ѷ¾W�f�^ͫ��NEN��S�ւ��q�V�{v�j�^�Q��69���2^�u�@�F�i��	ra$d|���������֊�w�U�����'� �� �0q2�b[�Ɗ��r�U����m�6a BG�#+{s�sD��'�	�e��]$�b_iĒp$���9к<F�y����uK[\���\uf�#hs�wB;vhQp:���mm$�x�RG�	�{>�Z\��]_z�r�z���?
�*������{��2�>E[����+=�T�a�,�;脥'� �={C�zi%�Cۤݰ�b��\�R:>�E�%���t�JfQa����� C�m��#;a��F�h�Bl(8��u�Wx�Kw��Ib^^�(r���pd�	�s\�2��c(��D����0���Fr;��,��MO��[$�7��7��a�4o���lli��p�=�g��Um_�aJ�`�?�mPf�\$��!�E��P�Dȗ�ĉ�O����#`Y��ʯ,��i��-�(E�l�Ч�vA'�(}v���x'Zq�m�5D�S�)j�9p��Vt��Fyj��IHN�A�2s
�{s��JT�	W�l�?x�������r�z_�)�V�L⛮�H��5���(f�`����bf2�zc���d���@��cK�������c�XA�i���K���O�M��b��������9�*8z�-���o|��4�Cj[�����x�yCħ{p��y�;�|�5����j��Zt��L�� :�K�ӻ���Ғq����|K�N�^a(|�ƿ}���,�j�q��Z3�  ����ɪ��Tq�gb�u\8V�Ά�/�1�NQ��\(��=���̶6[�����È7�}a�a1���{�
v��	��9���ڜ������ì���6��h� �z}K��N{��K�K����֬jsӎ8L��2 ����Ac��r�ȑf�Z�F�b'�tA�g�+������h�u@ϧ1,CC��Z41��w��{%M�GY2N��ݕ�
��-T��y�ܾ�&�k~�lR��?f��ϯ@)��@�%�z��8imϨ��������.5�	)��S��㣚T�����sʇ�WI_�*f�fl����Z�ʅz=v91��Gϵ���Y�}�"4`x����%��&���S����]�	��R��)e=p��l��XCX!�};v�A(�@ٳ���,���̍��d{h4�*#�D�Y��+JreqU{+�i'�*�����-2�7)���N��/��gN-$�k ���w�:�������Os�*^ư�������A:�9�����xS�5&�,��v�chg�l��K>Y�<�K�j9��"ޓ���&���ԡH ����0@hX ��[�b-�;��Ra�=�
A��]8���j|�b��IEH�R~�T���l�_���ST�:}ke�O��Xc��������ZnH���C�Ndv#��<��e���-�G����E�H�r%tZ`���_
�6u�2\���Ճ��ε����9�;���>ԙln�ZB������N�_n�A�<��֡Վ���e�D��t7q�~�SI�MZ0Jǫ8:���c���M�:�֩xQ*~ؚ�-��L��n�����Z�L8Ħ ���Cݩ)����h�]�����W�XHy�6zZU��Ew������;�,�t��8B��+�0��(϶�,�<y`j)���(]������59��]��7�e���bp���'0�T��y�T��1x�s��a�Zݻ����9�S�$,%|/�Xk����HQ ���yy���\��8� ���� �1uX�0㏵�Z�k⪠�k$��P�7����9��]���'����ɝ"�%��s#q��F�vg�K�<�[�K E�0�h�oK�9���hzqx%9��|����������5��.��}��G
^�>w��Z�8�j�D�*ﻅc�PcQp߈��d��yF8a�.*��ҎBX(ˮ)��xa�������=�f��6�6CE#�B�2�Z�AƐ�h��}C����aC��W�Z�?��i"p��1J�=&&�|�_l?&U�cޡ͜iv��]c�����|�G�>�6�Y�M�c:H��C�y3��7��-&����V̀��"a�����qs=�*���i�G轴�n� С���g�b
J�H���0�H;�����ozf|�xn�
@j��P3ow�7�Y�uRJ�Xq��ފ΋h��� 7�b�O� Ǒ�A�>n����=,���:P ��L=�6;sF�x<Q�zK�`BV�ϡB|���߸S�Ӎ&����)|�Cs��C�� ��i�Z��g�%��l���8���}���J�ӷ[2���E~4V_�?�X�����urJc�T�t?�wFϪeU����Z$�K��X@��#���?��c��s1�땽��i�O�1�Um�}����Y�jw�=���'������aAv��l+��b>g*�=�bY��*sX�?E�N�����J����k�7���k�p��dg�1�ݑ�3��Ь����F�:�z�p�s3{��	�v��c��E|N%+'EG(�J-�Wա��U_�Q�1Mp��?6߲ %�f������2��´&}��{�pg!���R�s}�.���Y�����5o�ȋ� ��˚%'�/����[��#h#��N>�hc�)��2���YBt��S��$5M4���K����$i���:���V���ö7�F̠�e��[g,���T�B�l���wa'ڋ0��H�qB�!�bO܁��>�-6h�ATm��v5�g�T��5��M(jY<�+�&�,��fJ}��1�9D�p��G��l,������+����ѢM�����%I��Ձ<��MT��z�_�BH?+"S� ŷ�W��|��Ԯ?��?c]$۬:~�b�D�@عhX��� _�p0\	���SY���ڧ5QB����4��Xf8������o���d��V����s�t��!Q�Bp�@I�|=YdDE���b��'�0J Ȑ�3R>ci�f4�D�d�>r��a���eOh1��F������j��E� Wl�#�ci�կl$^5
�d��A��A۱~�;-�\+���k�qN�8lqFK���t���\�!L
����] �fꘜ�w�>��(g�h�S'M����(���0˩�3�˧�ߓ{�|���O��C����B̷��}nv\j�c���f	�^`�1p��{f2������]}��eŰ��۬f��j�H*	��1]0@t��Ї��3\c�A���2��e](w	�K��y߱ &
�u1{� McI^qwTCJ��_3��)0��F�a�z��;��[�� ��3g>���\B�t�������=4m ����3Hwa�����Rz��#���u#��ʛp}��R���b@Ƨ��I�u{ʥC�ؼg�E���%��5d�;A`�� T\\4P�h��#���8B�K �ϋR�2�q���)�����£�e�� ��D��8�M>6;݀x�ξϮ[;<�A0t���}q�D�7�0pF�Pu�']t��ρrq�/ְ��g�E�K�@��z~N�k%{\�8P"=���)�.��G�#=D�U����ۖE��|�BB�����A6y���a�"u���5��ow#=Q�Kn�s\~�%�^=i|ͪ:�7`�4�7�i�q�3	��'p]�F�!^�$%���C<�QC$����O&���'���O��觱�j�աP�S��n�WML�\T���'?a��p�=��;�A�����y�����63zXH9��Q_�u�@mf�f�Ʈ��'�Dϖd��kB��S�����>���wZ�v�a�eVgr�he�ކ����s�G���;x�����qMg0&�r1� ���V���b��.Y���t�z% �����\�R�2���������,�c6�c:��&���ͬ�֧EFU���aH�a�����!`\��w�w�Z������d�ztjZ8�t�Y��ʩ��S�7�dA�0���\wt����ԉn��bo@uw0��M�%-��=��4ƹ�QA�ne.0�{�ɏ����g��m&�'�H�;7�/����5F8�%�Q��.d
w2���g���Y�P��yk\�6Y_�~���s��-;+}�]MP��<.A��k�����gϴ�����qݽz�}20Mi�G���K��1Ç�8
�c�"å�(����8��0 ���2��w4�&^ I+��LX�X<P������Ǥ�$Ɩ�x�W�	�����9ċg��藎@N���n�`ʵDv�#^"�"�\�u�V��:+�Hk���w��f"��E�Q��Ʒ�a�W�#�[��1#�$�v��ږf��ё��֤�N���௱�.���g�}x�̒��R-�����l�b?��M�b���}�U�R�|���־�y���� �0���V��k�U��G��-W}P5 !��?J�@�0���:�9p,;��� �'>B�%��>�ڭIy\�Eä�%���cDv��
U98hvvpC��z.�~z6yY��ԍ25����nX7�5�p��8�T_�N��(_"8(C��@�6z�3T0�o�S5�M��;0���Q(�c߰'���n�uQ�l�w�S��-��t�M�3{����c%� 6ܡ�����H����V����E�4ӵ^r�'
��u�P����tp��j9(ک#�m���a4%�v�j�2��۾�X�m(p]H����g�#����槑�`F��e�e6=!x�^���
 ۥ0��<!�D5}�?��\�C�?q���A��m�y�˚�Z����4�m���&�4=/�sg]Brq�L��4K&cL��	��M��yYxv�[�I�.�&_�<�����XH�`YS{z x&�	��C�iM�����a�!�%��BXd �tΆ�L�ޚu:?	 R��y����2dha��.����yލ����&�!rD�s,��a�"�k[����B�����l�G�2^�1r7�Ś��w�`�����2��Ϫq����^�M����Wk���`��l�;yj
�I���\��9����U������l�$dɁ
��@�K7�LO�e-X6X~�����Ϛ�q�!��\���:�[Q@�e��BW.����S%!�NJ��z��Ԋ�}_҉��ٴ�f^��_�R<���?����)�n(���b?�!�P�CrY-Mk��S�f�Ɍ�DY��߫G,c��|1E����H��*�,���|r�K{�rv]�x��U�\�\a��K�?�������ߔ���Z�.�]�G�4���A�� ��į݁ ����8�2zTY���@�v�"��]$����I�m�Y�U��.���	u
�uOc�r��%�	�ʪ��Z}x��Hn|�\�������n���3�Ó�H����-ꨬo��(�wϨd8s�K���\�<��Ϙxk��j��L$!�	�o��5\�՛���dZ���hN��mo���I������M�E��]C3d
-d�2��i6R �Za�Xۻ3����7]&��j��\+5�M �d���{�������s�䥚�
ks��U�O��]9��9���_(5�s?��Ξ�=�]bY ����EV��L�ilqN�u� ���nTb��6}��a��/��qEg�I
-�Vs��u���_V;�xc���ACe�F�$eR�P����f��M��`x�u�D�t�<��_F2�%�e��U��x��
I3���zT���P�av�&�%�e �uP�5d*j�����F�}Wv��¸���Xcu�7X�Y-����Kp��0.9,�M^�Ev���ܥ�/��.P�x����bH64	�b��q�|:�O<���i�<��۝|N����\���Qa��eO4SŮ��ܲ�2���S4`�>(�C��0Ϋ�y��qۓ��3�W�Oi�x�
7Oo��9y��r� ��K���H�*P�����?v��<�	 ��̩h��>>x&⍪���4�%��ub;�T��ߡ�Z�f��,�W��/�s�Hx��5j�`�LLF6�"gˇQp����%ϕ)ki��%��\������Y�b�yK˜2r�i�jX`�ꪋ��DI�V1'iI�����pC��ԗQG�3�M��gD���w��矆X&=�94��,���r�R� >}�
��=��e�4��n������7����J�y&H�P ���}ڈ�"�;Y[:M
�o&X���M��o��@J�%��g4\W`rQ�O	"H��OS��r�ϗ�3����9^0Ů��89��Fe����+��X��GC��;�~���<Oa��-�I��f[�]��Vᐎ��܈����S^��AҼ�`Fڈ$T�>��O>��i�a[��(d�j�Bm�˥�VZN�
�{�F|zW�~�|�v/7�ޔ-�c��,{sZo��h5$=���zs���w��
�����_�5�n�/��-m	}�~�\\��H�k$�lH��7�g��=s�3�󔾆�K�t�v/6�2"U��QpZUE�Hښ-W��D1��C���&�n���Ԇ'տ$^E��¢jW�m��U�6�D�p�YK��V��,L�h0� 
��3&��y[&\�3f�.����7�m���xzSq�ߠ�b�F�	�� ���� ��/Ɔ^|�=�"3A��C�]X/�Zx ��L\Ο@��ng����x�:��q�>O��2��E�ZBYk�BH_P�k��{MKd���� -�V�F�o�i˚���g�6��[�����&-��mO�p��6�q��*[��0����2`�,��6����4X���7��U:��u���i�N�qu���f���ک�G9[Ӳ�&y�v����D��܎�q��V��ω���Cfʊ	7a��y,�>Ҷ�wg�Pi��b�>����/a���[G�p��!sԈ��ޘ��,�B��%\ɩ���4�gw�x���X�/�y|���JoĖ����% Z�G���T�^G���v���f�?�]�+�j���nI]��:"��P�0@��������[����u�#�
O�Ű,2)Z���kS��\m���/ˤb��ɏ����S4�L��=f|k܊'>�K���z�$-
�����d(? �a26H?���������S7�vz��=1�s�HFBHMj�=��*�u�Q�p�؟=���c"��Ō��{\�]�yiȶ0�u?l�,�8�s�T�v3T�n<�.U�C\W���ыf�!pN%�}M:�I�~c)V��5(�d��(6F8Z��@^�s���EM
��q�F.&3Ϝ���f�!�l���� f2��vO�՞M�ƫ	!��v�SO'����Ǣ���?H�x)3��R]!�v��$�Ytٴ5����P��,�N�*����gI��0Ѕ[���fX�{�G�Um����ޚ��lY_�[x��{��㛞@��ɳ#�a��/s�����ph�k)��d�	L�Zjz���I�Y�%�
��R���ڲ���D¤��ɬ~p�ȹ�`⨅��hŴ�rh�P��}`��X�f�'�'�m;�NkK��,�rޡ!�^)	G|�V��x"F�T�?��r�gI�kl��]���@Oz�VJ���8<�̺�<��f-0N��e}�8\�gр�|���C�@G�Mڻd����o4O����m�f;B��<�Ѯ"䊃���Q����q��(�,>��b�\�x�J�_���[��hj�����74o�|��I�0���0�M����3��F�� ch���\0`U��_��_{�*O�T�^�ʧ�s!]��-��u�O:�ל�=��]~�5A�"��Mr=!-�ֶsp�
�Y��ڏ�j��u��L���i�)�a/�i xmlSyvrB�E{��?�p�Aqb(��V��l>�43�Tz�3��hQv5M*�'�][����?��]���H�vjA��*��;���Ԝku�)9w/MOK	={ +m>}��=�:�o�n�2��z�4c��6�>ˋ��2.��$�4v���3�׼�S�ֺΐ�Knt����ǎ����� |�+#�+�9u�<�{?m��s�@F�D�3��ͣ5t��+V9��'��dI��υ�k��j�Wu�v(�b��A���w����H�����zb��mq�;S�ƚYH�s�Im�iQ�/(�4�x�ߥV�E�o�g:=r����q:�X.l��6&5�ĕxW��G�fC����_p�����i
���� e�w"{���XX����ʘo��qgі&�M�?s�l=���۽���c����B|���Ԗ��d;�5_��b<����]��#,�$-�(=��/�lcRx͘[�\��� o�;m��T�U|�\�C�!]껪�)|;=6ʄw��%�<l��	�~�<m�Pi��-�⪣��!�""���圲�؏�A����Yګ���c�Iq���BY*Ǣ�Q�:�/�ʦ2��:W�sR�N��í�)��e&PeU�(F�G)����{���XQw@dT�'���+��Ug�&��#�P��Ȇ���< 7���"����A��jD�3�m���Y���#}~��F2����)tX+�|I\��d�
�J��ؓgr�/�(���������( �P��#j��R(��z�շ�����H�3��,��>�7hϟ�erI�N	^�\jSc��H��G�y�]+!OF��c���߁Tq/�1�4H��*$�l�[z!C�A�����++~	�2�4�[�)5��H\Rq�t=#��؞�05n����ň�,"̮% I� (h���5޻��X,�藨�mFC��=�� ����K����q��������$xf�f�N���vp`�@:D���·u���z��wU��=5�H>�� ���p,wT˅�>ߣ�	p�r�+�D��g�.8��ƻJ|�8tJm+��)����㚂����FŴ�=�h�B<cR]i��#!�sv^~\��R��#���k(�(,bKʛN��=��5ǽZ;�E�}�3fZ���e��[�1�p�-T��h8��mq��t�u$!�mDBz�g��=E�5�z���)띵���u1��&��[ߣ��R:\Y��.���_B���LZ���%2L#s�B�Y�6L��.��܂2�Ӹdǝ�Q��6B-Cg̭+kp�f�!� g4�X���S���ie��>dn�L{��m&�R��B��i�-Z�9��,ZU4I���m���e���jC�Z�Su�-��|;����T�Sd��kWn˲W*G����n�S��{.�]�Z��zo{�p�|wM�s�7�2	���xL�������1�Q�%r��b � n��y.{Sx�z�Ӏ�;��'�t�5�~=k�zf���sIfs;u��*Dh��da�Uf��Dd]r�]����O���9뼯 /`��=�9���]����l�!�'��~(C ԰&�"y�Z��C�v2b�� ��)�Ў�}�4ƨA�!H�^r��/9�r*��Ź0A���}�`덶ک�X<��M,��`b�f�n��jLk�xPhIsCu�3[�{E��B�d�����8�����!�!��o��Q�M{��D�4'������%a����5@h�!�O��~������FƤ�O�gV�z͍:�g�I@"�jv�~y<f#{5�=<�L����ML�˄:���9�{KR�	�-$��G�b�s�9���;)�d��<���w�0��X�,���G��)INr~����6z�Y=E�7��-�AZ��'V.���aڷ�Yd�X;��2.����s��� k��+���0g�B�#$+��(r�G8YMtR�g �{�gg��!T�M�V���[�6{�<���^?�<��s�4��}�U�ZN��H�4�V��!s���U�9[{�����QP�؍��`�^�Uw���-�W/�E)�����sY�L���6!g�o����
(OU���_��,����l�S2$�������ժ�v � o�`72c�.�f�Ɍ����U�)�K���^^�����o0�	���t+t�Z�.�c}�f�ȚS�@�c޷�� �7�e�(6���������f��X�!|ĥ�C �K��E�l-�h �lTt��['k��mWQai�ʽgP{��ε������$vWK�<�g����j���/�IA~��5����֮k�S{�te��@ӠR8��E �)����P�gp@ڛy��t�������C�Z͌��=�E�J��"Ν-8�%7NGu�S{R)���OrH�X��K�X��E7nT�����L���J�/(�(�v�U��N�`�iqEu������	�����T�F��B�3.��7�tE\�T��L�%�JR ��C%�(!T��t #�v����\���a&����?&�r�V��!r6��)h�����h�z#�P�0�}jo�+`��I�m����;�U%��Aq�	E6�$���0��W3E��������*�M�  �AC��{�Y~{�֊ؿ-G/k�3�-�+;�3����Fɳh{�x�\#�5�0��6pn��T6�$ժRy����u�;~�X���a��/ B�������P���Ț{ӿ��^#_�/V�M*��]�^�M�(��G%�T��ã����<a�8E�0(:(Î!>Q�X0c��r�WꭏP��D�6Ш-����f(0�ئ@d��>6��z�W�v�)h�6��.��S�l���3��k~E���:�(SV�	����RSs=���nD���dً�l�	�r��� Hݽ�%_��
�4t���#��Ra��A�kU7s��-�J5�O�ݒ3�=~P�0��8�#>����`�Uղ�������&��<1,��$3r�J�"	vZ�������\Sp�z���Tݵ��ڂ�,s�M8-����\���9�:TN��-�Do���ƕ��c�'�k�;�/�
���g�������� M�o�Id��Z}��T��@7�/<wG�vgO.�F��v&�lg4U�])�6����1F3���������}Jv�^#�,�)F�F��b��-��hXh�!�U��9	�T���#a;��N"��O9T�5*�G^�7�t��l��m��B���E��m(e��#?:*��zG� {D=L�1�d��d�W(,�͢��י�RN�5`�������Ē�#v8��z�T��D�����~CH�^	|���R̓�ۥ��q�z�o�����tC6[��25�d�v�n3?�/� �M+�\�y_�UxO L h��qJ9lR�s�M��������)Vۅ��p��k��_i�$[���&w��W|���1�y��H��^��la{`[G�$I�s���P~�+N韦�7�nh�=�I�ґ�"���U�۠,]T�!�E����qX`X�?��1 DU6����D�ߕef�Q��s�4��|�PJF��z��n���W�����E�D�g��[��{Jg�`�q�%G*��df��1��wS7mWhG�Sn�@~H�#|�Q��VO�V�!���i��k0�zȹf5(�C���֬�L�w��;�|�)LNG���"�2�/yr�&q�/�v�WL�Y�Ew�el�	�&�A~T���F6�r5>y�&\*��Y�f�+�i��IX�t�p�y.��r]* �(������Y�x!�dvE�����%<�t�gsg^��ŭ�rjb��I>���ޅ/�'�|y�H}�������i�h��ѐp`�QN�J�F����Y����r���&)��ة�:/�3����w��&1�.V��쵉{���%NQ�ډb�PEg�d�䇸 `���m C�rݯw�E�0�K�_�M�^D�wٕ��h%#f�c��(��� Ѣ�m�F�7a\��'�wzJ�r����g�yZ�p�Q_�R<1���"�[*|�YQt/����ϨH=j�.񰴁��O5(CC:M���C�+�{����}W�G���Ǡ�~��]��A�r���E�Q���N:u��#�&(�
���O�*�QG �"������*�O�@-�p!��_�Ң�4�$c���xYކ�F��w �&�bNӮ�}u�>4����C��
���'�=tW��W
��O�6��vR[���0jG\��c�a�q:�ު1��֞W�O�J1�fLI6�]�9ْ�Υ�k��EL��HdY�-P�ނc���$�&H��,ut17)Ëqhb%�|1ɽI(�ɬh?�Ov���/LA�,S��'�T(Y��_�����&FM]C_�w��&����M��JL *<y.!]����,��ٽT[1�!����z�B�q�����󓽴���Z�Q���g���1 �X��h�?���7|���6��XT��E���)���,l�y&��:���{`��厫0
�e�R�.Ϧ!�!��ԗD�G�,O��᪫�&�zCE������`6��dqM�J%����v�7��@����|��A�a�n��g��~�kU^�_he+ۇ�AN�tTg���uKHϦh���3��@3ҩ�����a���e�>���t���h1��m�T+�*2�	"�*eZQ,�y�n؟�0P�v!�:�T%����	��yx�>%�Gl,?>0��ql&`��4��C�u[��<�[�~���\��d��fԄ�
>A
��Ǔ$����Q��9��>���,5v���.�F0z�	jҧJ�y7�8-��C���1,�|D-�0����ϐ���{���h���-7��I>��s+��{ߋ��d!���P�:C�P!��t2zbl�a���$�G�4��tt�)���8j�CQh�_?w���X�������؝n�P����N0C`���K%���}MS� �_>E�/���5b�y[�y��g�*�S��g�1�G��s�.OO���� <�`�$����W��ͻ5*�����ż�m90�@���l�b_�+S�nBm��P�5,MSl�VY�6`zl�����lwc:l�u���I_��v�y!)
�^�P�a�{���P~_S7��$[�sX�Nw�����c(���j����ldt�Ix+�w�(�������xU.�^N��	J���T(1A�13 Ĳa���bD��������=�R�E�l	�`���SC�L��!\���}D�����2eS������u�٘��������y�ssu�y��C�o��~�}�u����WY��. �j���^|]!)tJ�����ϫ���&���� ���P�J
l$����Ȁ�o�� NS9��o<Վ�����.!]s���<��d^|j��?ϴHk�O$�H�Gn$�!*aG4M��I+O�U�l�D��4M�I0$�41)4��=z�T�8@؟׍����$�g֪��)r`VY��J����J�� �h����O�	:��:�@�5ӹ�{2�4q�/b���Ԃ�gd�M��r"g �U�z$���� ��_�Su��h�B�ĉ��{<3H����Y�X�&��݃�e3�P�o(Cc���0��T���u0и�}-��v�XqϬ6w5�~�j��� Sۊ<��3#�ݰ��։�X�u�&="������@l_������J�i��eXH�6D��o�
!��J��&Rb|��=h`�g�����x5G[މ����E�6���OV���'�G�2��A㊾2\��9�L�
T�3�G�~k8ȏt��� |��Y�U�*R��;8߳�������M̜�� ��M2ժ/[�`�-$��g����>2Y����ɞ�sm�y�R����f� �cea+fIh�ralH/-��Nc��(c �և�>^�Dͫ��Q,���n,i4�gY����IU�Z���ëY�2Q�G��G��;��WO��`�*$ `��o~�p}��&;A�8l'#��cٜ�Ow��	$[kD%ɍ+����ׂx��l��^3R?��i��z���U��f�B�|�!��P��w�a�Q1�#��0�I�s�jX]Λ
��YYF�G��8��i�ŵj�����E�|(��K�n1�����U������|$*s:���ޥ����,��Z��LfG�Vӝ�O�,���;`�ߠ�q�J���ٷ\=*�^�N^ݿ���>��!��}���N�cڂ�;���/m�&�X��Sh9-(��	����u�����ϳ)u�����\�-i���W+���<޷���rD��-���AE"�Jp� �E˷(��X��A\bj_��Y�bxO0�Zs�>{U�s����(���{3p��:���i���K1����\nv�&�7I3��UJ��HD� ���~����T�?zn�(�a���N�F��������M�Xc��F�;L ��t�!�i/��5�;��F�aծ�Y=vs��шs~=�)�J,��td��d����=hjS�P*���zJ�o����sT�{h�����l)��0��=��������uđLUZ����p�B�">�������u:Z�^!�qcɥ�#�G����V�sѮ�~"C��M�+7[5E_��6��6i�KҎ*r)v)>�:	�%OԆ	w��ML��tgzr�U=l̈́�ĶR�,���0���;B���
�S�D��sa�cت�����j����\�*�Kd��!=��i��b��	�;����K��������b�.X�G���yv�{�?[�=<yO�dx�╷�Ekq��X�{8b��+��a���ȷŊ�
N�d��8A�.���������q�}���ps����#��{׻���I��T�i�"�+�����a
58�Y�X�<ac0�,_I�״�G­Y1��^�ci���6��|ʉ�t�P���G��e�Ŀ�H-Qz�6�s�h����5�}� 	�T�?�E�e�ܭ[ ��j)���i|��F-`N����t��,�����U����Vw�_m��[ܭEP�O�?�+9��;.�Q�����b��:g:�'���^�N6� 2,����.�Y*�F���ll!���A7ė��O�HT�f������*�8`Cn.�Rǈ�EO�����M+}�Z�������=�9=��Ŋ��T��%�ϥ9����0�*<��Ɠ?� <. y7��&x_ؑ5��t��L!"-i
�i ��4tL
4�y3�n��?�G���� �Y���a8A���C� ��g ��LE���в�9k.'i"�]��/�X��͵b9�]�Z2(�.�^K
k��D`K�!��O!y^�� t���d�eKP�솭���v�n\�����9!�������e��Y.�aVFe���DǤ֞��p����&�������Ub����υ��|J���� ,m3�����>�5�w���I�ƒ6�ï_���j&���40��̲r\�-�$���E8��7 �Kދ���z���Cf�^K�>H}�M���Ȑ_5�'���;�d�K�u�q�Q���N�Z{Ss`���맖/���\݁W IxU�΁@�o!0��|y=R�!�Q%eϘޔ99�7 ����B�@ŃK�&�'F?�g�%�N�n.zfKp�I�����8N>r���7��fL�U,c��hm]�?�)�Rx��&T[�[�ϩd��t#�0F�	�^[i��s�H�㐵;�) 1y|��Z]�1�o>�eƒ0U�=���Q�� �ϖ�N:M��xuk���TZ�H�=���CM�š�[ư�=<��_Sf���K_%9ѻ�]�V���Oÿ�Ѭ�Ӈ=cz �NV�i�uP�;�N�N�&��yǪL�3G�2����CD_o��d
\foJu4��{}Yx�ɪ�2���׮W�T�cLv �ki<(��(��������_�wB���yC�B�ި����'�D]�`+�b����1B��p?�:�oS�T5����E� S˭�f��̴��9��q�ߢ����д�m�b�~���FB�����hWg����C-�8	�"Re81;�ʸ���L`=��+O��p��ue �d�Eկ�L?ci~�����;^ߐK^�e�'	5+TV�'�罌ڝ_dQJ���ā䅗��?#�\�sߎ�B��,�*�Z���j��]L�K��,&��ߕ��д��k-nj�������P��� u��/u)�`5���no����FU��  �Ȼ4 _ �?�ZYt��7BV�Gz$���K.��_��.ŏr�+ ᘡ> G1z������˫na����K����a�u���f����G���k��͟u���*�% YOL]��%�ӂ��^?ey�jC���.i�xԸ�i�M���4�PP#TXI��ZGЖ֠�t�(2�Kv��ģ��	�bJ��Gs�ס�ù���`P��x��6��LI���Wg�Զ��C����[j�2Dba�!i�ƪ�L;ѕ�KHq	w,I���k�����f4P�g]����P=�4��\����c||�|%}��%�@��H�6ߤ���:��]/�L��q�0}ڳ~a�����c�� ��\)�zҮs����n�e}j�/��kE���:?�FA� ��0i�-��]I좎��!�k�2��(Gy�j�2��z�T��;%���v�z��\��*�4[�����$����&02"'{�_=�5d�Ժ����y2w�E�ӗT_�(�	X��mJ��HG#���VC��e�'��=b@r��NN?ᇉ)r��V,��S�nK��:�"�+��o�"�,���`M�L�{��f�%�M�����2{v����S\�p&.���{ �8������>~iKX�O�Zqx��4�,Ο�%�a��ץ0��Y����Tƛ�%�q��䙥7.�.�y�ˍ]7����Jg�E��&��f�b���g����a�g�k�V�C7�3��:聂N���'��������v��@hط�:t������r�7,��[	���o�l#�G�z����@�/���q܄��8�aW�av[28r�h�/�3� ��#zI��.N�ʂ�:x��[6�w�Z8���곖 ���}�)
AzKm:e�Y�L�������`b�˧����sp�����` ��+��\cdf���T>�d���mf��������DMb$�oT���/1Z{e���jMt�+�.���R8af3��y�n�U��#|��E��{��E1����#���I�nR��� ������I��>���@�����bd��th�<�أ!$�%ն�Z�%�׮�� �8BЂ�E~uG����?��a�"�v���}���#i����-� ���n��F�<��)�T^����V���]�:�q�
tn9����r��و���>�P�r*=qi�|�E}d=�yM6���q��=�a�Z���go����"�'�Φy7'�l�
q�(�q{=�+|;?��2Ǹ��SY��M �?�Ox\���hu[K[A���"�	�coi��y9�am7��[$�Ј�^Uÿ�]>r6�;.���)��~J�c������Ѽ�z}V������|y3r���i�uV�-"��a����>��z��^��w0�Qh<r�c?�}(M;)j����_���z��b[��æ=���6%��](z_��Ju?CB�bR]��Պ� 	�{��5�@1������_LL!Ȓ<㻮b!3�t�E7��h}"�e=��,ࡠQ�".�˴�<�(�+�+t[��Q?����eʣ���t��@���@�����9ಃ]⢖��$;���@�
��UEV.���XQb+(��_l.�x�$� �>�#�f�Co	 �����ioo����ga9p��(��K�B����&G��;��d�r�5��-���2"ܴ5[4^0�B�
� ����D>:���O��\�;޸9��r���/�mi� O9*�	�D�=�V����e��	����@}f���* ÿsP���1
��zJ8��*�kǑc��l��Ì�]L<k�D+Q�e�h�}�R<&R�L�L���W��S|&F!�u>jn3l�\�I/�Q#�1�|��,4(��2��	c�*�q��pf
�k"�t2���\~!��n�w5�|��r�)��0�ҭF�\�^�	a8}9���6n\y�d��S���	������ǃTU���Rl�T ��A�)<���V9R0��@��VԻ��OK{��7N(��I��+W �x_,-���'g������Ox~ɸ�j����Ln��JEx���9�����T�:������<k����:;�v�H�Hq���?�6�r⮼��Gw~̗�Q��ˇI\��l/�m��KQ`��ѱ�������ǎK��T��2I��}Ilj�w�w�",���\n����1�R��=�X�Q�6�oݽ
� �o���	�� �ȱuʍ�'�+�b�C��\2o����f?��!z�OD��
yo�0^)�Vt/�B,�o�^�<ʲ��%]���� ���DQS3Z��ץ�����b���T��r���M_�b���[��H����Y�g���^;���ۚ�GϘ<塱sw@}��_@�*�9�_6f��%��|���m�ܬE87�ZsZ��[>Z��^�6"���*I�5U�#ز�w�[��H¹M�)�ky=A`z	zz�ޜ�p(,.�	�Vuњ���&�ޛ�����t���z<�C��\He�\E3��A����w���輩V6��Y��Y��;I��HT�?e�	��YX��m��\>��z�*�0�h@�t��s��L4U+�	�s1�� �%b��:'q�0RB������Ȃ�U6�#��dF^�L���|};�fbB��B4�ۋE\�jp�6
]L�[��	�p�P�jc��o3��8H��F~�����	T��XQ�V������Ol�^۝�,�:�����i���.�(,{-F�z�C׷�W�2��a'�YC�1�u��B������W=���$��>) q�mP��:�CV���i�Y2=��exYL��L "�E��Jn��ȴ*������:�`�̡&8��\�����Z~H��1Ӂ�<a��-B����U���x��J���\����{ò�e;�~3|RJ�qB��e�Oݔ�H�EjƓ�������2wɑ�~�[d~��K������x��}N��c�I���@�'3���߯�7��`�_{�1J=�P�t%O��b:��6�~fI����i	�1o"���dX7���;�]�[|�`��`w��{���XC�̬ ����W�0I����:H��d���.�:!��7�9�p��L9��9T��soз���G�9*���{�ΩƮc�oI��˱&Vj��v	˵P� wz�F��ֻˁ9$�qBp
�%�I~�w�6����V�E��[�P�CwX�}Ȯ�m���[Vn��y;����a@��
�_l9��1�Ҥ�"U0}^�]]�V	yc���m�jZ>�?�x����1sτ�h�L�?ջ�:p~�9Q���/SA���IK�H��B�u��\ar1i��S�W�%� ���� I���P5:�ִ5��ץv1ڙ��}�1'K��)y��Ieֲrp����������?��f�T����{@�ޢ���>8�%���7��l�%~�w�W��=A ����Pb�_<���ZC�"Mc�nB~�����d��� ���e1���,��!^��&��Wʊ���aRl�B�zC�L7*b�s�⎼��g6ѽc�1��
������pgkx(M���D1.��f�f�7�.����+ec(-ʚ�z���lq��8�{�����s�߿�Ȥ��V�!���kqj��MA����Z�7������5%¤F6P 
2yŶOǕ)����tm�k�EB�+?�v]�<��h�՘v��PvX���؜�<�(��v��3�KB-�1��]&���56	.�'�\�*�G��m������fZD0��TO�ž�I��Kv�}2]ͪ䔾��@~�Ê�Ԭי:�*�Ŭ������ƾ�<b����� К'Z̉�I¿�IKP��_x )ax+%�-�#���b�O���� �ļ������T��`����U�z9}1�t���Pt	��&��p�P-��V�P�4`c�������m�]a�-{�g�G���ՠ��X��xkw��cط����Sr{��v������S�_\��F��:n��I$�<�HBI"ό@�0ּ�����篦�9�U��t��\�@�s4-yi*I;.�a#��Z$��K���0 ��(=deR4��F�Ak�:=F~��6��M��p5Y�e4;���p����ݱ�>&'V+5=���D!��D�.4>�q/*<�J��T;�� ?&y��:������u2��XpЖ5��G���;Y��w ]���$�y�_���wߍ�ÜM�Z��Ù_�4#qc���"� P��hlcWQ�-���UQ�x��
���d�0��0l�<5��#���CU߃��Ō�	��͉z�j�~:8��@�r_<����+�x�W�:4�I�*�¤Ee�=h^](�қ������f�J[���w���/��X�;9Xt����1rB�:��'J���Ɠ��Ehp.��XPC��L'%���ĸ9�������Z|-���`23Ob8=,��G�=*�}����:�ˢf�Hl�N�kJ���:z�f�L�ۦꨵ���i\��Ȗ%+D�=Y����p?1�� �2nn�b?S�Y)is���l$�Xu�o<?a	�4�c����2�*��]/��^�6��V9�����tF^�F�	�U����� h��I����Q���S�m�0E��Հ����C�}��rR@�(DJ�����lOj�l������|�s����R��Ã�ճqN��h$2���)�8�߮��r�B������F�3Z��a�w��z��>d�%�<�A%a���g�|	��؁����+�)�
pZ |�sr�	�0�_��'�kg%�5u|w��uc���vHG��@�b7Ke�O���J�_�3|�<�bW�
��ܳ�U��[S@#�jZ�>��u⫯�\�4����,��y�f�S��v����;|�gT�Sv:lc�XU������^a���V��P�ֈ�tC\�ѐU�n{��#@S8�G|�X��]c'q����V��>|��P����p0�[u������iD �FYT*��瘲1������={��*����JAl��!D�(��7F�I6|�?���Ҝ�[�Bآ����{��܏�2o��&��*5� a�6�U~A�	�_��-+�mxM!��+X����4"m֔��)͍̃\%>U��3t'��6���@\��+|�mU��4y��I-hl�v��~ؔ�	�@�*�w�uC3�����ܫ�4��N��cn�M�j�|
��MeQ-����٢W�T4|� �7��9G����Q���ʘ���H�o���A��`%�@9a*iX�������|,|i��ݍ�E�,W����\�v�e�j",�M����L `Q���8gҀ��J.���$���{b�&쒱��K��Ae�y�fd��xue�lc��<V�4�Y�N���0~�C������g�Xؐ�S���w�
���@?��R�	���}F�d���?�+qZ�v�3YG�~.d���P�bpdt��}�O��<��b1��L����o�=ѡV2o�c�����P���ϴ��<�»���� X�4_K�bb���g��폫�te��� ������ǅ�6>��Jw�=���_wkskw2P�J:4[�0�.YӅz�HM!����_�������ؤ|�7HP��I��+�XP�RkHk)�3v&�H���"��*
H�!�]�գ�NO0���ʬ�4	㱹wg�#Jv�=�Qm�5�����a��v�\�0
�r����6ǵ4}���ϥ��jٳ�xρ7G��'���m�h_;96=I�B��]er�:�*��K����$�D��,��(�|=GqSg���6&�9�a�ƴ\@^���F��ُ��k��ʾ������|_p��EoQgE��LI�wu�"������l|0T��g:�>�e���/7�uv�7/�\ �f�<u7����q��^�ڠ��7h��H������q�)�>E��t�BQ�Өf�Bu^=ŃG`7� ���&@.κ��z3z�a$��̲��E���!���]�j6:?�&ƨazl'5!�7]?H�Q��.)��#VzW��AeW3݉�N����8q�ul��~�{Ξ�6}���AE���'�b����B�x0Xˌ�l�J�k�NZ��lucӹ����q�[�CL�~`ԏ&/�)�|�X�&i�.o�O�s�EP��~��o[�iƢ��'�%*�~c��� ���|A�yЇ�,+��Fo�*jT r�:�F�fέ���[z��9�Y6��ai&����K�7̠������Z.��X�q�!�7��L=��9�Hk�q�N`y��бN�k��J�ǡ�E�`W��O��� �@�*�ۻEg�F�'5���6�sa�L�g�]�����V�wf��G>/Y� �<~����6��?�>j�{��G������T�s�%i�e]�.�/\�I4���f��T:'|����7r����RG֮���=I�Ӯvj&|(�e�6� �r
$IZ��7���@/[��`XtƮ�x����4RP�s�p��(�.�_��:ʱ�H�gE}�K �R/qrg:m��+��&EVb>�b[m����7���e	aǃ�$�ѱ��i����S=�{�WqMg`"��C�4������Ik2�X���� ��}?���U���zz�/؝��f�$ҿI���4��.������`o����^_�@��"�5TAp}��"D[[b�xq�1�AI�"�2��x01-eB}��kG�V���/7 ?b4_�y�ힷ�VZp��u������}�����i?[�|�-���W���:*s)�Y�-��G�s��u���2O�A�l�t<�V�ֽ8L_��8�;�$f���7�S�v� O��7�ì��I��+�)�~�:����Ē;5"��5 iɋƦC����R
�:�݀�AN����e<۩�uBV�
˃�RLe'�;�Ob 1�_�����_΄ᝃ"r�"��|�o�p^|���X[q�����r{���%+7�ݮO�� \��#$6��i0�ϵ/6g����i~������1/���f6�v7	�시�-�`�J	�}ө�q^�{���V�u��`��_��4Lc]�t2�s��3����WPFS/�#��_�`n�~�2�z�����'�eG�89�|a/������i;\��s(��c#�j�[��g�&~�47��d����'�S,B�"��
�������f���Ý��!M圌hҍ w5p�S�!Ec-��zYl����{��6r����V��7�"M�\쬰���ޢ��-�؝k�s�{�����w7UxTc_OE���_>��Qz�8��ɒ��MO3�z�qhf|="إ��������e�k�~i�oJ�|���#�N�r�3m�9��˛P���ѽ��U��(�q��M�����0� v=�˿|*HGH)���[/�U�A�&C��t��}i���5�$|�{_�aF�=��_SkHx�jz�Qd�+�D�E�T0��
R���4�k��Y	�B�h�s�u�j0Ɋ��W�b���C��9,�����4��������EF	9��-��^)��ˑ{aG�"����k�"7���:�R���p9������4�+6C����P���sxhX�gs->��sAnMX_�W����dO�^d��k�=v�J�@~�o������nW���ͽ ^hIe�����Vl�� !lIj��2������f]z����o��]ݝxDy���[G�`�}��W�p `Z�l�均o����q�����:/nz��,]i�DkX8^�'�2n�g�y�	�����J{sh��aS7 �K��D�?���U1Co���T�5�g�\��.VK�~xfE,5�k�5�j|uz�3V�d��N�=���y�F��Cn��-�3N�g�҂���t������J��(H��jQ��H-[�k���\+�.8����?mP$.�R�\/�SW����!�)S:$F���^���C��#��	-:T���)'K�ד)2�=�:���j�b~6��̈����)��o�i!@d/�s�ڬ̸�o��w�K�
=���iy�[@E����0'@�*tC��q/�a;��)����"��a�B����d�ￆl�S���T���6��rB�u��5��h��#�I�"+"_�^�����w|8�_��*$v`{��;�`<��+�@7s|�k�~$-/Y��O�R-˪�O!���,�ӽI�#lw�5Kc�3�f䩩��#M��WYB��](:ti�mRNĥG?[sxH�QpS�4�y�K[�`=^~Ji�.8G�xB�g�� ?Lh�zE&@�<��#F�c����r�F@��\>��CړA-�#ԭeH�Q{�X��]6�b�ׅ!���;r�~s�m�|�)����H��M꯼����It\���L�kU�-D���kg�ݷg�pv��q�1�_4e5��-�<�*B���g)�/�M���EV�+�������N7�:�!0�M!8��p��R� �s�a�QKl���w郭�3���K���.a�y8��oo�Fk-"А�)U7)�O$�:�ʠֵ�zi�./��W]����z?t�!�(�$F���z�l�#���'=n�����h�d�Xԛts-�M���_F="&'N�ҧ����e9��<�#�ps�q�]u�kI�����0���T?�6F���bҋ�dt(�mz�ŵ7 ���;�Z�A���x�z���̆<2k41ؖ����6��tN�{�
z  �.���8����vmo
���u��}���t}�p%\��9e:B�m���)���A�(��e��Ҋ=�TR,@1�bx��S��*��6����i���O��d/��đ�?�K&['��:��ϩ	+Z�*���$.YVJ���9�ב��B��8a��ꖼ�w�&c #�8��$M��'�$�7���}=Ӧ��f<,e���e�(��}�-��-�J�
a�m��ӈ!E�ӹ�J����"p��� `<w���ݐ��Ҿmh�ڄ�^���0"B��\V�cR[�k^�������&Ƿ��(�s.B;-��-��4�C��`6p���q|�����;H�>K�j��&.u[A� ��ӛ�Z
�֒2 AX��)${���̛��(H(1 ��X"%�m!#5�cW�n8vB����NA7�n�T�f,	̄N��9���]3���d뜒A��)��R�k�*�|@����)o[��$���5��}��Ԛ��'rI�'[<�
����Cz!wײ��S��b�"x7�-�2^j(,��.���ʷ-p�#�X�V���\�$�u�ߏ�����i�Q*���iϨ��|.���d�y��:V� ��n��؄J�7�'�]GU���-�C"�U�Z0�F~Eic��[(V@͓s�3<����i7¹R�*O��7�|��G��5ÚA1�n�L��R�QY:��F����9�ѫ�zc�Un~��L7�Q�sCB�K�� JÚn
x7	\��#�aa�p4���Fka�ې��e;��~ͱ �
�l90��ɽ�Cr����H��e�7H��P8gبf�³�Ws9�E�!/M0:kJ_�vYA�Ɲ�,�'Ux���mM�"�n�ZKYY1j��k�@�ҽ:b`0-����TT�Q�NW0���5�@���y\F�Q�N�%g5�����qٙ�(���T�ߢq�f߬ڇ���<��V�J�޺�Z��ɖJ��o��3�!F.�s�3xfr��c�6�k0����t�(S�#�S,�Z��)p��`o'���(8%�lf�,j��8���Bf�~|����	H�#����+ F�1_�u��V'Ŭ�jϴhK�݈ĭ��_
��"�ą7�Iٷ�����٬_�A#;e��>d"����H�3G�sz��D�}!�Ǭ׳j�;˾�יz�1��;��bRU�X�<��lR`��P��	�C���~P<,�������D��(Xҁ.HY�'1:J�|������r��Qq~���Տ��fdv^>'�dP�um(��|-�D]��R���"ty�r�f�m&��� Fxw��_uw�+G;;ĝ�i i����FgV?���b������-^��Wԏ7;�5�E��̇,Ԙ�_�z	r��s��Mۂ�_�&b�p?z�du��X#|���M����U?x\��c��>�>���"N�1^_F�r������2��/�����nS�0���Q*�1G�m)����/q+���g΋���68J/b`��&g+͌���׼5���nfSsp��k����@����UD���/�jn������a�O˦J����[^�c���hmK�4���(^a'�5�������ةt�7wkf�м�W���Ka�Zb��1�D	kAM�y��Yn��3Ud��el�M��"��%0��:+cb�4l4 ���5\��f|/O����e&���j�qrYS�5%���Ȅb�Ɇi+{�4šQI�R��Yp�
f6.L"��I�4eD�I����R�S�~*2�3S,��	��R��g��=��Z����=�r����ʰhD7�ߐ��W�H��/�_#s]�(��e����6F^�rM�HǺo�Z�V��m˃��>��jg<��i�C���	�u��Ƿ!X�੄$�fXɱ����!
.3rV=[P�ĩ��Dk�W�5D�܀]�g�#Zh��70��i\7�0���Ic�~'���؞ ���P�Ld��A=��(xp;��0��#�*a&�HT�dI�#������%����v�<?��!��^D���zHUg����㶴�e�F5��`�Z��P^<�Qpq���G�;w�M��䗆���Y�l;ȇ�)dVh j�S�����3�0��k�g���3ix���s1�C�o}���rl�얎=?8>~Jt�q1�:q����,�UB"5���{ЅY����s�����W����dM��Ü�dM�W3pI���M*Í��&e�� �} ���{��I�}Z�ϊnd~e��� ��k�Y8��
�;�"Ua��k9��Ma���2�S�G�) ��M�ی���� #{���ÞG�hS���h'�VX5���+m�osF����pʟ��xmt�ϛ�y�,ݭf����/���:u�p,��L���,���l-yi���^=���G�ʲ4�r�d��,5}襐��&�Ʒ�����06�L���νÓ.��e:�ln*�\�X�j����LB��ȾyC�As��Bmr<��{��5�pm�!8l ߛ�8�>���.��S�(��Y�?�a�~���������1����7k��\(���qrr�ѫ�h	l��g�td�_����B$a�Py�U��O,��Q�8-�?&��hs����������W�)�
�\�Mk6(�V�Q��^�ˆ=�42.��-�9If�#��aql��ͧ+g�si@�DHi:օ�%�����
$q�����*6�A��p�:aJ�&~�Q�Sz�g��'H�xG��c}���S���F�:��:��|�y,��Ӛ�3wQaᶝ��	�9C��jF�s��	��Nq=`sg������g�jN�"L\j�?,!E1�d���%�_EC �,@��]��>r��%'�Y��E���P�#�_��h�	dK��d�	��N� ^=vcʣD| k�v�"���H��1�K^#����!2c��h#���ᚗO�ה��ڨ,�Y��$���k%l��80�Ť���������PD���Z�M�Jh��q~���wn��+���v�Z�J�"�4��P�+�4�����j@����<��6e�p㤩#>>%v�֕BE��YL��,��G�׷ю���ء����dv.��eU�=_�J�)�����d� �p���"�i�>�������	�=���-�1�Oܵ��DR)D���ɷ�!�$ї=����>����(�H������e,���vuYn��kX�Ma�Dv�ݴڹ�����d�xS4�gd��}f>Rm��];1xq�Qm��X�ETt[:lo�,TóEs-&��$�L2��g���-������L�<X�D�,�Z9���L���YQx�X���$����\���֖b�>�L5�e���֠V���eې�D�p�H��Vށ�Y
q��+��l�~ܕ���t�X1<oP��?�v"�Ԣ�Ub� �LM�Gm_R��-xoP�H^ ��������ѷ�P��m�ó-���e��C	�Z?V��ȤG�K������N�{j�M�γP띤�1F �햾�oPY{K��8���?�W�-����4�F[�fnr����TzJ�w9΂�:����j��K".Z4��BZ�0P�^�J��I�{ap��̃�D�ػ��w��J�.V����$��fyWy����S����O��c�`��t��z:R�ZC������ ��6�Ƨ���A�_��}�E?!'v�4�=������R�P��	�y�����(O)�fc�萠j'����w0�U�������T'�F=2�׿z��BY�?ه�d���PRx@\[E���/�(�k��7)ľ�+6�`�*����F�~��!h�����0ac�c�� "��҉iW�^U�پBK�]��>��.R~$��Jd)�K�����w�h �$ ��}�l����g�U��
�����r��DI�KK�
�����)ܔW��Q�
fbb��#��\8�`ּ*�N��ǖ�Nk~"F�JV�SȰ�F�e�4Fi>y�|T�@�u��{�<�i���������B~�B'M��2�T�|��0�Q����}��>;��� �-��nuRmn�(��$��� j����0'(�ņvh.c-
�� >�����: 3-09��6� �:���5	�՘`�jo��b�=��P���z���+�+����_�h>�"ΦP=�x��r��dώ�w�E�'O�������⹻g����z�Ni�R�c�J������k �/*���A��Q�f�D~����
�&�K�R�o�j���� #<^�A�߽f�,�κr;��W���h���-�c�`(d��*#�l�M(�*C���V�v(|�B��Q��3d4N�V�䯁7��Q��W�b	��CYbvP��O���~�kԫ�����O�V�Z�PdH�X'3���a�F	�Ip�<\|�v�fd���K�ܪ|1��u��nd~���>����)���Zm��l��ؕ�W6������d��j헍9�H�����L\C%o�F:%bYSQ�V��i?e�X7O#.mʴ}����!s�����ԝ�ì�@��mc��s�ԛ��&I�������݊�I�M�Ȃ�vݬO�~��vY}~���#)��6Xz���+�m�ZXt>�M�E�Tn5��u�Ua�T�\k2̢�7��h������y
��CiP_�P:Z�d�0��{��Ƣ&�2 'Y����e";s&G �tIi�摶5zA�[探L/�u��jjr���(W�*��SiX%��n�:�V���/9²>�v��ܕ�<��H��큛e�k����!J~�����������S�LU�i��e{Vٱ��#�'��ɉN
�:����}-3֒ �\s��W/�l�؞W��T
����\�s�Gui��֖o���Mi�#�uD�������|AD�� ��P�)�j8�i7ц@_�\�F�X�i�oW<7܊���hq�` �;n���;fCƞ^޺ʇ�w�����)�VE����
�'0f�7�̹oR��رc�28����F}g���D��Ɨ��G���
2$�2�T�ȣ_X4���6����"���t!P9vq����Xg��b7�����E��p��N�mt��;����v���Į�ڽt��G�nMV��F�de�D(Q�,| w]C�4��Xq�K�T��SB��3 Lt��
0��O[ȉ�5Ryt;���N�Kij6�wJ����N�qa��Ga Qa)5�9Q
7��������4k�Ԍ��:+剬}���'8�gXMۢ����+��v�ڛ_�x�R5�3�:F>-t����c�ڤ^Կ)t5	T|O����I�a'-�� ��uuXrU*�/��Ii�������)�$n�.�s��t�wA��ʤ�պ�m������Ͼt��PH��G���y&4Q�� �i3�fa2��y����� �g	<�@��=���o�����2��^��~���8V�_� [b��!�:�9��_����
��(L,�ݬk�"6�gzbu��k:����ݺ����o�}��SOR9۳r6�-���( `M%U��8�DM��p��3`���	�R���Q+�Nl��u����Bł0͍�[�"U���S�
�FD�"GH+��Fg�!��	�g�fe�PşL_��-z�Ғ���ţQh������?��˲@L�&��V��-��}�>a:���wV�з^��:�إ� $U�4m�^Y�~᠋�v�!�d���!�����H���Kk�pg1�Mw��r�݌�(�.�i�,�NQ[ �����H<p�a�)B'T��=z ����B=[�w��H+���%rj���S����BEz��{�y��5|�PB�����k�Z5�X`=Ċ�s��nmfM7�Z�a�OL,�r�bD/�P�U�J�W��)�Q�yR�G9����%x��-˞���٦+��>
�a6�cݳ��ڈXmP���@�iW�t�oN��1�|~��ɇ��e��.O��j�~�v�Woi���Y�Z-V��m�g�s�3tA�je�r� Q6�ө%*=t�PLv��ht�I*�q@v���[MC��q�v#�x�m�b+<1K-F��$r��̚�	�:X0#�4>��ގt�a8ru^fS{G�fiЭk�Z���"ƴ��%�#Ro�h}q�8>�b�H��	 �5�E�k�����{1tx� "���^�U�p��%���ǜ��lyl��v��Ӳ;���ɤO�� ��.)���Q��_��R��)}O��;zy(x����o9�kB����5֢:}	B�❶*��#����k�E��,���[�b��P�]G���C��<�1Q�O��`QFԛ���]�눐zϦ�ᕻ�8��f�o:��h9�ӯv�.#�4ٔ��Rv>�4	7�_����c@n$ۣؠ�6O�j��#�ח&P�o6fP�"���2�a�����jYWz�)|=Ϫ��H���Zo�/b��B�8=�{�a�8W�-�a�!�T��Q*�[R��n�Vu6$b3���=�?���N���?��K?�U=Z�X����ُ֡�#�i�p��@�ؓr6YE#�Imj��������tw|��E�4h��p�jR��uy��Y:���l�����c
�nu����5C]C3Q,&i�p�������:�g>�Q����r �`{UJ�w�;$�0x�G]b�9�ȣJ֙Mzm��.E��,�>0ҟ��2焳&롿>vTH��tZ8?Kya�Bwk2����u�*�hTd�H�X��������=)N��?w����p-F19����p��}m����W���eЗ�[��4�W�W�'�6�HiazLU�c�7NЕT	o�[&0E��ff��0��#�mM�k��C� �����j���%������uw�M�?��C��jfL�&�\�IZR�F��%�끲\���re�u�v��+�'�:Vb8?C���Ry�ɛ���x8�2���(u畡!k�
Q�SK����aUm�K�Cf!߳���3S�����,]���	KL~�U㨀�i��'�XҮ�E�?�*Q���=�W� |(�c��t'���;���Ǌ���\�&s�]?�m��y���~%&%Y��k4�J7�K ^��<�C��+>Ǎ�8����Vd[L���ů���U��!�VUL@���b�̮��^��朎`��!�lA�AC��5C,�^���f��%�a�$�#�i�H��T�����t����D�+�_\銿(�R�����c{���g���nƹ���'�2`x�T\Pߵ��6�tC`���ԇ�6g�܈Wd�q%v��Y����^@��>5"�zL�O��`�7F��K�Y�ڭt��Zap�͕��c�.0�}�,Lޣ�޼XA���#��� �~�佐�j��\��D�cb��!���KCs)]PϨm�@&��p��
2��iӊ�JЛ�*(j�DBe������E�-x�j'���S��WL�}A��6L���,mR>O��OdEnh�/[����:���>��u_U�\��s�w��-|����k�	�L鄯����Q�����C.o��E��}V2Q�Gu�O���Z���ߏk�JͽsZdI>3O9:����bƜ:���Ќ�0lğ>P�Ê��]I�CӪ�TZ���2�$�X\Rl�y�^�&b,u�`۔�>ÖP�H�$�Z����Qɚa,+��M���qk�*�g׭�c�?{�gjD��$��ͅ:���d�+��utJLexª�v<��1�Ϝ�Y�7��P|>��r�M$_��������lqY:b�t�Np���d�_�������4ϼ_��)�Lќ@|��ZK�Pw��i��Z�o.�ww�Z*��L�����M�_T-	C�y��G��K\Z�Ӽ�o.jln
����ԩ���0x� �g�6�8�gV�*�Eߑ>k9cC=��X��������r����2�Q�J�3P �g�}�Q*l����<���^�gUUR���n� m����E��T��H16�����5}0!Bx~�Sm[/�k$F�e��e��^H��^哧� ݨ��Z
�tԽ�D�����FA�Kw��j
�I�f�?]�$r�F���g�?3Ӵs��c�p8�Ĉ6I	gH�V�e;Y�U���zw�*eT8�)���Z��.Ѝ��ċ�	�-�=^i��Cn����pI����^%����O��}M_���n�q��ǰ2��T����d�,�\?%�io���R�������.��)�5�yؚҁ~��T���F�|`Do��S�0Rv�`O�;Moՙ�el�>�v`�G�sj ÌC¹�Q��8�Q\�&��K��\�v\�����K_��q�U
".Xx�O%C�Qu��hġ��6M�a��X|��+�H�k҉tdkN��*�#/��ԋB�x(h�g�E>���}{ὁ��gN)���?�!�K�����`*�̃6�gh��̓�2[Rr��Blzb}�f�N[�0�ٟZ2�mWeRG����nX���nq�W���������
��]4,�S�M�A._���\���Yp��^����Uhh}���y)἖Zs��>G�09�߭����xH5 %���Ew~�Gg�O!�w�)�JG=nb�Tp�W�h
sG���Ҳ�	gW�D�S��K��.�����"k@�B�Bj{�S.�û�a\��&�@jm��B�O����k��3�޸���yߙmP1���i��Z��f���ؚ��4��ߐ`�٩G��X���]*��}i��J����y��lR @���RkeOD��&E>�z�শickL��9���WC?|שs��H.O����^W���*1'1 ��ʪ�Rr�*[5�Wh_I�i���ڰZ�6?2 Cn��v��V�O�$��W�0��*bb�_UO�M&�/J���|����&����A�>W;�4�)ʯ)��d��R����%�Q�p�{)kK�z�$���Y,�1$!���+00�&��cx������xXj�R���ʠ�'��Zݨ��܃[Rx~�:���u���ת �7xP�����S�lR8��No��P�j�a��.�fU�����+��pߌ1��?8���!.�-p����mLx
��r�W�1�'~�F�a�M�.�0ք�@	�X�+}q-�i�Ⱦ�tU=��v@?�Bv�;39&.�@R= �Sтǵ�����{�X),��H�����l���vx�O��Z fwP���y���xi�����Qճ����(��0_?�v�����5��^�%���:@�h�P�2a����V�׌Z ���[��Ua5�l�i=����n�*E\� E 6$a�麖����.;�:_ԙ��C����4D=�ӄ���Я)�=�V��w�X���W�~��d�o']�+����-�[0�DηBD����׏�R�ϷJ8�2���f)�#�n!k05��2W�xq�c���`y='��k�>����5z�c�$kT}I��J@g��7dOo�P�Eu`	ġqp�S����ٮ��c>��A��`�H��<���cuV��L�xB'm 2�B4��@F��^�3��%����]��7A'a4>����&�L��8:4>V��!z���%

k�� *�����%IE�� fL�t��5|���܊E>\z[k��7�֧Ԗh�0�.�M<���#t�,'�w���i��M�������w��7}�B� i�H���Rݢ�_ ���ޗ/�5�G	lJP�Q����h��T
H�.�uK�T<l�w[�yO�W�L�su0;Q
�9��V��7���^�=��ߚ�~�b MA�6�v�>�ф9�c�V��<��?����;��vzp����ZI��2�j^���;�gR�_� �rAf�5�0Ι�L�qR��9i�F[�:�I�~��ګ}ݧ̇1�&I�G5�r���V�;i��ywa�J@�1�l!O�e���cv��:�K�'��~��6��0�ݫ���f�@�2�ޚ?�O:h�\���M��u��8~.�o	&�(Bin:s�M�ރ�O�QHdt-b�D�Y+],gu�k4�u��ǋ�贄g�+v�{EB�;C��e]����)e7��ſs�U��i��-%
C۶�3`S1��nr{o�wi
Ŷ�/{B;%O�@��^��l�+t�0k޲x���Y�x��4�D�>���ֻ9��40$Ǥ�f�2ً�����6�H�nui������YU�rC�8�8c2z�&z���H0AAm��f~DG�ق��\x��+�9����P�^��� .�+B� 5���mi�����V�Fg��[��k���|��W컱@Tc�%VwD���vg3�΂�,tQ��(Ip,͐�d`���N�.��b�@!Q����W����_Fɿ�U��g: ���S �CO�I�E�?�����x�[��F��	:�oU��k��:�;^2Et��ŘǼ_X~���q�ʝ�#����հ=_�ؐ��=R�w�_i;ɕL �=	4BN�
��Y\��M2��
#T0
����!ךiH��_7���ȶ��_��X���0\GOl�,R�S�G2���>$Y'$7w�x�r�qk�i�������+��1s��KpW�N�U�U�F��<�K*��!�M�UT3v�l?��E>�.�:$��s`nd��t
L�4��&����*N��!��d����$V�"' �`�ڔ���o?��<TM�&2�$K��$1���x�eEԜ׾1);�Y�c�:�ZC��5�FӆA�)>aץ�ʒ�a	��$|�װv�G\z�>U����>FPT��f��J�2��A����/#�7���; SO>�3����AM��(3�Q�/��"��f�wY��'�DW�,%��ڸS熅����F���{���6��ƗdTi��37r6����&�&˩Yr��c��/L���k5�W-�ᆟ.��u��x6�Z�,�ޭ��o:��JlF1U����*��X�,�>����E����Ƥ�k�L�Y�k�A�K|��_��xg��2Q�-:��"�.L��ZX���}|*���H����e�e���i�}����oې�'Ճ�pRq��]A�ղu���	*f�k1�c��ra���%���6�_��)���~���2 M���r_3�'8�؀� ���=���jK9,�\��0a�/<
�B"ҴQQv��i;��9��C�0$� >�����>�6RfZ�6f6�����B��M���D��SJBƔ����PFR�B�i����6��m��6u���~)�	v0YU
���WB;���|}^�qŽ�<X��D;2dV�}����~8�63=d><�.#�"1�KCߠ�ip���-U��-ǻ�?�}��D��nM[�QB�5� (��V�|p������%�Iy�����:(�'1>����jc��2��3��;�~ҳ\��3E���J��2(:>Ň�����7�#�
�X�e���R~x�ZX�چ�;��o��N=U�R9���$�ˆ�"~!��쨗���Ԃ��![�a�:�"0��y�mi6��ߘ/w�K��	y���=O��F�z�{˂-�x�d���<NZw;�D'���Tֻ0��"6�c��
�P�@/�.]�17�6K�dZ[�|��I, ���$�� ^(�����M�o�h�k-��%�g�
ʟ(M
�H����^njb#H%ҷݎƜ�טw=/7M�d��Pk�n!���x+Z6�)��Y_�Y����ݽ|X����q�tx+F4���SF�>��&����V�2�`xA�T�x���k�k=�����jC$V#:'�+7*^�=���3
*����p�~���$�z�VG��6���mX���E�����P�HV��f��{���S6Xr�h�#�>*�T�ئ�z�o�x�JQ�Zؚ]|\B����T����f">�tM��,�`i^5��2���^M2��6"�h���[�t�tƔ��ҟj�uF�{��j�ذ5xf듡����'�r":x��
�+_����U���w�ֻ����^�\9m��]�YN'x����_E�±��zG[���~~���U�����?�Ba?��ЕW	�c����6�;ڇ�e�,��	�O�(�c�)J�=f�qp��ݺ%j��U�j�8��НW����5H������	 �����l��J13�q�j�(67��XJ�M����y0�A�f�ػ�5��a��W�Rz����91H9�z�Dbu�\0���')�ݱ *�c��_|F]U���U'y��81������`���_��p��*n�4~3�.�P���@L{��Z�6q���KO�H+��:���Th��	���`J�{bR���YS��9[�������%�k���R���[�J�9O�te�,)s=�(NcJ��\RE��9��ƨ�N3eF�?u��ޑ�d/�0]H�7Hh�(�o��0J��"hh�"�@��`����xm:�V��~SoYs�3��fΈMAvU�S"Yy$EF���4v*N>!Ǣ�8!�dr�~â�^=WNp[���K���Ql�	������!3�
DM. ��<�Dș����ms�$��F��2�÷�i��];Q��\��c(����um��y�i�RZ��k�4�^�=�j4���X��P��t��`�=cjD���LO*-�I�E����RF��Cf(�^��R/�%�h��W���|b�e�ƶ�;�;�L����D+���7���8Y�_N��?N쿿����V�2��n�G9i���b��@�qZ�H�<%{�{��џ%D����c.�����c㫜ϣ@�m?	d��~��R�iyd�ԲMf�F��������#!p_�u�(�Z6�h��w��)b����?í�'����٤�t�����������D���*�\.Tg�9���w ��đVZ}R3Х��J������X9M��*ʠ�`R½�F���+���r����w�|�0ڸU�ZSXa'Z��e�ZM�>��a>�V�{�78{��}Y f�����B�y�7d���f8}��⩡���f�;���	{�Y�.�&�P��w�XwNY�Ne7��f��d�Pu9C]����b���D�r�˘�ԟ�P�Iс�� ��Gz�id�ьB���/Xg��*)(��m%*�fި�ु�z�K�eh��{���{ �z���Փ�P_=] 0�6&�]ܢ�>Fbݞ��Ы*�&�$�'�ӎ�[9�³I�q��2R�略�,<H��M�o�#S�6Dɶ���u{�_r��9t~Z�q�=h�ZTd&������MC'����L�d���kWH��Ui\Vܕ��M�I�J�n�)�7�m6�-�C�l�)H��/
�����o�"I����[\�x���dZ�Sz#�M0�t�RQ<!ω���$z{��`[�Z��"��S#�UQ-�uw?�'o�Cn��[��P-�}�߄A�2��Z�(\d6	` >Ł��V�g��� ͢v�4���~�GZi;8Q$��9��B7���z��3���DK� �8��:ޯ�-�2�<w}AA�����hB��ٱ����X��ѧ��C(c8b^R���t&C�
�Z�g{��t���}O�&sIoӦ;ZjҝYO��a�%K����E���zGѸ�U�9��o2�+� R̻�(vD�,	nt���_Q/�Nt��8Sޛ:�wu�,}�UU�+��YɊ�����VO)���0�v �ٞKZECR!���hMI����"[�g������'�z�=z������vs	��!�y��G~���z���x�t���hcY��{���=��zF$�?��i=�X��i��h��(O4�#\��z0 γ	��k9ަ���·�Z��qv1�]%H ��Z�G^�
>�j�Ř[�D�y楟X.1d���;���{�D�C0�D�c���Y��MnѺ� ��{ ���s�1��ά�L�ْ��L���~~yDv�,��Z^xӓ׹1��s�2t������B���?Oa�B\y#cݞKd���]ߜ,����r��mI1G�i�S�"C�Vk��l���»g�	�ԕ˧���Ი�z[�}:���Ş���u�E�19��Kk�����?�2}W8o��7�������T/�y���E˘� l'O��,۱�Oq�k���G�~R����+�+?3�o��Ô��=љ��Nȟ�a}��,\7���լ�GJ�q3�"��	j����+l�Sԥ�(f|o}V�^��K[/1ئgR>��.�:��s���|�Y�d=Vz��7��$����(�ak��ԩ�,o�Ax�
�ǚ�u m �I+���s��Wix|����䄿1��H��-CO����֚��·�6�$�`h6t�S�2N�̿���!*��Z�Ujb �q�y���p_���΢6s�|y��o.��m�<�]�N����31����>�+�BS�/�(\�~W׌��l���Ό1�0v��&����i����j���c���CX��u��������n8�)��<+L�]�nl����a�f�8��a�7��y�����3J1n6,:s&Yw��"�$ �;d+J�")�����u�c�"����3�|���z�b�$ʫ.��F�؉Ҝ�H�"��k>���"����ɫ��P������xҽ��V!����Dϑ�f|�4�p#*����N�/�H���9��+"Z��v��xfM&�w{�2F~�I���;�z9�W�����uhhRZ�Ԙ�,}��@DyD���\�2[�����a=�Ѵv����BQϦ�M�%�+L��W{�L$�\��+%�K@ITM�Y�Y���#/��c�W����+�Rk��bt�D7�8޳N�d@���Y�殾X���j�7:=�V����\<������)���6�|�c��|b�Vxa�K3��J�iژխ� �v�4����Z����w�X�3��RB�H��}�:|ĬOc6ۜ_`7����nOA��3�y@�5��� A��M1No��kJ���e@\�T��J�Z=�X�����6vp�}����kc�β��v:d��9�����}��/�q��ӷ�U-G��\����!t}q�Z�ո,��6��>��$�̙x;��ߪ��N{|ͺs�_+f'��57q�O�u6)d� l6X�[R��K}���"t��<�pܧ���Td j�Q���$u�>��o�	Ԑm�u���_˟>[5F�A6Q�I�6'���#�e[���;]�e�`
6sޝ���a�Q�� ����.�dN8ʱq�9*�P��T[8[s����!������ ��]������;~���Lkk��K^!�$)<���S++���E��`�0#K��˭PF���8Go<0���%=4��̂&�RB#ž��j����%9���&f�z���s�oe��<U
��Sz��:A�2}3b(��4�-�2FU!�}G4*$p%�����Xr[����F���p[ϭ)=�8,����윬3q�i&��%����K��Dsnn&w޽xQ9ޖx;�h���OT[���R}`�D�!���蒍�x�>��F'g}�>���8��?~���mT��߿n�2n
���V�O�I�?�/Iw [��:��$ʝ��=����!���K͇ÌI����I?6>��25>Ej7�����p�w���Y�w�ZX	n�h�g�`h��'�m�Z[7�ۥ��k֦��4L?(<�_����~�kP"fk�����h䷹��.����ߓLQϑO�������`�.�2��|*��&\�Y��z�x$�Fv�!>Ғ}�����=n}��	�Lo�y���*�$�ȒI����9�8���?��N��e21�Gy3�Oa��≀SqJ�RVk��v�*kS�-��0l��o�$�<�������s�0&���y��������$�{��/�և,�O�I��+e�87��"B�TGO	��4������-�4oy
u��3%S���6���C�hy�ݒ^V�ؓ_���6�`G�&����.�-6g��fِzۗ��.�;]V���D��Ŷ�'%����]�x������~G�RM�,f��P������d�*�ܗ��>B:X_<r���\/�e���y�H�٪����hgr.w ���a#[d��"H�+�O�:�����ho8<[ö����lf��s%ꥉ���J�������}2�EN� C(O7�Ln�=Sl�T�D����>���ג��!�A�~���|]B�L���TEBz��hf؛�=�����6}���\�T6���R<���j�ͧ�c	`L�-���Md����r�cU�!KM@Ƌ�{1�&�/�ؼ�ʀZ�V_��Q�G�Ǡ #a���D�� �zp�zvG���-.���;�����Z��k�l����^3C��C>�_��8�u�j���^�� ~��V�� �	7>9��Z�v���BKŲ��,/Rمg�O��k��w1��9G��M���ǣ��b#tu� �9GB�PV$�i��'&Wʶ2��Ye����٦������Mh�U����}��DPO7(�~�h]�kd1���cqd�*�ۆi\������2�����ws[5���"�:�r�q]�[�*���6�� ܄ ��Q�.P��XI���&,�������z.~:���}޻�^���|��2�i�9!�Z����_B�\.�#v����u���A��%Ox�l�^�2����J�q��?������� �x�,A�+l��Ab�?��q�Y�������1O^["���!��(������-�F߻ǻ���X>X�~)x�c�{e�G݄|�>����l{�|5H@zo'$c!�
H6�%�5?˱��M����.I"�p$�1��K�SP�q��W���$	^1�E8�l1�[���(���d��H�3�˱o���)�@fn��.�Ȏ�vv��3��C!�����lv�Ql��ƻ�" ZL$�L,�ެ�%u�=A	q`=wJ�	Ɯ��' ��5H���ddz>�҄"�>2��cv�W�i,�x3��F�0��k�Va�j��;F��aD̼fȄ|�r|��u.�]�s��{z������O����wb>�m��+�����d�I��4��9:B�]I?>>��1	AA��B�����]	�@7����t4���@Q\Y�B'S�	��u�-r>S�F��j4֖3I$�+69�b���UJ$w�W�3*\�!N�X�hlu:<�|� J�D�+Ѡ5�W�g���j��h�4�W������!:�4]0~�,7�")r�g~�^����&���R��.�L�=�팭�����μ�����e�'x39��= 9x:� ��.
�PI�1�u}���@ZeЉ��!����-D<3$|C:�����xU�٭���k�R�)AaT�/�뮵����/�/'�f�I|,�����<��N�z7��=Mb  C9����e�J���p�SJ�	��	4V�W����`e�e$���Ӹ�7T�HJ��X2>���`�c���ť�2� ��V�ެ��^Y�]�+��1H�;1ޗ����(�q���b�l%"���� ���+S^/�S)�P�r� >
���hcF���1�Դ���Y�>?Ҏ�̭d�_�ס#���_j�Q��rpa��s���Y�n��U\���P��=��J�5���뀣(���=�D�|^��Dն�C	�k3g���G�b�b�\+A�2�\��'\�ڞВ�%#8-G��@+V~zϕ�����Ձ~���[G�y����z�Z��K�'P`�N��Z��й�	�����*��Ɇ:�0l�7u�p'T�
4��{�S�'��Z���C,T���S�r�2�r�<n�](��4e�ڳZ $a#l��Z-a	\)�?{a�*㛗�Xٽ}��pn�.KN3����X�3�:�ec���JA�n`5����;�x�:�9hI���h���Ot�T%*����fsT��`�.�H���C�1l��V��n8v�yD�_fq}F��=�Z^;�=�����X�]���?D���_����3��U�ץ�ָ,bxt���<&r��5����*\EK�a��C
V�:��c�)��������q��qi�
��
=����H;``� C���/�l�>�mcz����������I*�y�"��<$��>2!�gAF�w�uj�\�d,긫���&{�	rk<�8+����K��@!����OlP�;�����}���OX�j6JE����w�@ƞFqG�x����|����ES�Ɋ����`�6���D}�ǳ��M��xz�9]�7d�~�$�'��"�q��c:B��c�y�o�u�q��k�}!�PBR��/�3]5���(0���XU�6bF`�Fg�Pn:���N�P����UHr���#���8�ǅK<�3�۸�uB�H R[e���_9�4����5=�ľK�	�`�F��P� @Ɋ�)4`m�s|�wEc���|kɑ�\C�'D+ @�p��&��ZD�����+�����n�w!���55�X`䴰�R�\<Kf-��VK�3X���[Ɔ�̗g���
��h�
�]��E(��Ui�V\�2:8i�F��J�`�ϣ%�E��S�Q���3q��+Et�U]���;�/ա�_��z�psM%�h��`GL���* 0�Nkc���HS0�܃R�wG�ĝ>Cs!����]�T���m�2��+)B���c�Ny]�<1��"Z���U��6B���/�:P�[B�Նؖ$�K
��:��!��r[���!s)m'$����w��/�i6�${�u��T�#�\��ew��k�rq�~�g�*�m�Sz�5�|�2P��E�wxٸ1�H�#��uO�����x������$�yB,E�{��*r�5�Z��?�Wȡ������������WL|F�h^���c cd�f��1�3^ۧ'��|jY�}�h�e�NsQbI��=���pR��,^��۝�F�%e\�{�l{�PQ��`�,�;���uI�CE�Q�I���Ak)+�'Kj�d���#�	�����H������_0��׭�_�-��I]$���"�bf�_5�w�z�I��%�8?X�oHY\@����,%?��D�d�U"l�8T�y\��<���#�gc�X=�_9�7�[-,m�2Mm�Ïb��0>��o���b�]P���/�(:�kT�����SK�m�04���$�Jz6�"X����X��&���x��b��� Pgɖ�Hr����_�PБ!:w�׻V�H�����m��vfB���`��3������="��T�ШϦ�Pkn+K�Wqo���)(���ྯf��iW��NR����apx��"*��.��2���B}=�J�����,����)K�����=�z1�0pnOUy��01��0� �2��bՈ�
��mY'zl������fӻ�Ƚ!+.ȪYP��v��H��w8Hۀ�e��Tp�9�p�.����E�V�g�O��j
j�X�T�3��x�W��5��) ��!��Z�a�o&�`�������;p�{'���r��͋3s�=��c��r�%Wїx�Y]y�I�p�gW�|g��_��e���!��j9���9�J�͌��=��o�d� �f���I	�%��޵��-�'�-�|	�K�:"������̑}�T��Gt?���2aZ-ci�$���ǃuBQY�m��T�{��|�S�1�T�������e����k� ��V�؋�x�פ��/�U�P[�}����Jr�2�e e溊��_�ĉ���m��e�q��9��V\�y`�1��O)���r@ǆ)b�����N���n�wc��)o��Pd��z'�w��<s	<Z��R��4�@����Πn�B��z�}�sm���cK�`GĒuM�� �qp��AM�6oNߣ���'r�r���h3�OA|��U�ަ$��@@�)�S�y��R��W�i�+�>L�;}���wʊ����m~��I�f2)��9�q	'�t�2��H������v�^���s
^�c�b;����Jݶ�^�oEd�
`����v3���y�ȿ��+9aY��y\[-�	�[��qW��e��z��<��y�d���{�X�
!�:];)��
O)o��w;s@�� p��lѬ�bX������r!h�ā!%z5{�LI�t]	��|nDq�.����͝f%����Vo��XE����uܰ�q#�vR��Y$x���u�Rю������y� A�(I�)�b�/j�����>����0b"�ܔD��AoP��m{ɛأ��$TmBj_q��0^�s�JA�,	�G�4e}Y�q����9�z;-�����U�p�G�o�\� �s{��MφI!����E���i����Oz�.�9+���e�ޭ���4(�.�) �'�Po�9�����{��ל��
�y[��IF,<	4�<�������UM%��r�I����m|:+:�e?�
 {C�nm`c#�0�V�Wo	B�̸�d�aj��1wFؾr���tJ�Ί�J��BU,&:���BIU�YQiH�¹�z@���v�XF׉g�`�Ӏ���Υ��]��"|��J��4���J��-z��W���ܯG�L�@������r]����'�Ҟ� r%V�
�}̇�g�Y����؏g����5��Ga`�f�ɲ���F˨cEn.Ju#�0˭�{a5.�~�e�.P06kk���Z�7ʓ�����>ְ�����E�f�� u +�W':��̕�ͬ�����>���݊��3����u�n>F�|i���\1
�,��W���o��(�ZO�ewsޜ¬����M���k#Hɱ�V(�H��<�+�5��}�;L���)?mD~�����ޛ�.��"��N��a�t��fPVE�N��3�،��J�Y���t���aZ���1�@�g�8�ao�/b�V�5��O2WIs�
O]����f\���8����ҹ�?���.v�\w?+C��z�\�o�w������ݘ�H[u����5�����2��u�%/Y�A
���� gJ�$H��mc�n�͚LV��dM���_�ѽ_�RB~�'�2E��xO0��8���[r�ӽ6Jwu�-���4>��
��*�пC�d��6��<�c�\[�w\c(�{�XS�V�&V�U�Q�&��ٝs�4�EJ�޻�8�H]�_�%s5*v���s��xYa�3����1gzI�"�W�����*q�I�+��-�}Z��L  ������v��,�/;�8�~�']����#�%Qb3e�TG��5v����E^���ec���|/62�C�dI�twE�����< �/���)r�@2���)�*җ<���PE���V��[4�����.���6��O�������4I���	0�0�J|�aZ��@�z��Z���J^Jx�n�:a�(�\ܡ*r�-�+�bee���Y ���19�Y0
�(4m��y�YF(�����[DTm����2U�|�1&1�d�/}Uw�0��\��{�����t��>�q�����R�Qc�, c����*d��s���|%k(���������5����=��b���6j��8g9=Ns���e����r����.#%n앝�Uc����0ʠ��Ǘ)1=��a��55>W�n&!Htܗ��c���f7G��j�˷o!��\��ɚe�V�@�O���<K�����g?���f�9�yhz8�:�>������1�	Cy��%��T��w�wg�O7�ڏ �~�㸥cw��lU}z��"��_�4�n��R�ú�(���{��}�k��Dꆯ��ۚ[x��n`��4 =�n�B���z=�-�ŷ�~�x<�Zؤ��-YA�ݷ�7�ŕ��h�ep�-�
ւ҄�-��,����C�|\�1��emD����ܖvN�R|�W�E�6v}!�h#[�Θ���j���b�iyO��� V�9�-)kZ����0Mn��m�Q$4L�|>7u����Y�/��?n�Fch�Ti]z� �������{]�'�R
a�&�T�@��b����e��џ �.K��<K�� k�X����	ϓ�E�8��/�Q��8 �<kT@e�x�P���ζ�ds�7U^+�h�]�纫;|��'I<����7�(���=��Mwa���pD;8��*��a%���-fKE³ ��8���`�Y�Ҋ�q���� ������ů��7"$mR6��w���Yl �;��DW[��-\���G�p ���
��n�������jD�`�@~��_j���M��
�-Q-�@9� z�R�ipBK�+�sc&�0�������q�T7�ࢵꐄ�7�h;�,��(��[reK���y뙟Qef�3Px����W��U
b���0��Mw@�̬�CG��љZ��O`ol��d�k�8BOhd�<sB�ZaO�_d(]��w��� �
�S�8��>��Om����N� �U��*�׃l�����`��@+�l��2�ZK�-w��0��T��H��)�|Ϟ��|(g|'�% y���6,�m����6W�ڃ�pf�N�g��P�.%���@�@%��\݃�C�S����y�AZ�"o�s�(�q���w ��-y��G�Q��gqn�f*Ku=\-�"֑0����'Ф]2�+��$5wz!���f����W:s'�zE�_�O��XU�!v`��ͫOtJ�w:_E�*�s~��n���hO�ݖ$��� �����^&@���e-n�e2(��`q_IƳ����_|t�?�S81zS�2��7mN��ʭ���E��V̒�l$8����*c\�B��?�*y��*���rZ&��CW"s�����h$��:K�.���3���	���3���%�&�)Yd�F}��݁��Uh����"������2貢E\�V���q���7[ĕ��:�q�Ēv��^:���� �pL079
b��u3j"�`���M��f�<<S�Gu?t��^s�͟h�
.̺ο�<�`�1����U}��"�"3VęF�.�|��޳�#��G�,+5�jqP[`K�Q3O�r��i�)Z�YБN�գ���c|�̂�<�A�U��&.��]{�b��O��p3�7�a������(0a�����:�L�̂7q�C�W��}������`7�m��R Y*��,���wi��Ӂ�K�p�� :X˗Lw�6�q�Zq�TY'
|���E,�x�\����Կ[Z['~`yQ�G��ŗU�o2t�x��.�W�w�����x��ɲX�w��]�ML���|�68�&���JF9J�o	E�L��T�.
N��o_z~��VyP��>�c2�ca
��'��5ȫ���J٥;Բ!L�����G@�X����a��/@�>�S�xzy��c����Q�Z�n���?���,��V>'a�1l�[��[�/�1��±�y����7�m̚Y������A��L�̖c?�Q�ȅRN�"	�(�|}}�9�x�!Mq>o}�l��cVic���:4��d��C�a�U��A��t����
E����D��]���/��A��)k*h�0��_\�HE!�8�Үf�'$sQ��%ت90"C©��YJS؂!ѧ���@�R�{�3��H�M��޳��#d
iͺq��WI��o�5�x.ch�RS�ȭZ^W;�ٷ$̜��}�6�m�}����&���+G&�Z�5H-���Um���Ek����g�;ڵ܉�����ݘT��ӱ#	�����;�S�i%� 9��i�=?���pa:v����-(���wĀ�l��=�_cF$�LN8�B���k;�3��R~3̚���ZK;�Q�>��xp��g�'����/��hV�%b#�io��þ�2=a�İqw?�����bAJo6��X�c�T�xk�3���d{����do�Ю��B$�!��}�#�ɓ,��]��.a�
� �=W����h
�/��<�g$N�ǭVJ6`˥ݺ�ߢ�Q_��F/E��azP��=�Y&[�V�2�8'�E;�5�C�¹��iJq�ء;��/'eRmh�R%�fas�/5��QTn�����L�} ��S5�g�����T����+�4�H�
�pmD��I(@-����n�P��'z�Z��e��t5����`�h/-E|�.J�N�	!�[�Ԕ��y9Ӗ�#�>�I��8ml�x��ay�����E��"�1� �`A}�ì�P65���C��]�bu���{�딾q]*�mQ�u�E][�όqE��GN�d�i���Jn����F�0#m�߶{^g��(ʵ�e@6��M��[��1���CDC��5Ng�z������e�E�k����� ���R�Ysԕh���9$���jd�y�D�r��Q��hd1ѭ��� Չ�t�t^*��Z��E��YxU��B�p�+���8�<?�Y%5��V��ۜ?��[��i�ߜ�<���S�v ����:�HZ|�j��{gLƎ�����
�3�mx���7Hj�~ءq6sX,:Fgor�Vb�ۃ��ٱ��Xf2-j���B%<
~\�|��O�����(#1C�Ȏ�ǹ��֏�.ܑ׃�T��d�`�rK�/`h�A��F���o��Y�q��B��z�柧�2]�<m��������Ul3(��Gs�g,ڴ|*rc�� �U8�6�G3��?����D݇��Ya�7bS�~]���,�p�9[�ĠI����Bt����?�\�!/l!�|��%���	�;�,֝eeg�(=�۴� �鸇���D�!P
����Y ��y(ms^��j���[�81��|���*G+i������9���+�o_�������*im5/w������u��1^��1�#�N���.�V�_v�5�RB�\��(o?�q�� L�3�Ϊ`����Ӆ?m�}�9��f�Wo|��[�*�'��T2��Ԙ���W��j�t䔵w�:n��s�9��� ���!�{ W��#��g�� �{_a;��Y�>�ԛ�!��K��9v�4
�i�B4^��P<�m�1��Q�cNO�4�&�9��\ȸo~)dM�|�����>P�}jH.N�.�:�n+� �^r-�`�>�jm�HO���l		Cxc6�U�n�$�p?7�>���:�X�+T�n6[�~���c�P!1r�ރ��"��#��t��^��~�Iﰚ����?ڑ�RŜ<�7���Eht��*���;�9�ߊ#��뎳"_�(�(��%h70F�ӽ�J p��&õcr��>/KK��E�&Y昹eZ�c�i��F���#~v�Ay�U��KzO���ԄY�:3F����_��kz�������|����<x,�T@���`ЎoT��\���u�9|��3�*>�<�AQi�LTk2���s�V��9��N_":D�Q:������p���[�W�f�0���!༌�R�:[���e)�Ȑ�q;:\&4���V7���O��x�}��!�����w
�A"W��g lGa�̏kܐ6l�������,�S�0QK�_pjr�J��emN���aP�zB�����I�-HI|
,�����򙴙~�-.k�����~�-�T�[3p$��5DKE��_�l5�h��V�N�����m�~gr�˒��
HX��D�>�]#{�d�e�o~�W��ԭZ�&C�8���b}{:�E��>
���
]�B����=C�uv([|�f7����'h��AkY����6�A��s�M�]��۠i�^;��iO���v0�<h�� ���F6�=����Ha�q�ߡ�ޡ��D~����h=�ī~[e�q~P���<�'Un��_�z�w��̋J,���b���յY���Q)M�f�p�ۙM˟�IC�+�38x]��OهK��R���	�LE^�ʰ��2��3z��z�D�R�0jE+��-E�/ X�pv��"��!��ǝ����u;mv�@W֮}����eDA��ӓʼ���(,Lksx��u��E>2N� a����'�;t�-'�-L�'�}��j�G3E����2��G��OWQ{��%�q�zAa�xR��f�=��l/��~9�b�LV'7&[]a��N$��F��j�.�s��h��q�<��n�]`����b|�5�P�q��c�֧#�w�g�I���%$�A����Rb��n���¨���P�%ɪ*4���(znAXÌ�'<�{��k���~/�I%��fn�\�=Mʩ@�������hz]���8��qڤ��ĭ-?�ͭ�3���.�`���<�V��=l��R	_��_s�$;<��;�6b)@�����񊆑�xa4�����|J
���_�#%� �C��^�AM���k7�z:$�E�Z}4������T�� "*�����э�U��M�zf�5D����Ȝ�_��� i	En��#tunmEDK͆��=&�����ܦ�\{�����ö��O��G�Wng��w���Q���XoƆ��\�aiD��}�7��+�D�z׼,��?��JK/�=�����{}��c�_*x=� �	w���B?$9ޟ���=մ�I�?,��6�QN�[�b�����LX���s9�P��&C�^F8u���V\z������8rl]�9�û>,S''�0��?�n*�x����s ��ƛ�{tT�)OU�o���Rl���o@����c�n��
���*�QQ�~-��ꮇ6�F�hQ����=?9���o�5o���8�0g7���]�;���#��Gv+?��Zۛ򌩓f�1���eI;V��y�)�%�i椦�F�,F�ES��J��M�~e��� _�����,8�4��U��eQ$D�vW�a��_ϰv6���LɧƔ����!iC��N+g��&���6������R
�B�>΃Ї8�r����ys1rG%�&<¶�K���$K���@�.�Yg�4��(4h�]���Bʢ��9�D&N1���D�M�'5��8�����9�Ė�����$�Y��{A$���f�䆨!�?��� +{mY�U&	K	�DM'I��!xN! Tw��0`���41Tj��|�V�dr��@?ϩ�5ͥ���l�벟��h�����] �{�Br5�K�5�[S.���Q���딵i&�\�R*�H*�t�U:B�$��Xj���s1Z��b����zz�V��/���W����~e����9Ք�m���X���/�X'S���m\=<�ǰa�CK9��1��=Q���������q��	&��	ʟ"Ɏ����;��z��#s�P�����)v�B����7��Z����kQ˙~>�KgL���EȓL"o���.��<����̂zj�ާS��1O����r���W�$h0k5a�.4���N�� <#JW_��0&�M��ݵ��Q�eB6������-^>����y��y ��^;uiQ���xԱ(Zjޚ�1�,�R1��R �u{Dyd�Q����P������a-�Mj�, cޝZ�)����|�����ɸ����jq�@i��FZ-,|�@�����5�[K�E�F9���v�G����A'���;����;��	Sak�2H`t�v�lˎ4�H�X��@rh�I=^(+gF^A?�͍�1ق=0H���X�E�����N0�=
�fk����H?Fl'���F��u;�4A%t.��\8�*�E���1xR��E'$C���̯�%��<]n;E�y�j�3
(d�g8�a�� ��
�g�f)��Qx�Y
s훊��ZX�q�{�e%S`w���N��PȌ	[^�Bsl�,�/��b �ZK��e���$p �o��:����DO5=s�$Y$Ų�-��X@��V
1R��W�'���7GDy��f�G=��q]'ǽ�b�B1��]#�x��ء.�׺>�h�ҩ0��2m-3����E\	W_N	�Ed��R�R��p¨�AvW��ǧ'׀��tr���@���� o�����Y�S��;_XF��#�`u[xq���(����v�Σ)
�郊'��Y�QY�<��]�)~]��z��'�2jo�T��6�|aY��M��Y�>����&�1T� �bL<Ъ�orP�b�q`�T�����Q�B4�����lY��\8�}�����L��G�8���6(�5�3ǚ��w�!Û ����|��վ}�&������l��]_���2[=�%��E�!&�%��^x�G�8˒�IP�����JL5��)}��A���ov���^F�?�s����j�(A�a�?�TE�}�$��1�ؓ�f}�n� I�~�8O���PV�Q��8��F�Ć9у2w��?a���=ZUge��~~\m�{~���rnsayx��D�'y���@��!��څM�;+1�x�]��SS}v�wqW�p��7ܜa��>�RnpF�|G��� �XN<Ѭ��&V���?:��C��J{2�)f���o���^.���u����Y�Hvi��Ǒ��C��>��Y�I+�v�uS���]�}��H�*�{Z�>Z��x"�ED�q�T�H��X�8�[� :X ��ā���,�wf���]���"/��7��wn����mߎ_����=�y��5e#⼤4��r�F9iyoǂ��*�[SP:/��V�2���`_�Bg���ͼ�H-I��v�_�
�1�tU{��E�Om�^��oҷ�n\���0�KБ@�D�=k�U�_q](�հ�$|�q#��S�O��~~GU���Z��5i�Beݽ �b=n  �$�U'���c�g?�[n���c�R9y�x���~R>pw����
S���4��ǃ���S����}]�|��w�C��,�c�s��c��K��5r����&�Ct�������U	
�YR3��^B�XKU
7QC��E���^�آ�")��ܵ��� ����)��X�-ۺ���H2��#Ҁ1V�'�?�]��8�=��[`��4�[��J?eM	�/юS��r	����TMC���z�-B�0	����"�`�m�k�?i�4�eKPy2���6zn�a��#���0"�T9)�9|<�A�������2�V�굂�?��������2W	��f�t܆�^��l����󭗷N2筷�M�;��}�&=����k��F�$�*ܯ�}�ě��ٶџ��9Z�4LV�9�
�xo^P�����O��b>����)�.�馩Z543��K�YNYs�-���
	|��!��AZ|:G�xy�F �'��K���`���J�aIj'sM�x��}�#���H.xl)TI���3��0��t++�-���~+�g���Y���lW�A�#���X�b��JY��P�I�������7(�)��g=�*�_S�IG�庶ę�w.dP�2�;G^�EK�2�wg{(�l�74�C;h�xo�PF���@k�^�D�����l�#��=In�u����J�(�:jc�e��w�=}�0����yQ�躽���Pb�*����\$pVn�aN�]�Ay��g��h��(�3�4�t.nZʢf�e8X=�x,=U��}"��	�������tH8��o�]�y����Y����B��kLdd�ʣe���@�\AH�F�y���%�2��#P���~q#�v�$�/vլ�@ԾEh�Y;����0�Iֹ��O ��/��s~��v��)��3�ga�EWY�WuP��;\H�����>� ������%�+��Z�l�¿�8~@�q7,�Q��G1#��3��9����QQD}�AO�Fou hn�V=q��'�߮6ǖ��]�ETF�T�"S��x�(�k� �&��Ր"�1Mm8 1�wk��p�8Q�
�AY��Gqv/��^����m,���{o�ts���#ל�AГ<w�/)�r�|�����E�o���+���(��m���:)���+�jfx�0:�q#l�0�r�`�MhP�Mq�#|�P��.�Y�����5��� ��R���W���&G���AˌbNՁ��e.	�㊤YE�|LEj����U,����q�����18͇�53L(�N�Om��K�v�k�R�7�n0ދ}я)i��<���[�G�Ś�q'Z7$�����8����X"����,$��S0?S$�aك�s�vE����R��:��E���m(�w�OWf��O߯�@�`<�Z|D0g�6�����A�?u̹;)��7�U@�t=��.��{��,�A�5mC��\�%�H��P*�q�&�f����5��YOf��J�1b2�k1Hݽ!(�|�%d�ի��#�s.�{�4
�X褣�/(�]�TGr$�M�d��_&��ӿ�Ԍ�ܥj�K=Ӂ&����\σ1�Jbs,:C�k}�:i�/�6v���;%-V�&*�#�r���:��������Lr���y�;ό�l
���.<��r�{�젒�C{�r�] q_X9��-'o�ZƠ�W\�v���L7�a@���i��:Wu��	���/�-ˠ�N�F\]���a~�;<��as�tar�����9�6�� Gm����[���W�Pފe�bu��hҬ���P>�`	�&ð���V��!�I�LdF,��^��jv���f�U"1��`�O?H<2fc�}�΁n��&Wpm�vwO�	��4:��������GTY9ޞ<�n����aw>�_�BPt6�K �p$�19��#wO�!.B� )�I,x�+�5� �j��
�řf %��V��P0���_SbOr������"n��l�I�R)u'2[�V�l��*@��Q5�� v�?��u
��FG�d�_ek��I�/����kM�u_i��Y�w:�e�bv�p.� m��y�����kʛM�s�o�wYF��jnH�Nʚ�|������.��zC����	r�K�����w�1����'oա����D���Vb������~0�B ����+�\��h����1�6������M�C� Kv���?�b��S��!<�L���X��k�.�B�[�q�R�+��:��A���/��Z��<~m��?��\����T���݄4��j���q��g&
:Ѽ������]Z�)n1a�$Ѣ�䲌C�e�0������ӿӾۮ���+�d��/����7�L�Q_;��z;�=/�1~{�)3���U��~q���WP��]t�:",p��C�mA*τ���ʳ:��4a$�G*�2�5��iSA�*|��T�+����nܝ���[����������FP��=:�z������9�#�̣NÊ�ia�
���q~n����g|�f�M��H�8�Q�pd�&˶��*����$�K<%J$�y��8A�x�A_�^Wb\�̨��M�G`����}���	�S
�;���4�>20�v!���L:�KW<��;�˱�a˦�n������.'�md}ӣNg�PF&��&}�)֜�������&c�@Z��4IT|rr�W@��A��\W4�tl�V��a'`�섴R�7|� dn���H��f��*#����f�kTo�_Ƥ�'
�V0�5��(	���
�[Ɗ��n=��.�iy �~���	7 x�%:�+�#��f}
�	;	~�����:�H�P�$G�~ՊZbxب_G;E[�z��m]_�nǄ_&�L���e��6�q���j���㙋ml%V5.��޼�[�2�Ӥ�)��[����Y���T�<�7馴�*��q��]�ԙ�HC�49.yp����A�'`��4�c6�pk c���*׮���e#.woZ�sC�?\gk0^Qre`C����P.ˁ�o(��6�
�+]��;a�Y��8��<_a�����6M�1�o�D��b��"7J�1�|/���]�r�ӾdW�.�����p�|�@
�'C��;oM%lk#�����RDm;A���Y��j��a�����H�N�|�[»aF��jnrVU�l��JX�#��r_zt��*�V�����Q�X5�ܹJ��[/�_w� �����Y�;�<�>h�'�\Cl�d�����\^�T�_1�+r�>*e``<�WH�C������cU���M�Y�T��d*M���K���G�:����h��*H���G��(�t]�;����a�8S����t�{���Kh���߇dFO�
���y�A�I�Lz���BH���K��
���x�l쨥Vt�V�k��8�u��\�k�6��-ZgC�r�fw���	4���� ��aԓ�dwJT�(Ř���JY��)��ن�E��A�%�8�)b�|(
.V���k*[�����E��>9I/N:�uc��HZ��j&L����Yz[u]��m�NV���!�B���������::vtaQߐ�@2�葾�j)j}G�4A�;P�mա�*���ղ��� [-˒�'�ܩ���"dz�y�R`5V�T��p<��%~������+��Yp!;1�y��
Gr)U�������ݙ�#�`�^�`�(�ڄ��E`RGNj=-����2�7�v��@��R���v��*f)�ڨ��܇����������G܅�<�"e��3��z��8�C\K0=ln?��18X$�+���.Y%7�Ny�1!�J0_���j �W��9v.�s4�Y%̘���F2[�K�ɮ*�7i��R�E|}/�<�F�Ą��
B�sf�)mCT���2�\Ҧ1��ם�I��'a�-88����T~�T�/�pG�3��n�R����uF�k7�ly�,���n񕖸Y���@�v�x��b�r����V����,��(9SQӐ�s�J��d��w�-X[Zf}�!�V��O�q�L��:^r?~�����(�^�G���s���=�ǿg�RX����_�)�1W�N�x��whrq#��A8��"Rǟ�$ ݹF��-u��/1�R�C��3�
ޤ(�^�}E��)rL/�Xw���h�G.����W.����U/adQ�b�?���(�O����e�;j�H�͓)��f�k��ˌv^�i�u������d_�h�)r'�[�r�����U�O�'����@ HK���1��W���{W�����ޯ���~���o���U2Ȼ��h�y&��F�?q��Q�xW~rX& |�?�����1�����p�:M%�D.otߟ?WڤB?��������� y~�V!��м�|�p3EʺH�*Ɇ9�1��!,��o���Gg�u�E�V��	���/�T������y�	>����Jff���.��u�	N�l�\�RF�����0����S��C?�l��H�+�%���t�$��st�|��2s�2>&���Ԓ+��3����X%�f)����ˮ[#P��T�ы|ּ�fVs`��Lg[@�$�QwKƠ�H'd'���"0{���d/^�1��z�D�2Vʅ���麣���I�7P�ᲄ���S"�Q+�����p&�y���XeoȉNf�ͥ�]�u���Ĳ�V�f���r�[��9u�6�W�T.���[̧s�����y��C�G��]�h�� ZR `[c3�-�x)��� �������+n�gHJ�����n5� �W~ݩg��ai> ���P��`�L��D�zOz�2�%�AlM:�9�^�bw����Z!��6��8����=j0��3�1"���	�C�Dћf�ī�ʡ)�
����n'"�
��!�^o�g��'l������V�C���s7�칠~t����%W^%i��.�K�>(���9���qZ�Bo^m�gd��m������>���PH�� �� ���~ٹ�9j�h�>����A��U��EXQ�%f�h���״�(~䤂~*�wJ�I �c��Z���5�y�I�_��U�x(�G}gM;����%�$�zx����g0�G	"��k2~/���H]Z�'9�s�6��=�U1>3�}���Uמ~p���c���h/��Q�Hܜf��Ҟ��J`�yv	X4��p��A�����eg����0�[i���J������9/�Ӕ ��`���q���ӝ�3^,�7𩐦���K�O*p/��*�������py���t��Q���h�b=���W3^L�wG����U�q9A�A(�P�I�#�P(��4In�* [������/v��w�',@���V��\�t����KV��M�ۄі�P���t�.`$�N���$�0kfC �ś��)�>O/�=_�8z���^�qsU}�M@����Q�ʝ��њ�Xq;���N�v<O˾�`�p|9GKX�0�G6��|wp\������j���o�Ã��<�,��)S���d�'
Ee�
�a�ǳ��������bJ ��mQ�&?��,%86	Tc�;q(.Tf����PM�<P;'䎏T0��^�wv��G�?^,� �K>��5�T��&k$N�ħ��"��́�t��]�mNͶ-n�騙�6�=Q�)j�	j@�$0P�A�}�uQ$�.F2+�O^��U����'Tyظ�@�����-eB�||ؗ+M���,�ӡ����M&e�8����N�����$��ƥ�����3gǇ���~w����>�����8������p���ۈ亲��0�H(^e��sB�!h��؎J�����;ȯg��I-^�u2�4�n]�
{D��gGv�	���j�Œq  ht$5�1�*���;����!�e|~��.z!y������͌����!A����Ym�!����=^�� w�h�w�E�i{�BgΖ��v�x��l�5��HA��?�B�y������?�\rR�%���n䫙Xm���.�qd����K�3�g�Sa��I�x�f:OŽS�"�ߵ��;g�T��qg�I�2�R�M3饞R�`�*J�m��>_�����~jCJ�uk�6p��i� ��H�Ä�u8&��{C�.���נ�5�cǳ>�n����2.�W�\��<�rV>��R VE�^��(!{��
�&ET��K�k�t� ���؁ug��Hf�>D�-��?�\��#D[����͢~�`����1-�8������=;�u�
�,����	�-�Lw��X]��~�q�pg��2-%H�����D4T� ��L�Wv��Z;���m1�O�M ���5ˎ�m�
G�n#߹v�,���㯆��_}6���(���/�`����>zc(�zU ����_$]�`��a�(�� �>x^Ώ����� ��tY]%+�$oL.���_��A'����{D+��������+s���uI�����Ex�T_]��M�#_#��n�y�����<0�aR�֥�d���:4!���ڳ����Q���B�B��� �X1���N�f��o�V�ts����~tp>O1��D�Q�����6����,-z<܅ ��%R�������$ѵ�v�Y��9q,��B#�Y���{D�y��,�CE�!�Z�_�#��"�d(��=�I���:�8�@�#�dlb�ƴ�P꾝�iX�C�_��U��S_�r�o�E��X{���Z"��ӽ馕��I�B�3m����a�Ce��8�+��Ղ,v����77�"]�#J�����XMm��#	 ��;�˭s@\\z�<�R���+c��?P$�b+0��k]g���Ji��H�_�zH�GM����UI@�yz�<�U
�Ɛ[�>�_�m��8nt%��3�|-�%��8ͷ��aR�~�:�1g�+_�R����Џ��&EzZ_[�<,�X�P`��l, ����c��R�D
B�iM���i>*@���aD�=�yDmg�v�0=�ZŲ�[�Z���"����&�И�EU�����j�i�xWn?�BT�q��AR��w��Q�§��B�39OTygHWK��[��z��_ ���W͙gFpД�7�P?)���6�|�19"���K���)����q�J�l���lJ��F�;K�.��-����ݽ�juk����]D��ã%߲,��<�pE�UX#Bz��H�`��'��B��.����d,p�z͟��g��A��@�q�����,of4���rƐ��FB(N��b���
�m2BO�)�/ᬖY�Re���V���7�x���}!6��$j|�&%���(qMkwxL���p.!��j�$�!?8�Jfl����(M� d3+�iG��L���~y��_�������?1ɓ/ �J� ��sQ��y��z�#VRٌ����Ӑc�X��}��Q��`[�to)�e�K�l��<�c.H ��O�:�9i�w��v�]:������°a�f�۴������A
��-���mI�q/�B�C���AR>�b��I��1s�����طF����EQ�|��	������-\me$g:Q
ݕ:s���@u�t�[iċ��Q=��7�N�	��;+P���D�5�畄��H��V4��F��"C����� �=+�����g\j� |2���<�b&�6���@�j+6���9R|唼��;�E��ǯ+Dʂ�w�|��{Ox���l�ઞ�"j�VW�0 ���+�&&�	��fxF;�W�*�e�o>�O���m@|�AY��/�����
���k���m��aX8��qW�7*<�F1��Y��$��'��	{c_������ ���)2'|3�ј��M��~
`��3ףl�sೆK�ؤ,���,Y̐wUL�W�T��7�[Ip&st��t���_`�Y,Xi�j��GmL�(-l���]Q��`S�Q�5s�RW-{��Aݧ(�Lv1r�]����`��3�r%�3\�
ov��̕�;6|"JS�9�����n=�-eP�]#i�_P}��������Po0Wˣp`D�Iq����:K��O���������!v.g�x,f�!
�rN9��^1������)�� �E��	O��C۹���pIth�_�'�p{B��D2���&t�ȏ��nw�ڛ,Tn�Kх�p��c�_3�L�G?%��	�V�4��eZ�b0_� ���[.@��?��nZ��1��@�p����t����~��sٞ�a��=͞S�*����c���7%qR��pjj��w�-�����_������ɂ�"��MV����uGM��_0��vx��
l�
D=]�o}�-�/� ٤�+��\}���}��o8�r��.ȶ�[��P�騇J2��U�	��^�'B���f���А��z><��d	��O���W���E��MyC��U�f���4j�f����7��|�ZѯS#�o9E��Tr�+C�@�\���e�Qs*7����J���2JJ����}��6��PL^釁��z�|������y�������|'�E�������'�S��@c�.A�J��/�5h����[�������v�@y:\����Yf�A_p��� "�h�K�=U�m��<h�u�N���ܺ��B�5{�i�j�8���5�Y��V����Y�1�!���\O�j���"8�N�>�B�<_�ў��A@,�W��??%j�m��~�<����o"f�&f̑IR�x��"�M�
\m� ���~/�Ȧp3��k4k�V0�ǵ�j5��{+�+��/��03�&CH��&�:�ƿJ�gu�T���#�����<�o}���(�2���Ǿ�������*���[��9KaR�H�ҙ�zY��⯁}�ц�G�[�����ǆBx3���Dim�/���qf�0&5����/��/�~d�1m~]�?�}�v_�C�g>�o�r���#���Z�=�Z��}c��b�3����a�A�^���6�s�㑑'.g��:Ӿ����0z|�ܓ�ַ^��nI������R�fT=�u���NT�y70��_k�YY-��e��7oN�/����N�X�Ki����{V�grǑ�ߓn>x?h[.��f=����^�^T�Xi��^��������DQ�7)3��7���Z*1P`NRє�
�c,[=��J��`6�Ȃ֞(�@�HTp�w��hb�y�h���b�X˝@��YBk����y�Ѥ�����kP��I&��'�:��/�K�&haMG@#�V�qI���&ř�$d�aT���1X&=�2b����8�P!�?7���H���?�����9~��׽[ �q�v���ѽ��7��$���ͺ�L@oK�����*
��>"���P\�o��n�>x��kQi���;�oc�;^�PBhd�/��A"���=��Ԙ���;�&T(��uR�+��1��_>jG������H&Q�/�.�h,�|8��\u}�/`x#�@��5�kw�smK�p��'���r��3ɔ����_�����(T��io�եc��Z'��izg����X������Wp-.�����$C���@��V�[.�$� -}�(��}�`uC��O ���U���ǰ��*�I��l~'K�����p0��&;H��(��C��	e��ؗw̨E������7�#�<�gPũ�o�H�#�i���س��d�j�w���4֯VS�/�������-.�Qw1v_�1�;���Щ~�˷�5{�f:O��TG��(�-ɒ��T���S/�,_>�/�4�>�_�s�(������� ���g�Z׳^�en�D��U�\\V��]�3E���A�d<�$`"��f��_�߳s����