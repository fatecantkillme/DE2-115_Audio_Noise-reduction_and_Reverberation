��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<���=a�bm�kM�#��k�.hJ���s{?)R'#M���ŭ���Yʤ�ϖa~�Ed0&�a��RޭO�*Ar-�xeA�b�Z���(��Y/BhO��ӎ����0뭣��IOi�.��h�P�U)��2Q��)�L��Ԣ�d�u&��%9�]��v��[�O��L�%�DD��/zj��'�Me�	3m6t�+ay��l>lS30w~ݿB��#���-â$����q3���y��
k%!÷�O��qUÚ��}>�\�U/Q�D��>+^����N�~����G���"W�T�`�q�_*���$�e�X����3X��kG[�����O�7�����3e&�ZFK�sL�t�����/?i�1�՛)��PJ�hx޽v�e/���-�EC�[���:��	b��D
;~V��Tў:�f��������<��8�p��!~��*������,7��~��kpq��
�P�=�ޖX�U�}�d=�o\�{�oJ�QB'�=5��/��i��ݕ�75@א���k�Z��P �4>���-#�;�K����V���]eAj)��ɉ�^ꟁA��/H��QoF
y?R�"e�7g������lQ 
3/�\��I5h�fs��W�YM��H΂)�m�C����Oi!f�yWJ���k�s1��43�vޥ�0���fW�M=8pU_9fX��V�sq�4ix|Q��ɰ*"Sb�p�E��1�E��T����������������������5ap$W8��:9���ޝ�.eB��r�w[�_�سWRa�m��4K�;%�f�< ���UN\�N���H��H�A|Z�)�ػG3#��p�@|�P9�KT���l�1D�dA��?f O>��S�E:.5W�����\r�
5�v۴�WOB{�lZ׈b:�}�=p�0���\����<yj%"���*���y�Z.�����S��	�
'��)�6�>@�	:b?oG�>G�um�l�l���&ϥot�A\�'�	�%�Q脗��tR��e^��=��O�lf�)/:0��.D��DY%:�@:�T�#C��S�%-N2��lm/o�A����L�G�cS��X�2DD1{>L9��O]:�'�$p>lW�ޢ�D>SSt�&�G�m��x�+y$�I*N:(;Ԁe��(+����!3Qz�����-*n5�NҺ��e�e���/��8*�.8#��������6kΑ���i��>�M9��ֹ��a�Rc١�y�|��'R�����Ł�*�7d���:we��Z?�no�#O��*́@����&�u�O1�Y}C�\H�G���߫�r6�K�J�'�C���Д~B:��8���P�3h��4�ˑەqCd��x��c��TAl��4|j��[ʛ�`	J=�Wߔ!_;L�,��
�Q���K�-��H+N�n�Y�7�T�Z<��iI�ൠa�n����h�#fi���R��$9�oKQn�Ő��z�岳�a��oۊ�
4�3��&�p�+��fF*{#�FY�F`4#s�O��A��h����cjRLOGv�;(��j�$�p��:_�n��_�)$Vdk�б�L�$���j(wy��1�Gc '�KM	g�x�%� /�9'�;�a��T� �H���nOV����IcHjDB��5��6���b\5O��}����'g�5�3w�;0�{��|�beS^��TJ�OG�fYl�G �{V����8��c����h��?
�>��M�&�'�,�N+"?���7�'�Z<���3i�g�];]1��!h'�p�~�>�U����h'��U��$ �7T�ф�nwL��yi��ߒ����i�����LE�%$��[��!U�b��q���a��MY19=+*3�jO';;]�(�.�d�u���&��~�{�<� �Y�~P��vZ���$�h���*$�#��y�Z#����5kCMv���?4�rm��+S$-��18�� ����q�s�FL���ŷa���j;�9�Ǎ>�#�0*�ر�6ޕ��,l��-E����*a5��t?���2������� 43��z�}���DΫ�k
���4�dC"M?���6�<�
U��8��A�d�ͷQ��ha��P����/es��Q:t{b����󪤛y{t�%U�y�e"	�������@'c�g3-S8�dY�Uwթi�#�O^�Up��c�\E1
�P��b��<�r��rR]ڈ��큔�/5w�p�RÑ}_�a_8>g�5�@%�[��e��0�d����!�#�+�?�LJ�a��JV]2�mL_$g}���M�bU�|ǒ��8����u���=&P&-
��A���5Y��v��[��u������ ����`Y�-ET�}��+A�L��P\T��1̃C�y~M|0�8k'�������ɻ�`�jQ�A�l��Y����5Ý%�f/���=ֶ,��(Ö� M<�ͯ���|�'�K���T8���%��<j(�Y������ͼ9�����x�@�g!#ͳ���4�eD��c�EѢ���Z�2B�o�p�@W�4����{��b�Z�!�ł�>ב�HJ#Q��mP�`�p\fa�X�*�<΍��*�Aa��P��h�K��7���bI�%�Vj�Z�C��U_Ј3�_g��h�~�d#���������O�Ŕ܎�����ع�:��>���y�k����/XA����Ri�%��(x��e�:+��}����K�t��U~i;��UR»���>҂�V.��6H&9Fu�H��XPY��|.�F}��r$b��[ߋ���UE1,B	�,�1!�����}�E�,�7�2WGr�BG����Н�����iwV���yJ#��Kg�dč�x{�#���BGc��!�|�\?�t�PlB��AF��A�k{l�qsn���Z*�諳i�NY�"،���rc8R���J�q��%GL���
FE� ���|�3�#N~&�Q�d��*!l�G�Q*G'���N����a�y�cu1�SW�$�����p�Hqh��������m݄��T({�������ݛ�����EUX�E0PS�ҾX���({k����U��$�B,+�ػ�����������R����)�Dl��M��T���a�}R�:���D���v���͟(�2�����k����tX���_��W.�N1�ǜ8����� 0Շ��u�`�F��]�n�u"r�t�Y2������j������K7s.��a�|fĤ	6�:6�1�Us��G8`�)|�K�ǥ0)a9�f��x�T���S�J��1R�1W�#�2�Є�����7���	�o)��h�T��X�?a�-�7���dD��=���;)[��~�5M-@�C8�v��JP��ȪF�d�ؐ����Jh�����&.LyM��]V�i1��Y������[�ŕ4�y\�7B�3�L�+h,豿�#�����P�;+>�@����/c���H�,��iY6k���w�t��Ki�)1�3�*�?)'�^3�^�vJ�i��'%�b ���'KOE�2�f�:V+���vM��p�C�Ly$��{?r�	>�2j8,�^�7�nk�յ��)%W]�%5�'7�"ܸ-�req�W�)]]tu���{(��<Iܬ?tG�&�'Q�V����.�?��n��
Y��-��%*�*-�5����r�>7���n�-F�*;&.���!���g֚>�ڤ\k�=��\g4^��Q��LqF!p+��(�g)�9�;C����0�0-���(V=T.d346�S�D�M"�K����ye3�'P�s��SU���Bw�8&&ob����0��!���`E���@ ��Ӌ��SG9ሗ�����~�U������Zi���$>XA�jd�(�%�R�u��~�Betj2���@H��H��nC�Bk��S����۽UԻy��OMQ�Y)�~�H|:��<E�#�0��L�Až{����	��}7�Tƪ�qs`��������Z����J#�T���»��I
ڒ��(�Q��n���}_���T.Y�G��v��1��� �ITG�c��TiT]��M?I��O���A}[�*a;�H���t%I�%���6�P���h�[P���4�0855�N:��R����u�u��l6�^P"+�.��}G�/�0��'�X���:A�$��k��ev��(
��Q1��)4��>`�	"�A\�J��ݸjq2�EЇG�o\/?O��z��_�ص�\�6�?���9��D��P ]i�%�eV�3��N��Z�ye�嗼�8^�+�)�H�V4G���B�0(�\���mBb/�%��fH��;��]�{�M����j)y���� 8���ؤ�����}�	ْ(�7����.!Z�PXp��yD�O�3����Y��|�"L�Ҟ�ӽ��>��(�b��V	��탄�B�TF�[|��"��R��c��''@&��w��y�@Jϝ�IC���(+mռ�&�ĭ��њ�3�6߁q�
��E���d&��܈��C�x��f]��.�ű��r[��e���*�L/�|Ȱ)%Z_}���S&��p9$SM�/�=˛;᩶�2B xlMq��FU!���eղ�Nm'�(�SɒQDL�d�����&�Z#8��\�duz��uȁ�h�+�Im�x���H�ԕ�)^+���F��-:�A$&��'ي���.H�"z�֯Ԍ�+��eǬ!����j�̭�(8���;���r�ꐀ�V&�
�s���doi�^V�-��2�O3/�����U��0�xe�n�W���1%���́�)/�`��@��*?����U��� ��O"����it@���l��:�.��<a��|�T|v�?�;n0ɄSg�bh��5I�cǙ�����Zx�+�g����.B�|�����Hb��Q[�:x����;�����tHc���.mO���a$�>����17DT��z5�:3�X�~�CzW\��px�zp黶����c��y�Q����Vy_�T8��_�	��9�x�%��֗�PL�������X�~� �/���7��[67��>�2t�kǰ'���;kH�F��iS�(�
�hIMu��ޓ�ơx�K
��g�{������亭�0�H�(�]�]!`�ZO��,���w��x���.*�[��3A-j����w�EInU*ȹ��R?x=ۯ����֭��d-	�5%�o*�B����W�D�@�?��V��&���f7���$�Cj��VPk�	�/�>0=?�t�j�l�99WLE�&��u��/b.���������l��r��#,����,���W���1F�V4z��Hj�CPK]n?�}A:Jaѧ/�q����ܔcgU2y���f���N�3�"�V��!R7r./��a�#��t<��gP#��^� p���g)�w�S�eR�`D��_^����*ż�+�F	c��a(�(ii���Б1��+sO�"�V�����Wɿ�U6{/_)I0ŕIlK@��`U:�-Xy������
J�B�����k�%Kl�k(U:g_�J�f`�z��+d��c&�D���F�gn�5]|���;po��Vȴ|S� ��� ��B\���{3W ���b�?~ W���>O�-rS�9w�}I�zB��fJg�o�T|�*G��Y�T�s%��I�P�ޡp͢�f*cT5UT>v�:�ّ�`Ѝ��F�X2���(�F@1^��QV:#q�_د���Ÿ�/D]�hl��Z/*�{p׊�-z��i{-�0 WR��������{lgq<9�H�o����[M,���x�7M������7U�-y����R	%�T��83I΂� �+����C2�8�#�^N�L�m����Â��P�Cy�̼�-������<�	��T=���9v��E�ɢ�T�>�ۼ�Cjh����B8��`O�Q��Z%��l�<��b��b��$e]9fȥ������,�"U�6JiI{j��\�d������g��z�V�ڱAi��Ljk���w�&S4������I�q(	�K��*k�[���9��H��y��y��F,�a������bu�D����&�E��v��v񴯱b�5�h��dgQҾ��T�X����];�h��R�}�>U-��*��x�Q��(o�ICˏ+V;���Ԃ�㳝�}ʺpV��"�k�!��f��!�v4�.&�>N���Ӷ��*� �k�9��)�	q���L��2:Yj���{%6��,���,:C(�z�K>����=o(}=�$� f,��I� �u���h���7��i�k�X�ct
6�gY~�%�j���|�.j���f��v��,��mmwU1����%���oK�	η@�W��������_7^�
�$���FbW���$�T0A��w���fP%��Z��u֪�O��, {ls#]u�<�gPjd�g��h�I��`���=ʙ7��b� �����д�>�pF#����bٹ��.��#a�Їƽ����^'�D����O��_�E��OR!}�B2����Ku���h�� �T�����	(��ptgg�Lǜ������P�	���2�^+3Ydy��j5���D�b��0~��%&�͛����R�E<bYŁ/j������F�F6G����-W~	�Ei3\M�7��H�w�ޗ �����未�b�t���� â!�;��N���!Dמկ>�b�G�
 �/6FK��#/�撚P�y�+����?�ܜ�vܙ2��Ё���1a/Ж���ȳij?C�_\]%�� ��i�I^7��aݡ�7��~nSB�n�ɴ� I� ����J6j�/8wZ�a����y�.k�c����Hu=I��Tj�	Ǥ-�9��1RM%Y�Y�)���͌�o�@�,���,1I�H����d���Q�{�{��;߱��g�^c���Ő�����?�[^À��]rfZ���C����+W��3�rP���I1��_� �2BM�Ft�/����V�]n�-l+Ey�=�>DΜu���~�
���Q�S�K�W��`ۮ�Un�e&#^<��I۷>��R}V�<$q��x��=?��Pe�k�-�f�z���pH�Z��V��(����	<ͯ�z�p�a����[���$�[��6dv]?rjs:tuS���	�C��TEXϓ��p�?��β8�Y�.`K�M6g<��MW^�f*iy6'�^�V3sJ*�5.�]���J.���|�A�ai~����U
��X��jGHprC�ö��c�45�L "�4|�2v��+�8Y=m�DMt>�Bn�be\Aa�q�_�^,w�
]T��xk��Fq�V(��<��� 7��OV��������I�K�\�YfD��kF��AP���7ϓ�a�l*�j�SOvp�r�����Z1��7~���9��k]�.�Ռӫ�FЇ��&\X�B�� Cb-���cS�7�����DNW��w�;�.�l1�/]�V��W����12Eb.�d��ёB�ߔ��JmbV"tݖ?��'��(�g���9_.7?޵��y�X#w��T�.<U�5U�1Й'j�䥆=��O��A��|Mi�c`ӛ����o��x�Ηь"�T�����?���2��c6�v\���ˑ��V
گ��G�r�����[/p�x�&(@ef�vPp��~cc�\��."�6�ۗ��z^}
\$��kC�;��-��mZx�8PH��q+U{�������2�pT��w.	e�� �9�*5ơ
S*�-��!-�jG����ј�d��}�՟�<烦xp�(�x؈}1�8�ay8�Zfr,�'���O��aJ���?�����'3��,���X2o��D�+X�w��X�Ё��������>\������ܼ�ą��Y�p^Y\�7yג�"g��E�&B�v1��L@'|&{<(�Nn��BX&8�+��L*&�jL#�+b3���Du�)W!��cO߼��v�1�ϐ=^�b�-9���IO.�刳< �}�M�^�h�6��]z�-��_p�'�K�=>����kӪ��π��m����)E���(�be�6Oa�Z�,{n�Y����փ�,v��$H�<�aRv����PFV/E�*�R�a����>\��y&r{�c��ґﶁYz����;׮�EZOpU��д�6|e8�-E�$���N�n�>��3������&�~�e�c�>~>tT��*>���$k����d��ˊ/�z,��bax�����^O{b�@�n��KK;�A*���ؕ�:�� zB�0bMeWO�fގ��E�"d3~�
���(��Wᥩה�輕N4:�©�@�W�al�b�y<�.i[ar��1����?]W�Y$H�{\|	���/�hܚm07{���s����ǳI���8*@%�7c�$T�?�0=�y���%ն�-9�@���	��7I�k�c���R0?M
c�~?�I�G#Nd�j�Q��z�M�x�M���m�4�UÅej�:�����`i������^}��L����~�l��L� ��Y�J�|�ه��׻���+���u����/V���Q���$ ��'�t}�3&��?2cf.��0rq�< �'k�O
��\(���7[L�G�����: XTX��Mw~cV,;�Ϲ�*gs#�#؜��X�Z���]j_L~$������\E�5�NS5��yLD�O��]Tk�*�\���ݰ_��Qߎw��{_�d�������Nv�� ;��sA'�ʌ�N�$}#
�`t,7f��5c����]���X��-�8QCȟ��)*�U ��ծ\��p��jR��]�S�#,��'?%�|Dh��B����/�\�|r���m���a8o���G�O��L��f�.Jbξ	W
)�,�̻"qm�i�d�� D�