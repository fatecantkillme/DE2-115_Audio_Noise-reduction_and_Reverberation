��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<DU����PG}�
����}�����q5��э? ����&��\��RE�5!�x�.���eOm�\E[ٖ�W��!� d����zD\
�嘽�*me���H�YxsA����S+���6irhz+{Cx�o�(-��9���1�}<�,��,j��}��-Y�@'M�-v#��!�1���ք�g
&�^�����s��F��~tL.��a}��e���р��B -��_��n����ݪ�B7�R:d�-ԷGV6��F��dm�$]}������
\MBw�5@(��a���`XG��g�O�5�����I,�[f��O�nq2��$ti�`��nm�/>1a2�#�К�;�PG�S��E��@��4 ��b/��KF@� :��w��y|�]�6���Y�B�0γ/�!�z��j�KՐ)��(�(���J���R�H���Y��<��smH�fS�}�ʧ�Ȼ&�,l#��1 q\�&����3FCJХ���]md�~�;�}��C,��`�`0����Hė���k^� �&��	禳uF{e[���X�"���o8* `Wu�YN�F����{U���eS�!)�|�'��#��6�IE^�tܚ�f��~�U��4 �FZ��%��]�1Zf'�S�c��q���DK�8M�6���<���ґ)�����+wyw���}��M=O��Q�ħ��ߘ㣃�cF��v-�n$67=�ㄧ1,B)^���}3\�S�}����J��5�����S,�P�6A>!��>�nEJ�Ü���r�b�|��_���AjU�\�7r,�66�<���6������L��Q�
2ȥ���@'�����s�.���]��B�,Ĉv����0b�W��p�������r�楨���Ĉ��#��r����DjD'��ȿ�B(n|"xtL"c��Ox��Kr��1�����`B7[c�w�T��&V8k�ƛ�;{+����e둑zz��#(��/Igwt⃄}s�ݸZ��g�h�U�v��EP|*kW"	q�?�5����j��M7���m�*2�,y"po�M���k��P4�)���A��H[���?��,�rSW������8H"�H�k=
 �C���y���<I�n��*�*"/�!;�M�|M�,��BH���]*:_6&����Ō���]Ǌ`������R��e^%``W5���4�&��ΫFx�9]�:�� d��5���F�$�*E��M3|NO[�So�c��2 ��hZɂ��N$�&އ~^v�b�aq�9�"�V��Hތ��}���c&����:q%Ĝ�o�ٙ����-���&�� r]w.��w��k�bo��Q�y�^�w�cÏ1�-9yY��ynz��~�u�6by�Q%G_&ĻC~�E-�o�7�i`���	�gq��]eNA78���`z�TZ�ͦGY�3볘�>Wt���9��}��7?y^�K�ޖ['�1w5��+�טS�y�w@��2��l$Pp4	sw������qٜ������s�X5�QdJ��Z�C�[�' 
y���"��� ���{�ӕ���n��ۈ��3c[83EE�\�� �<�̜�_�8io��_�ռ;>�(C�AY*)2>�,��5X.@| Br4��b_Iv͗�Bt�d�ד��//�4�Y)�t[Tf�_`綧���cƴ�]��G�/�s�EG���݉��bgF�����Ԟ���=�����Ȃ?��W9{��#,N�7Jm��kFS/�]��ES�g�сߝ�� xd�Hѓ.h%	r���Q�\������쁴鬅�mbi�z���i��~�t)u���2+��[�>ю���!��}�6�+�V���Ѿ@�R��͸�ke�(�XD��A����}������k�۰u�p�۵<���%�X�{��@��Q���J�z�z�,����g��L�4�B���q� j~#����8�a�J�RJَf@�T�r˃b`Q�&���SPC�J�;GUX�;=b��#�v�ϟ�.R�́o���2�s����͕qm��@R� x�[vݱ\}�IoI���,'Ϩ�H�������*���Me%O9�X������2��bW�����XbW=,v#���0�x��M�7^s؆��iЎnDh����{��ӡ���H���o�`�_�IX�����xY��+P�u��4Wg�������5B�b�ۥ@v>~s7������Ģm�ǋ^|$��t�`�������(jX�;�H��TAH�1u1�"Z����_��ؠMˡK�iS�A���'ؕc���CJ����2x�xiW�hN��n�nOLj3�-�+��e�k�?�nyA����������|�TƆ�:��.�[�S���A�qp���K��z'�_-��O��?�Â������eu-<���ʡ�n̄B�2�����M۴��}����V?LH�N��"���5l4�ɠN#��&5.�z�+��eT�+7�C �0�#�%5c�iv^�qy��'�>�'g��A
6�4c��@ǀ}$��'�R0),�(���*S1�xq�RTx���ͥG�#��q�yx
iL�!~�׬���)St�X�_��3�\��tǒ]�	�N?�cr.��H��!<59�v�iPu�;k����75�^�&�M^��)S�����I��q���WD�ZZ ��w�d�q�	ͯ"O5���`����8,O��,��q�*i�W)�2�������Lc���9<��X����A
��ae�^eA�F+�UЖH���'���h��џaV 
���=�K���������N��&7`"���U�'�IJ��q��[�άx����������F�Y���|!��ܪEmP���^5�!x�sO����j�A�z6�4r]�V�����xC�v��~Ê��?����;���%ဋ��y�el��&��\����_���~H8��u��~+l� ;�m4yߩ��Ƞ�O��%���K!�L=f�KxV��:�|�J5M]�o��+')�IAba�m�甋���2�=5R�~,�o��|�w��Ɛ���VT7Q�2bےk<�٫e����641��Bq3���]�Od2�v�d���\'��S=N�+V�n���