��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<Ph���כ��`"���LαL�JM��=�m�um�9^�t�C ��ZT�ar@�|�&��u������?ܞn��h���Y�T6
 �P������L����*8Ԭ7[]��ε�@Z>�7�睠>l�%�R'�����l�IT���w�1R��5]�*��|�4��<5d�#���'(sR��hM���<Ɵ0���i��=�͊dFcH9��-��D�p�uO��e�>�!AmV,b��Z'.]�/���Uz�qoZ�W%���P��9������jS�3�Is(��m0@4�n-����rRe@*���z� �Wt��,7��7,���,���Y��������s�QӁ�`4�y6�L�i����֙�[���'x�V��mv�s$9C��x���4�r{��ɡJ�=�֠��LE���$x�NC\xf�Ib�_bKO���Td����gD4c}U��t<��Uhd����E��^Y�*�9�y�$\O�|C���A�o^y��n�	"/��/�.P!�S*���O8a��&�8�T/O\>���|3=/�H�g��Aul�e���QХ����?���
�?7)Xx.�����ٌ�����u[M1�H���4�Yղ������#t���ѣ�--������v1�\-���fP�ւ�*ү��0SX�Q�M���ҁ.e�)4�R굘��������َ�:'�j�ЭH��:C�Z�)��Je�{ qB����w�& ��v�
���K�H��avVR�aa����d3%�'p�2�����ԭ���.	�v�'sϲ[�����WK�/1��Z.�Jk�7���ϣ~+�z�[X��ٕ�ˮI����.(�04V+8��^1]�3�h ���9�5�=�E(�*��"Cv.!��b��޺�6����"U�u4]f����f���xL 	�T%�G�������/e{�(�__;�_VH$��a��=P�85��RCW�j[+�6f#e�
ę��_�L�?{R�d����*4���������W�c*kIv9�4D�X��՟�s@ʷ��; {_��V��� ��T�X�S�4���?�j��լx ���d	���������c���`ܝ�C���6F
0�b�.��4R+P�(ұ�o��$l$��PUH��G����qL�	�VR�\�ņ�5|�d/k����M��'1�v!ٽB��ȾJ?!� �3]c��7wz�fJKk1�ݕ����AH]�e3y�����-�~�	��Ӄ(5��v���K;�|�3�xp�����!�Y��r�	�n���*V`q���94��!��:���J5���{!�Y�)�i�2�ڇ�i+����<�yٟ�^T�K!�jG3ԃ�4n��Z-��Z#a6�tL*��Vc<�Dc-������؀��FU|�z���a9�>*f{�;��m\}b�nd�w��åL���h]�j�*��,�Rbn�/�(��DD���柅@ 	�0W��#hY���h��-Mw��z߄w��n��)��W��6��l��;Щ�s=L�4N�z��^g���K�}G��e�?�j݅�>q�<�a�eq��i� �gIn������]Ŷ�l��NN4_��Fϗ���>�#��H���>*:܇j��9<^/K�0��I7I��;�Fz��&ԆZ���������	j�/jj�yy�F2�P&q�np��<��ӷ�S׉<C�x���|�fD}u���[��
�zM;DԲQP�-g��:�ԓ��E�"�6xӊXNX�0���2Г.�.5�n]�}�����7.�L��w�(�͐�L�/�~<}x���=�����i�'��#p���Θ%B�M�ƴA�w4��ݗ�D�ʗS�<���P{��3����!���M�����G����ý(]�QsɌ��Y09���H� �M�ˮ�56s^W�;=x�ս��7.���������,K�vJ��n�G�FC�Mk�h��:f�`���Ѧv~��f��>�G�&��,�G*(�Ep5	տ��3�8<�h�L�p�����ۈ�E7�X=I<"�����\Y_��ş�3`���(��y<!g4w9\B�L3!Dt����S����G��Efr�4-�5�)�Q�N����/�|�xg\���:_?��%F��дS`�^8����c�M?�{[��ԅ��Ts}!�����l��{�7� ������.�����%����Ts�4 ކ����2B2R�T�hv�$���dc�[g��h.{����t'0Bs�'b=���	  ��S���w�����ߩpv��\9mvh=g�~W����!Oorݍm>cW�����#��әw���"D���&���;/�/�Y}���8�jz͑����:�;#1�ֱI���s��01��GTp�W�c����5P��W�Zʟۚ��w͵
�6�S�P��g�IjͰPQ,s�xg�������R�fb�K"A3]��Y�2��4�&�
&x*c7��`�m#��]���,NY�<h`'�D?xk"�s�b�k�Eu:��'��k��>��8���(�u�8s�2��Ͻ���r(%g�#�K>M�0��!�Z��c��8������֕�C��Lӳ���3}l����o�h}����@�J��B��J���j�
B�+���PA�"���v�AL��`}�����"UĴ���
9���W��`��!a#�333��4�B�t�e�������?�=��Y�FM��@�0�,�=��X�X�+����8�Ƕ�2�b|�9ir�J\��he���V�*�sp��E�+�@(`H���sE�?��wInBgk�Q梬�ۺ΁E�2��zI����l�pΙ����[���H��H���~�%��(da��:&��C?<��&<�����ȓ5j����U�dm|5�=���Hm �<��8e�ʔt�Y$�b���9����|����oD(��e�n+��|�ɐ���;�s��{WG�̌�4��<�������"b��Z�l_��T�����l�{S����$C���9E��*� �v�l�"e/��Ȯh?�Հ0p�7#�o��ڎ���'�~\�O��� 	�ш�Y�WB���s�[#E���y�L{{-�ܥ��ij��b�05��uC�=�[�i�D��Ar�M�0DI�8j��D���XO	��_�+��EV�/,��z�A�5[H�0+ל�zh���� �i��ϔ��>���g�&����準hz�.��昳�D�n��P(� ���O0����T���]��U�޷_Ui1�j���MC� 
��w�i!���{ٔ���P`1�J+���a���&��7VY��wZ���CF���`�c�� p�3��śh��k�����ma]>�	x0�F���{�,:l-[��O���S�� ��{��~�%ʭdW䓅��-8%�7�w���{�ͫ:�	���>_E&a��7�K�P4��;��&�I��L:M������S�f��ip�D��_t��ھU��p��ؓ�(��1���ԏ|�
��ʸH��5f"�<W)ט���|"t�B��YJM���:���+;�$���o���>
�jF�������7�9ۭ}Js��Y��}�;��I#p�р���r�Gf�c,�?E;���jk^OC��b����RyM
�Y�y�w�i&r���&�9u��G�a�$�eh^Z�{����:��62���U�����c�����e���7Л�t��"d��a�^�d��}�*���<V�~-��Hp��~f�'��0��7�H(�<�g�@ԝ��.aӞb�<�v�)��3蟘HX�f����I�������*����n�z�=t8ëQ�-��wlJ�Z��D�F�	��c�% m�*>�j��<ބ,ٽ7�������o˧B�V���<��I����x�9���7�h�qmy߃�v�����J�{��,�J�퐿�)��A�ݙsnܿAI���w B<���nm��u%&�/�5��v�b�,|13R�v�!?9|�|c;Q�	rB+��d�;��7uPK���~0,��= ����L����?��G�bN�B�Y�Ө���i,J�dH�5�Gk���aV�DJ���
��;ݲ.4�_�4�[�4�)R�fv�R���\�ˡ����+�yIM�V�O�i��{�
����݀�P@�	Ld-¢�'����E�k>���颩�.!e:��8�$n��:�����<��Q�{���)u*��X<Wų62y5I�>u9�?�!mQjQX�#��ZY�O(���V G��#A��иK�Rg�H��K�5@��5�`��v���x���Yv<{�;-yF]�g�!`��bܕ��?�`n�o��s?�ŴW�vC%���<fF2�ӆ5���o]x"�'s
�3�z_��ME<�F�6�8ƍ�J�X�s�x5��7�N��^LG ?�l��Ȃ�
{(Vg-#���Va,�)�bq�$�!n��pD����j�uU��|�V�땩{��J�D��ݾ@�[�]G>�^e涃��S���z~�H�rtMX�����_f��B�#E���6{��3���=�λ���ff�,��e�x�X ��JqO-��QC��I���ƦvX�-������F'��Xk҉�QMs�uZ+�2�%Nxi�N;Y!*oL�&� ���&w[�����gle��tXԹ�Q��K��@�mײ*���^*���c���p��7�0��f
���!��S_+M��=�?�e�Kd�VɁ��	�P:\U԰Y��nڡW�>"�g?v�=��AN�S��j��'GF=a���!�#�KG�oW4�֜����6bJj������y�퍚���	��9���H� �5��w��\rs��C- �Da*a�L��R�YAw�=d��4�?�o�8O!1��0����`�4��c���'n����u�T����} df{܏�e��I�������۵���d<6Y�u?<��1v���B������$�8�j����"k�R��b�DD������[ٴ�fmQI�Z0�U�հw��������A9[+��3.O]E�R�=+�㖱��7�M hC��]D����d���-���n̯�DB��#Ϗ���cJ�B����LaZ�����y>Dp�g0R�S����!�͉wKt�Xp�����Ȳ�˅�q���RֆUj�~�EG�YwMU r�hG��{b�!)�y�R�~RɅbj�ƍﱹ�,��t�ZW%�v�$ш�g?���l������K�H���!K�` ��a�s�"RD��>i�|n���*Q�(~�&�=��y�a�&�Λ;|����	3WK�����?J��$C�զ�	���Q/��##����M7���R,��ޮ��_��\�*+z���t=c�0��S&�4�|�U�Q�v�{>.�^�N��(���B�~IlQ���%E�Es-?}Z{��X�8��e�hYl5��!�M2�ّ?�858p��m�t�-v�X��1��W�����llP��I�S��v���׵��
�\=}qM���C*����|�g���@��I������ZQ^|)���h�ɍ�)��Jz�yU�%��v��܀l0#a���uFc�5A6�.��#�p�$ u���j��Gy%ߩ�C��50:zm`�U�{��6��wA�]� ��߂	4�^L0�篷��a�W �3ۄ��&߂!"$|�+q��rD����{���c��J2�:�Ep�`���1>�W��FŪ�lZkv�K���K����=�+C����h�*���$vQ+��$O��;�g&6w]|�Q����Fѥl��z��ԇ�{F؝N^�����C�W/zM9�O� J��P�bN�w�"P.~��������n��?�<0����D���(j�)DZ��6�B�k%~�I��ඥP~x�-B�{wk���r�0�Ċ�M=�w9���יB�j#����o���(:�p��1XM���hU�CZ�2˦�- �1�]<���$��.\���#R�Z��~���|!к,9$g�-ð�.3��J��َb�x_�KD��e���c�E��~�S�l"�[�9?y��T� ^G�6a�g���������3�y�\���m='ر��QHuj!>6�c�%�,��Q2ķ��poE7B9\Vv��X��b���l$v���܏��L[@�9ApǄ�u	���= qa�A�qnHiAfmG�S�fh.j��|�T���T�LɊ��NS�z� �D��F�2/��tY��V��%}���V�6�B8���<ubmi�������6k�Gg�؁�bm��I��n�0�~�گ�آ��@�cH�79����O��S=�Ack��2"k�j�Ɩ��@=lou��7�jW;�i�;S��P���ū��ǳ���28��MdF���� �48���ɠiFg�N�ջx�6iq� ��U��׶�C��&�2�݅��k�2<�]�5�~�W�l(��o!�`v��Ůx��up��`FU���o]�[��G��Z$�0g|����q�x��x��5�BFb���ٛ���hк���RV��mU��Fq���>�IcB0��K�<!��8�)<�	�>p��{�<�ҽ���9�@BB?>�O"�nj2Dh�ׄ͗u���+-I��OR���8�ᝪ���rڄb/0��H]KS�{����V�*��_�.���V�<�� ���ذ��Rj=��zإ1OJ�qK�/�z����Ԧ��Y��S}�U����L)LS9y�al�T&�X���U����$|o/F��<��FX?1�HC@KQӤq���_�6T��I�#z'(�TM��m:00U��{�x��G�b_Ň)��It@��&�b����c�/L���;͈٘F&*�~��\E��?[�q ?��96A�b����C|�a_�;���Z�jE����L�����W�D��J���ˇ_(�44�`m��^����3#Trʃ�e7o`�9��g�	�ܷZ��<�}��h���g�N��)�E�l�Z����Lb&��+�܌[�b�t9�B�f�2f`Nߓ�
1
"G
��J�P�Y󈸛� d�M=����q:6{�o?�>D6�iiM�;$�E��?���EzH�M�i׋[�֏�E��>!Ifq,8s>x���5!��7��Q�ϙf���Fs�yٵ������%�x� ��V�z�苫B=cXnf�9�&�ʽ�Wx�G��7���Qs�s����#������N����|X�1[���w�v����Er�Dh�0m��X�)�\�v$��}�v�Sp����X�f^o��ѝO^����Y��P��1ƴ�0�Š��71y�W5I�FBh/\z"�dw�0b���g��v�9��xء٦C�LƸpz�:V���M���Wh�!<.x���@�ޙ��;8h]U�n��^%��0�&�����A61��t��Wt�0$a�=��J�ܘ�)h(�T�&�ڢ��_�
1i�Ⱦ-B��@�q�`("��jE�
�<��D��N���,#�۲�aZ�o�6M���8��&��m�r�d7�B֤�gh�6
�hk���
��8|��L�K.�o��H Y�2փ8t���Dx;j�9��B��0�WpÝD��t_��>�}�î�U�R7�:��Rh%e}��G��+zI���P��||qb �������������3���%�H���(UbBw�/�:n7h����LvM��g�*�Y�x0�f�a��8�4~��3�sVJ/��6�xːEh�{@����Ds��a�f�S`+,�he�H~���Ps���-ܓ���P��C("e�߱g:P�GÕ.��8�c\s��HW��ځ��c\�mG�
�Y�(s�:�Ҵ�Jd�D;_�j���(>�,h���a>^��X�k*�[�j���oh���Ev"�{��j@��%���?A����`/�07[?p��%��!� &X��#�D�(xd����D5Y<��[����K@������-����c���Y����k�8h�.�i�횮o�ȧAG�]��[CI}���[���]��S�48n�{�K�=�0[��k)��c��������(��&]�Df���V\��)�Z�Xa)9�z�x,��I�$��������Z��3��f5g�xhj�������=L��i?L~+Y��p��B�
���X^����l��	Qa�Hߢ���G��]�s#yIb�o�z�$�f���6zp�4:&�Ӟ���}� ���9 �X�i;�y>��i�{�@^�|H-F�Z?���W�a'z[Aӡ�::foX5�����ε�RIΤ��g�O3L� {}�I^jB� ������;��_��n�g��*uVw��,	�G�N"b�3�8լ,�9El9=%p�c�:��|2��e��$�:1B�aX89h3����ົgzv��4~@"'�N+��ncqwP�f��3V~U&ߣ��7��n�{@�{5�9��Wf%���h�}�˧�Y��U�OA�s�s3�G������/LD�,�p��l��pk���┄����b�7%5�7
D������X���5fu2L��NkGȄ�
=ǓK��z�UO��d��C�N`w.����s��3<�n.�A�a�����g��,Y'�E��R7��0S2�$"v!�F����r���w<#a~O6��UH�n��4I��ZA�.M�@J7�q�0���ɠ^(���r��\�WPt5G�8fU�Pf�(f|a���?����S���Q��F�j�\c �֭�3G+pd~�Sj&x������Ĭ�r^�b��ĊkV�K�2�op~����j��F)�Ӱ�j:�A��PW<d��}�)���4F�4ŦsKJL	��1f�\�^hִN��k��P7�wW�+�GH���%��a8���G���aS�� ��*
Y�������on�K���*_D�� xT�z4�`��E��Ĳ|��I�'�yʹF4���S@k��ډ�B���c��K�[[@CaB��^��z�Qt�B��h/����6�>TWܤ�\�ْ�z�w���<���Os�L�5����c�$������hNl����|}���:�N2qב�(Il��ts��-�zs���u�al�9�8<%ï܈]�R��{��x1g�g�QO��F
6�M�;N��¿F2�� �,�!��zYĔ����9"�oC���<T\ZNW>j��(���Y�1<���i4�@�d�ud�ְYF��50�
�3�$0�)}��$�u�"Ug:�o[HW���@���*gۇn]䟽��Ɂ���� �fp�؈�Op�>���d?��i�>�̅;��P�A����Tl2s�d������C��(����rOի�zs��L���+��遑N�V_�3s����#��B>B4�/L����w�P��������0�l{��B9_ѺG��eK�,�oj�8� 0�m i�������7?&H��wΚ��h�K�X��|�Ӕ����Nd�@s/f`c�3v���;Wj�1�][��E��Ν������׽[^�0B�{O��<�j�߫�g��rz�G�b��(� P%�#����Ì��!f�q�#�Z΁y��k�[����ߖ�淠��w
	�����O�޹�R,�Z����Z@9d_o�k��{��?��?���ᖀB�sf05{+G;�G �xkT�(Z-gW�;��]�z���E�^��Ok��aLg�DnoV�*)������џ����/�j�{��w�YUL�xBuP�V.cY �鄝:���=��#��aDC��u��:�G�|l������A_zLG9��ۀ�K�(K�Wj�E~�D�݉�`L�|��3��1�BT��p��Yؼ��uS!eпh��=�Aہ�qF�����$�-, �;�(-�S#w�r�J�\C�T���[��m<͌%��k_K�Z�|7q,��ᜳ멕lu��[�y)YA^�~�+ g����PH�ßx���]�9�:���(o���28Q#�=:^SG�"{�����צ1ȯL���'���$��oGO�W�-��H|�<�	D�����
H=�\|m��$���l׎���&\�}a�Y�f+�Z.�3�|B�
��](��L�{B����o
����/���P�ZU� ��4���%6�< lkg�L?�p3zz�#��L��)n�R���~�H���N`�4,tv)(��d0!F���X�.tv�ٙ<,���{�9I��#���Mk�Mǰ�Ѓ߬�J�90w1ˆ.�"��H�K�̈́@��k�D+O8����g&,<sK�*.I��Y���TQ�4�K��Hn��p��Eq�Ҝ:�v"w��W5�c��tALi+	˿����=�j�
Z� �HX�3����q=�8Kv��*Z�h�)j�S,P��+؁���A��S��g��
wMu�f�`:M�8wM%�Os|��Ń��/V>4㵡#��<����~l[��E4L�n����t�\�����ٮP�z�����;�$����gEd �?W�n��l�@�צ�R��	�.=��7�i%Ey�"Ia ;X?A�}��]@a�l�>hkz~�5����n궞x��eVy9Mq�x���mHH�U&�@@��X�+��MG�����di%?Z�p�Ajp�>���ٴ���Ty*�G�������`��9���9��t^V�球��-�!�jn��-��N�ˆ�j��:X��З���Sa��R��E��
�?�)aE��(,Бt,�!{� ���1��Y��܉Vz}��u�SuÜ��e�,ls��W��a�#ɏ;�2�&6�	/\2i�|�\���.�=5|REq%75\��0��K�wk4���Vu,�����ȭE|����_�&����r�Cp:�uaϤ4]h/�ZNՁ;_eG���W��ր�b�����{�[h�Y��s�g߹��a�a����?z��cj�����:`@;���Hھv��c���h������b�D.��p��{6�$#�݄ۼ'5�M����z�}�j*�Ԡjα�^P�>QC5~�B8��8�7�`/VC����o��� ;y����0)+�9a1�:O�/O������	PT�<��	���d�?�f�![���'�&X2'�jVF1s���˶ �t�����_K���?\���:^��v��I��;�l;^`�i�"{�����K���y����U�r�ʆu-p��s��ְ��JB&_�%� ġh��J�W��m����C9^�|����s1X\�_u�GP/;�կ�ָ��,�.��+�P��f��N���rl�٫�{�l�>v�Z+�
=c"�d�X�s��A���E-k���Jt��=�BC��Uh�a�s0H��J�y`r�<ZxSk�>��2��;+.�:�V%�)��tLu��8��i���
 ��leAw6�����>����N�L�ѱz�E\�cg���B���"j�DF���m��4Ż���+�`4��5�h�m#�\�;�ilHZ�u��~y��;A�^��E���K��O8]��1D�F�b����J�}y�L\�
. ¹"�
p>�=�T��l�l�|V�h���-�!�W)ٻ�����A���A[�zk!�7=�<w�	Ֆe@�:��d|�'�l�_z�UHUZ5�,a>!�B����߁��F���,W��~��j�:��,C�5!y�^p�-WH�8b�3���$p��1�q�8&����6u��!L�i�Q� e�x�[�%}O bc��A�3�M�o7���Y��.�5�o�ӫ���/ue�ɍ�ͮ���v����� @Kj/���"'������0c���ڔ)�qS���|����7(m��oL�
.��ٟ�����i��cVahe&'b�x�X������a�aS��]eH��5n�����Z�Z)C7�H��Vg�"=5�3�L���M�� [��z˞F[T�cT	�z[�!+o��Plz�&�,4V��eyD�.q5f!�Ğ�u"��e�I�5
`L��u���TaVd+ǽ*,� �Ε���h�~y�W(ur�~���4f�
P��a��M�N���������@Y�`1v���{k��+%���e���1q��ع���wq�\�0Le4�ˏ��9N�z���b�fd���2[8�(�q���ز�z�v�Z[�԰3��� ��3|4I#26���ۀ81��nS���9S���"��4G/��?����99��4��p鄭��]d�LX�˓�Q7K���;X���`S��bT��F����gJ�w(<$/�	*J���$�%���S�d��\���Y1��~{�u���l�4��*�X-�'x�����Do�>AKS`���S��'�7��~d���\�|�S}��Ji��*ܯL�ި�*��4Tp���pFֆ��}_��������]D/�2oq�nE�ថ���b/<cq�|
&�+^�"�o��sV;S*�2=֞�\��∂w�h�6�8T/�
��=�$Ց3��g`�Ms7l4\͖]F�J��d�z���ۊ��!G�'s�7f�e+_�

K+�m��Ġo��X6��2��]�ET��t �^ �~&�
��$���-L��:5M>���<T�
���P���cw� ���ٖ�믣H�؏_���(��keesP��JF����f��oD ��$�-���"��a�� ���e;��>�� �2���V=���n�i�HOm6����[��a���0��P�4�Ȭ�����/�w1��L߶7W��]��#��R-�����ŭW�s�I�>N�
4��	L��v._CR�=7{U�r��G�Y�1 �ռv���Q�g�é�3�?c:��T�V����A�(�87�]k�n���y�
zE������G-˚U�J9�&��e������3b�V_4��x#	$��"d!ŎO����ɠ6s���%ȁ�[L��<ɏ�G�/Y�u��:�HH��؆Q���A,Gw����Q"�W�l�ֺ�2�)&+A)f>'�O�%��	]�d�����JjǶ�ݱA���b?���6��#��oɱk�T�M��C8�Gp�C�?����g		u�H�[Q�͂�x�?,n�/�a�X���rr�̬�k�?\)r�t�R��94!�"��f�@�+�o<}�sP*td�b�̠��׋&�`@ұ;����>�����گ��',(bw�(��Sh+0�5ҡDz����?M���V��H(�Uu�m�R3��a�A��Cr[���	|7�[�u��y�������#�� ��7`���Yv�t:Z�E��	L��8���P"D+��n��wr��9Q#��/Ư����/��<�b�C5��C$�yF����[FMrH@��,y��@<�g��-dĀ�y���~S�dT���=
�XrFtiG'�>vZ��<��iH,��#���i���J��d���|��sz<[q�\�O���ƙ�d,�-�"�|��ͷ��1��{�����r,��#��A. ��[J���;`}:Cs�i�]�"!E���z���i�cz{�R�1����4���Ϗ~\Hi�X�3TJ�n�;����c���ls_��Zah��&ɟ��U�����H��t�K^���Fd�x�$9�J��#xt&�k�\���6e��0��<��7�w��4�-���M{�6�Vd��81� �ѤW[,0�T��;���
vȀ�u�F�!��*Fðh�.����1ď#�=�#���Wd�/�+{[~7Q;�<g�����`"���������kyKAo"��lB5LK�Y�#C,x����3DSZ��|͎M�M����~���V��	V�/�����	Ta?|�v��bLjS�+��p�<\_&	,H5�xף�@��=3���M��T�dc�C@�Pv�{F'�VJ�U�1�˲���K�p�k�1_b�v��M��S9�/�I�;j͡U~G��ޭrA����JG��Y?�3o��X���Z|4�qի�4V���L92�����AK݃�i.@�k��#2��g6��4���p\�ٌ��_�cilx��r��xk�8�L�����7S&n�aLnk�C����r$bMCi��<�F�"E�TrK������jh7���*���s���~���X$����_�'����]�Z�W��˅h�9R��`�^� y@c��	��9 T� e��q�������1���>9�Q�R<�i����3�v�Mp�P�/.�d�"�ц�3�k?p��{����ܐ��3�,%_c��G(��Cy�"�z	p��d�%/�}*~m�>���W3��(f�w-�E.��>�W�v!� F�-DW�ߘ���E7*���K��|3e�Cw�m�����I�����"������MN���ٱ���}�k7D@~�j�F������J4��Zlfv"W՞Si��p���KI7M�a��;$�F�����F�^�V�\��e�_F����ɳ5�CV��Y�۷���W8�IavI�#۫�V,�ɍì�o{�՟�,,�����R�U��R~7�����^->p���2W��Y6��/���`�[���U�;y}J�S �Z�P�i�G�t� ]�U=9�f �8�������es��^�f �r����de!��A�}�w1��{��hY��E�8�;�
T�~D$6?�Nq�Ϙ��nȖ�1c��؉�H�7������!���k����#��c`����i�� �@e�S�X1%F�j:f��EI+��E�#5D�Q�
�ȩ{�~݊�n�$�������4p]栛�12�ֳ���:�AP\^�W}By0F%�"�k�u��ހ�B��hO���K�� wэ8�:D'k��:9�1e��)�<.B�����SU�8��>���a��K(aY�|&�)��cg�8/�@+�������Y���{>���*݁$ 6�Y��|a&$X�߆�=,�6���=t'ݪTo�`o�>����d<�l?��`w4E����8�%���DHw%����}X���۬���z V�	�k%F��P�1S�7�����k��#�����2��| �u�3�;u4G���'�B�>S�3?3�um!y�(��B����*��F"����o�h����T�=���F��aD�:����^�2o�*���h�2����h]9�!���� �������bk�{z|h+M��lE�����5���r��]�ᬊ]u��h�Ϥ�+(����n����{��ĕ��G	A�vba�f[�Ȯ6��R�FGG�"�%4�^�[67l�����v;���PK�N1]�L���a3j�k���j�s)����6�t�	*={���Y���[Ws�6�}Y�0��-�\�3Jٝކm��MU��qֶ�}�.��Y��!\+N\Y�1�� Ј;�� v n�
��Ɲ�^�m	�(�-��>��Wo�ᘶP�-Zb�1�&��6�-X�y��P���,��d3�r���}��2x���`�ş���̙RS{�֔��5��*D֦q��9S����4���ꤗ�͎���e@�=^q A:����v\�h4�sP�|Vh�	d�q�+�Ŧ����i4,Q����FC��|Q�ŇH�Z�~פ4� ËjR�,��w̹���v���A���W��.��L�uW���+sl��{λ��M��8�Oע1|�g=I ��+ȇb�{'31˒��~4�W�$�O'��uw@�o
Q�7�Z�b�W��'�xB[�\]m��j�/��0��+�q�_r���B��Î�H8o�L8|����}3�NzS;�ؤ���2��k����A�0�٤P��� 2�퐪T�;��p����>_�Hd��F���v�Wq|B��T1�	 tB8�Dˇ`c�.iw!e���u��`�t�S��D��ӕ��-B�#�V�OQ����G)��Jf(\i#^���������!���H�,Jq�ƹyL'�����2��GK1�Mtv˚�	s��"r�%�Łx=qzh0?5R��cY S"�R��o��{xƁ��'Q��ƚ٠��<>+�[��j.��r��>b� P��F&qr�g<���djڬa�ĩ}�1y�
��"�.`ή���9YK�A���l!	��6鼜�<��-^aO>�1���v��9c)L'	���+r�dvv�1�����	���"O��Dt�
v��蔌���0��{(=��W��$UłK��-���w@�E��:��PK�!�J�i<��נ���+����+�X$/��G�qݱ�FQ ~��������r���5��,f-ސt?������se}�����8PR�v�1�S4��IG7s�Fu6������6u㎳-�>'!�e������2av���{��r�Q���c��xvZ��I�٪ﬨ�6-SDu/��h9}�AQ�6)�ma<j)ɏtw�k�):,eAl��,şe���YUi�@tK���4��?�'�"O�ڍt�w�+Jk1� 	�j��EM�~�9��cCC��\.>s�����h�}�sf�ɛN�XZQb�����0�����z�,�kIJ�2-��o�1p���7���m����E!
M�����󋔴Ǚ�ď�	ۜ-Ge3�=B��s�W���e{_5۸�;�Y���?q=
�쓽�Ƴ������6��(���ee��]b����5��®<:�u8*��I�.�-��{�к�Z9}�/�7�٦���O�٠��y�%��͏qÖ!M�F$#�Rڈ"�7zS�+��+�]��,�%�dw��o|�)�
���Qa���̩��V��|�LAx�,�p~���f:0��ƭ
�Կ�*I������V����!�re[�l@;��q-u��n�ڀ!@I�{������)	Æ�������R���;osZ�=�����g��],4C��}�]o����fo����YG�
&$�q�6TT�bЀʛ�-*��~��\��\�9`p�����K�r��.�p\����X��#�  �)	t&.�,V����M�C���%}�����VZH�>#̷�86��sq��~��Y��Zu��V����R������ϻ7�v�/GZ|%�X��)�qx�g�d��-����K(��|�
F���@����x�0�Ï��&�I�t/���H�e��"K����uq�d���L��뀰��,�Υj��),�G�Qp�O�/��3�p7��!�Wv��5�Û8��ɕ�t����e���hp�8�U�<�djB��J�,?���$D¾������|�߀!:���d깃���l\	�,T	xp����A��BeU����y&�I����,�f�N����1m���S�Diҗp��j��Z1 �.xu*��F��H�K�'ى�R/�<Y�p~��/�?����(�;���K�o^�fd�*άL[C��	Ė�K����c�?\��^_"F!�00Yc�3ɹa�1�x�Tp�A���ƖU����e���`@?W~�ֱ���	�$��l����A���M�r��ȑ�$�jد̶T���)�ߎ�:ZǮ��>��LV}�"��^��՗%z��(y����}�#R� z�^�]������wSZ����_ğ�Y#�v����X
܇:�x�;��������2������_�O�]I��	?��w�_{�A�e�>�&<n������k*�z�gk�`h93?�[1�yŖ�B&6 t�s{�Ug�Ooю5��%�X ��w0����L�d�]��\�8M�`
�����Ĝ��߽�jGI]
lV K�>����ط�=8�U��>qvg;4Do�5P������`�$_���֫!�����E���$I&@���q!����Ƙo�������e;��[J�'�ƞ�x���:T>�-�G�	S�����A������7:MH�n��HȪ[���/�"t�o{��)�Ю}���O�U�di��;�'n`GA���B�
���FF�4�.�����f	�G��6m����wd�[��(�b�w.�
L"����S�8�vP�����#^?����X�6ً؟:�]X�KT�,��� &�3@Dn�����l>����೎�Տ�� W_eC��C�ԉf��q;�܍�"S7PR���)�ܾ-��˭��l]�OW~����Ԓ�L���l��Y�T�%q���7��נO��(7�w��4C�eb"W��4\�'j
�dޜ�~k�<����R��А�0����Z��3V/=	ha�Cܢ�l\�O��_A���0&�k	%�?S�~���$�����U���]�OC4��=��u.t�L3����E�f�\ҭ�?���o��l4*m�f�!x�f2���%C�ڤ<�·]��v9gz0��&�np~��S��h�&��@�}50F௯V�Y��15�3����gs��Bb��c�x��6wƳ��kh���Go�1�������e֘��h{Z��2��o�@�Y��N{9n��t��B/H,�0�/.��Ȭ5��.��3�%��ztC����
kD�l՝��}�;��JfE���� o�ʻ�+��ȔIP�a��m���%��[/c�u��3�V8�Z�0����m
}�Y�pP �����3�t�!�e�}�"�(���xꩧ��y��l��BLL|4��:m�0|��D�)526�ٟ*O~�qݾHP͝� �*��5�&��=�o�Y���D�&�qn%Y����>4C'sR����V7��͕�?��S�j�#���~��7Q�o6. �N(p_E���������F,�v ����fWT*�='��?XB�sN"�Xy]�P�����A�ecn�A��9���C�4G��:��!�{/0%�Y��8b�0��X*72�!S։htya���2�ri��h�k� {Ҥ���SHE�0hx,*$E�,��lE��m�4���-�N3����>�� �J�.2G��~��� 
�}���;�'v��(��Cݕr9}L�'u}��iW4��s����0�h? �3j�S�yQ\�55��9�l�:��ۧ�$$Q�¸Q�-�4����g�R���PM���>O=��8i�XW�*E��ĳ97��D���m��Px|�'���c��Nyl��~�R����p,1�D��L����La�ϰ��S_!y_]w���Hs���C7���d�ݦW2���џr2EͲ� ��E��65,9����5/�uє�y�/<Z���V��@@�ېkp͞(ʇ�)�WP��]И2���Ku�uz_��s��:壇P����~���wN��8���PA;
MR׊���,w>z(A�M7�#��h���(f��z����m3�����Q#��}K,|�>M�)iK�����y���W�7��b�w�K���\bH����,����9�^���d�m��$�c9j줭�(��Z'[��9'ygDL���=Vcy�	��Ն;b��Y$��]�Z�r�#��?�)�);g�9iG��<�K�^O�>C�b�`�)~ݦ��#���X�<~}z��+s!*~v�
/�Љ���Y	�(2�t���+�f��I��s ]��u�22�H*8����z�Q�U-F,u��.r��o�U����I�Č-R�_e�B=��x������ۇ9Wi�x�zIP1��otG,�ĩ��ɫ��n��1Ğ��i�5�0��&m��3�JD�DI�.v{��p�R (K���`xçN;O�*�& �"��=gj�˅�u���Bכ�0�"����b㒔Ծ�};V�K�IP_RТ�yX��Oo�a9满�z=�0L~�E��� `�n��%�H��$i4���>�5K[�]�U_�
�_�QJ�~DK�e���t� ���4=n��p?������26��Ў�ɤ�7:r>%&զ���#W�u���\	L(ڊ�g�����Ėg���=�&r�~���(�	_���e�
�2�/A|�V=�م�2lm믥z�ܪo_~kHӷb�IX�9����	��*�/&29O��w �����=�K?|̐��"[�{��d=c!�<�N[�sJ�M���X�J�x��WB<�\uk�W�2?���S;���e	�f2�v%�Xjd�P�R�x�P��8�<����n��Üy��ޞnV0��3^I�Jq�\Uf�1�����,�K�z�v�.�fx�Lk���������4�$mO'��}\��LxI�_uL�!�Q�O%�pt$�����2�l��$�� 8&]�*yͭ���/�(V�s���J�g��g�-��q�d�����)q!G�8����A^��hG�C�D	���X����˫��-����Q���L;0���~�2�Z�c-'Gm��IT�%���W�W
Hi�Jފ�*?���z�?p�J�
�w�P�0ЗH�p�su�H�����aHE`�6JR��%'X"��_ퟯ�mQ�$,Ye�߀uT9�j�\��/LC�VD� ��TbG�+�������u�X���Z"���K�`٣��	����(@��"�����߽��k�X��Y��.��/��	!�n�85�3�����1;�&��:��lޓ����P�$$ZG�O6���ZE����y� t9�Ku՝#S��
�������ڎ��(c4��:Co6Yhpo�4j(�P�+�5U=b�����ͧ|�(cC�n��OK��e�	��#8Y�l�ۥ��3����S��R��h�����|2���Vdyj�3��V~���P:_�g.$�Vёԥ" 98��	ƜN�M���N�D�?� 
�1*z
6���L�=��	I�/F��(/U�Cav���ㅂy����de�Z���¿�Hp��9��*����0zj�r'x�=_��U%�n6���:%lm>�?Y� ,v��]�a�
�N�c��'WJ[�٫a�ӷF��g�Hp$3Y�\�޽��d��
�<�z�ܽ\�3Stգ]�Q�~��	t���W�Y5�!헰e{��Ŝ�
�Pq��БoV���RY&�.�A�݊���U:PS)�H|<���@��&�ᖘ��?y��+�P�T���v_����5��Z�Y�g� ��F}�;�('�W�3h�E�m�B����LJ������{����A�s�,�����f5s{�Xq�%a�{�%���<O���.�w�3�ϫ�*�M��A�cp��2�T�׌�+]g��"pg��H�P���a����q|���L^p@�t+H�v�r2�f�fo���_��ŏzU�[�����1g���I� 9nB��X�u;&F����8����2�e����Y���TE��A�Ƀ��ڒ��S��87T�����!�x���r�IQ�]���zW �T3��p���N�bs Da�}yx6����J�-҄���L7 )�`P�p�� f)�D!NK%ۿz�c���q6�gl<��nC���j��4�?~yV8�L����ꚡ2�P� �TI{�r{_I��_�U�]���Lp�%���D����!�y���ҦI�Ʌ?���hFܠF^K�p���1�_�]��?:���\A��716�oԎN���Ǎ�Q�b����M��Ǿ��]q�r�Ш}��r�3���l�,��� �kfp����깟�C*������㳜�e<���.��@������[�Hy ��q��dX�Tt4�Z��.�A�l(Z�,�$S�8TkDR�GC���Nk�8���.3%�]� -�����R���*S�,\�d�#n�D\����X�
R��F��𺻲�{��5\	ϝу���YKk	�����
�wUn���s�.p�@� �u�I�C�F%u_�;'0QU'�)A==	 "@G��6��4�:�ecҠN��0�nT���?Bt�F}�e���{\繍��a�r�C�/����l;�n���X�[�w@�d��X����MxI��1vR��t���-U}-E�)��Nnd_b}�"-��j���!t�N��6��~��Z���=m'����f�|�'��6�F|�7"�_*{�5e-BS��F�
�X�f��?��;	뵪 Ům�ׯ��/<��h��4j8P�#5��ض�6q�Ka
�N���{�����<J�/����+��8��h�O�4����"�X��; ��uJ��}I4�����Y
�6Ss��,���Х޷�!K�s����"Iv��Q�O�<�5���0�*]�g����qP�;? z�!ƭ&�+5$<V[4;R
�U�\��M���l��d�+F�xP���$E� Qg"�sjAlçB���*��'�$�8W\��lX���1� �(j��?38_�g@�v��1P��3�4�-98-
� 0Nz�]�f"�|��
�i��#n�$l�(f�l�RQ޷�]C6����&���՜I{>UK�e*�-*�n8:��;z%�{~��+S�:����Mچ""�: D���Z?�|\�j�{�������z��	{���i	\X�j�G�Ee�������!���C�3�_4�`�H�F������;�P��$��+�]�F��_	N�b�p�<f�����v�$m���*�W%,��)�p����vux�~��֘3G �	6c�ґ`gD�/�1�k�:��+�1��\��CJ���ī#�/���c|�]D+�����̓*���"���2�#���������BK�X/�DIb�xPtp]{������K��z��W�-u�t0%�pr��"���h/l�W�z̦�o�F�1�֔�9&3�칥�3����t�?���=_{4���E�qZ|͛��x��$����z�f�(jK`%��S�s'�c�7��S�����Jc-��{�Z�ׇ�D}�v	m�SQT�nP�
�(A�C�P��zBք8(�����j� 	l<���{~�����s��� �Y]���n�4��. ]����>p��uTQ���^�"'�{>顯�3rEz�_mBe{JV|�����y@��iRT��Ŗ�+�C����Һ�<.�v���F��C�e�&,��m}K����*���� �q|�%O�z����(iĄZ��bh�3�H�&��?�--z��VQ���yC�D������㧱����nv'\{!��◝�������K�y�s������.��M�U�D��3��`��P*��=�dT���&�[��?VZ�9WtFTO�kz�po.���{�����i�S���W����FAV��ܘ�w���$��yu]+�;A��&����SacD�̽S�{w��^��
)�7�"<�<%�$�Aǌ�:�p��3���w����cDN[^|�W�3�&�T�z)YيG_\$��9VCę���3
9��ǧO�F�4 �	�7c��1�O��m8��Qi��R�-���^��G�9���1�d�-c�xj&>�v�[��C��U,Bج�e8#D�g(�A����vt���ix���eiB����ìp���^dy����_��6E�2�34�9%�"/�ų�H��Z ^���X"��^�G�$�u�F��˾����<�Rk��L��l�'�NO
���^���0O!�]��àa�[/�)�Č`�`>��'�֦l�84�	>!I��d����Ź
��s�21g���7�[ůBš�GMø�+�.zh'���,~یH$����A��rڥ���v��R?W���:�?�m��̙Mb��Ws�l�n��e2����j��(+�ѕ��|�XvslX���.�b�K�H��`h��O{I;g�[$:��B�%?l��7HE�#���T��ЀT��x�,�ժ���v�A�p���Bj���-�a�Ιۈ3vn.+�R���ӽu�� �U�8�����/"��֏�;��*��OH�Z�h1�_0Pݭ���C�)a�S'Xb�t��^�?��+N�|�5�Z�N��&�7��|	�4!#����d ({��c>�"ʲ��+��b��l۝��U�μ+�����]e���v�fΝ!��w[��c�����W������^̒G�Hg��P"�xb?��V��`)�@��z��u�z.��t<$��xt!��^b1+i)���sL��Hbڄl)b# ������1t����Z�
��q<¥�����r+�fϧp�2���8���T��l�`�<��I[�H"#��j���-Y)��W*p~�ё;f�,,>״Gd�ԣ�w��1n؆�'�Hwل`b�]|��n�������u��V7�1���ӿ�`����Q���^���K�� *j���%2�tD8<i�T��9+^x�����S��;|W�ߛA&[��Vh	�.�">�s�^J���;�@p\$�YF��U�{�ݖDr���HBS�*�7��=s5�g/���6ԯ�l��O����
�yg���bj���^ձ���JİI���c�c���mꬱ���̖�Q�΁�r��z�O�i�}� ��d��T�,o����=C�T��k�rb���zE���C����&�m����ID)@ўB����o&���,�V�N��E�Xw�VսR��<�J�V_Uw��*��[�ª$8?�ꇻ2�\ME���ˇj�����֤�7P�-(�ݪ�PY��x�6�đ����"�3�e?T�n5õ�;N��#8�F	�5��3�y��8NW�q� �A�5�ȥ,c��H��<��g4]P��|)(���fZ�L�yPN�d_'�hLb��D>�7��2?���-��oHί�U�����B���`��`�|�+�tq�ן�Ieyh���bH�7�faM/��ŉ��/= ���~߶����#���T��-˲\�v*׀�I5�]�d�`qmEg%N��{�!�]Ixy˵A��
�42���,J�����*E%5��/�_��z�X����N�;��:��d��E�2ખ��^;9����0E��\�9�׿�A��a�>@������s�@��R�lDM���K]'���y���͘���,+�bW�}xQ6���^y��O�PA#H�q�í��%(
�#̢ ���=O�� P�;'�@�����>z\g�q�n-z
�W;���ŝ���J-"o^�pM��ˊ.L5���T�49?/�~�=Rn��^�j��!]� b��[���s�"o���6"p�j��^�C�oXŵ9�҅ې"�Q>�6���1����16��V/P�$������e[��&��DRs{}��j��G�~f��ML������R+���<�ǻ�r���c\�����ۄK��~H8�:=�1��nP�������R1UX 8$��4�Eta+�*�� f�,�g&�ǌR�$Ɇ]�ƫ'"<)�5UR"S����YI��M��xO)�/�)�6�GNJ-R���a����\�iN�!}6�*�����iC��1����.��+���W�W�ӝ6u����f�d-��?Ο�##8�DA�<����<A��Z���F-����-~Y��[��M��TOS[Xo�(�j��g�k��� �ŝ��5kL��L��ob����IM�S]���$�ؚ�nmW�%j��8��=M�k��=�[�.,.�O��r���e�-3�$Y^����O}����gk�e�?�dH�E~��N"Y����'o`e���d�Y��M7�I�Y���7}�����0<{k{:�ԋ(L�$@b�p65B��sM��-���,�xwu�8���Q��c���8��j L��)ni���i����W*�o���(N���P�r��ጊFG8��׽֢,G	U`I``s.az�1;�	�g8�e�Z|���.U�zI���W+�(�-w5L�c�m��ą|ǽ�vhf�OS���v<�y�JT�9�H�w ��d��Õn��-\P�c���^C�^=�X��2}$9ž>���n0{d��9�Q�^�\-�#���fR�XR���ݮ.�y^�H�'�>C����߻z�bzp%��z�����-g�?�S�bzeg�E�����CO��s}cA�y�%<{2в��H?7�%fh��@~,��P��OX��*�j�:�>��SZ���#���OTk�|��������l�l���t�5��]����H���[�}k�\�ï�C��V��=E%G�;T��C��E�G̐�>�-ٚ����@
+bd܌��>��U�csXR��.��<�Bd� �����ABTΣ2mhO��CK�d}�֓��M�>�Ն��E�`��n�i>�m�~�t=?�w�!�u���!�YF@Aa���K�/8���x��hH�E����C-w��p�W������_	|�Ǉ�)<�I�YW��8�VrZ;Y�=�[^�Y���r��y�{|���G�O��V׏+7Ch_��"b�Ս�G��0-�~�b��,[��f�ps�oxު4K)ؠS����Ԕ��C�`���E6�H��̭A�4��I�=��O�c�S�rI/PQ�Ec��X׸�z�ڔ��k��ׯ8+���+s6ם�qE"����0;��(͑��Jq�h`kTE��(b]�b�P�iBHB�,�����+��Q����-�����4[�Y8�����|��Ƨ4� ����Clx��&�9�h#�Ul}�<�_�ͳ���y�+�*Q��h�����<tN�%�'/22||��R��x;�$n�?5S]�=�q���= s[��{T� ѵsi�^�uzX��7m��� ݠg�tc�L2�oKqХ�:�/����V����k��B(�O���4ł&���nY�g��!��!��)F?�V�{���4��ѽ�ZX*w���#�[*o���u�y�y�~+��t�:�JQZ$@ÞhW��i�m�j����L�m|[��,wg�(��yUal�f�D��H}�&˺�ج��d~�jD��9�:��mqZ]nlQا?[*'�%خ�F^xa8�c��󢮊�mAV�ڤB'C��b��	w>T��q3�r��2r�]��x�+m�h;t?_9��
���`'ͭr5�l�/��JQr�m��e�U�K��-�X���W3�#�~o%�Q�7��|����N��:�2�C��]]�F����r�"��[+�IT��}]��I:��.�o���+Z�S��D(/�ǁK��+��n���2���ؾp-g��5��(E�0B�]b����Ez����R�;���I�h�
�A��2?+D#*�R�jZr������Vw������+枍l��˽`8gR>���W�.�&�p�ٖ�O��O!�q����<VJ5#�5�:UJ'��}�S��C�CK|�8E#����t��NkiC��Qv6ϔ���u�$b�x�T��}P�T���|�ȿ�>�l�*O�C`6�GWd��>�
���逭_�G�Hm��6<)�C��̡(�9�a�U�m�����5�A���hKN�q���G����KB�WF��8�����̇QHL����IF�UI�ze���h_�o,�_��͸X�$\�VCc�$֧Xn���w�m���@�B��m@���$N_�w�"W��2R�o���&����`�k��p5����B:�H�l��&�Am�����&�e��g|�7Bo	l��n�����X5��zr���c�d=�}���h<�À�y	�.���I\h�c��`���n	�o��A�aa��?rjȧ��D�MZ+�٩�Yt�u�ʈّ��*)���[�R��-%W���j���A�k��]`S�Xq�.p��e�q�
мQ:}�~��Κ�����7�Ҋ:���ڧ������l��'y�
��$��Ƿ������/�#����^G��T���!��e��߯�2��۱|M$t�X!�u�/1&����hF�%�S,��i�-R��~�[:��G���S"#�0��B��f#�D�A�8�+#�3��3֖_����yWBאW���^�;@����ϥ�aԯ���[��^f?޽1wP=��k��v�m��O����\����Yz&AyG��[�ay��/L�V^�����p�rM�d<WJ����!T��0(ex���#D�ɼ8n�4�q&r:cA]�ʋ�'�u[�v�����x yg�ZI�t#A���L\AV��)��*��Qґzf1�S+Q?2Qr8Iz#P�� �Pe ԓE��7Re"1�9��&I=�B'�9��`��0���[��:~�Zx=/�
3��$�9��f�Y���O��C��e����:���n�����TD/��}��Uf�yg��Y�9g�[px"ph�.8�٨jd�$�7g��yQ�[f��]ÃY��5�^e�/��I��}��?��S�O��̻�A���L U��q�Z;������AËv�N�"�ƅ|Έ4bǲ|��F9[}B�L�6���LH�]����anJC��{%���<��w�1����ڊYLn�sy)�;0����F�5G� �bUu�C
��*2�\�0z�P���s�k<�8���M�!~�2c.$��v�9����3��⌹L�^��~���:%���M�\��b9�����$!�z����� ���Rs��x%08�:��y����f����uf򐀭y��l����?�7�q��ٞ�E
j6n��Cä́f1K�W���_k���8gj�T?�:��eJ�?�������.O�m���}�q�(�X눋����s11�ia��/������vO�� 4pv��rzL2r��Ti�)\}wO,�棶�I ���N
/K�V�Ρ�.��C�)-н�?���(�V��7s�)m����ϲ�H����&Ք.6}��2la^�Q��oI�i�P� �QD���P7��j��k�r]�I��Y7H2�	I��v��l�d=Vܺ�k����0쵈�Qd��y1M}�n�!wxD��W�!�8ȮU���w�Z^T>�jl�bf��*7 &h(�j`��E��=S��;X�������=axJ�^V�B`s�	у��B!oY���OE$��d���q]TM�r�_������-49b��8���j*�r�s��T?&��Q���u��-������e��wL�D_�K��L ���ܽ?�I�)�~VO �|lα"t���nEi����,� �*��F�(r)�X]�:�����qE�v�-3��*��Av�(u����q�+�ϐ��lU�"�ߣj�ꠉ%qUq=l���6���b+��8��g����`s�t\櫓/Vv����]��D�f�G����dh���$��J=2�5�ޕg"''�/.��|K�6XzA�hp��`X���D�|�dIYJ�q�l�
X��Y����9�W�q���'�S�D|��w+��{#:CW����7h���B܃�cqاYa�]��R�I'W0�VYf��h�Ee�¤�p�0��RO��m���<�^YV����^�@��z
��oW��1��"��BWtv�1�]Z�.���B�T����՘�fz��#�P	�D�N��,uV��d��$i*T9�4]�8N����4m�ψE��5�`C!1L�|L����|�e{��ӆp����ڥ������<?��,�1� dgm-�;-S�I^]���L���2�8�]������9�9��#I�����<��V�Pj����Ì����8����^��cq�F���WFҝ���+!���I�^��'Ʋ-n#?o�[���Q�e�_��p���ש���0����sE�u�ݝlr?�Y��f�*��X��խ���C�s����F9Z���/�/Ι���z���E�Ϸ ?E����GH��Ns�I՘��)a�Ff�J�6�+B�Z`�82�Ï�L�mXqs�$�D`@ˤ����_ȊF�H&�79=�ͦm�\?+�E�|Y7ބ�4��h]D��W9[��j_��$�G����d���2Yh�`�e��2lr$9]S�"~k��M�[�8��`Wz�����VP�۾����I!�ŗ��i?�&�Uu��ߪ�a��o�a+�uT�=%1�ڗ��Bj���������C������
*����EK����5��5�@'+b���h4�ۙ\��FԼ;������^�^�U��n q�ٻ�y?���6��I�����\c����F����$7�����(u F���q���J֕'uLBN�/�)�>�0�ɱ*��/�_ ��/ڑ�q����|I5OZ��*m�AS=�
���G��g�GH�S6�ʴ�dpWs\S\����s�Ҷ��F�Vb��k�յV��{	�49�2i=;J���~��ÿL��A��9�&g#R�q|'�/�6r��^�Vc����Y�ʥ1�5�Qr�Ӱ��͊+���d%��F�����r��n�ےqb+/�4���Ƚ�D#b���Y��Tճ]2G�*���M*X'�&��l+<1)pK~���]wV���C�5�T�!//�C���K�,T����(�:G��6�^/�f;p�3N�gu�^��a6Ӥ�>���>zX��"��-.�	g4�gv�xL<�j������� �o\��T s�����f�gٲg�"B�I)ʧ:�lw8۶qз�T�I��s2�T㳇����x�~�b��at������_��R��.�^��3n������ԋ�MT �'5a>`�2�Q�w��%����4�}�.nb1��7��vن�Z�G�q���^'XYġq�����Y3Z3,��eW��w2(T��6���	�J�k�K� L�/��_)� �@s�iw�����u2w�\����x���bwڻ��5�;jme��)_F��;u��++�T4n�h@�j�ߏw��S���P��MME������R�m����Mܒ�c�Նk�N*ujj=4�@)W�G�Sc:��<�����o��#qm��j]��R�bG&{G�6�Kuk@jS�k=AS2N�wH��d�^ͻ��kL�A��<��6�-_%���ǇW����ےwv�<��d+��N|K�SW�2	K��rO�=�{�T��#��s�Q�n��iUB�$8��Ψ�ݝ,wz�H|F�T/3��Sq�"и˗\�xxp�Z�J��W�(�̼j�
t��T��F����F��I1�̙ aw����#4���ϊ�m؎�R'�ʇK׺J���,�=���y�`���j�3�^G?K��[+D�\���%-���9s��H����slx�\.J�-�A�H���}*��p�Z=-m�Z�a����qZ��e��\؁�N��d�T�����Sm��慢7��H��y���c��[�Ե�.�r:��D�彍�oI�4H}�p	U���?�L��%
�4�MB6������obX^�lp;��A�8F���+U�N������\Ny.�	�����$9Ќ��$�M]INgJ��b���xC��Rs�bm���1GJ�G��w�H�R��I�eCR˽�N,Ճ:��br@2��\�Д�k����.��	�Џ>��|��(P@��-y��8��\��㥐X�4;$���N���	C=�Jd|��ы��X��'O��~�Y���_�,�L�s�����Hd~�:��BX��{rA{����j2�+4��N�O�]l��#�0?�z�u0���9�����~��-�@=�g8��zEi;V� ����HV'ԗf9��
1�k;P�	�n��\�U��jj�XF%ì?���l��������r1��N<��6!�H/c&ܷO�Rᣰ�+_, ������}���	2M�W�c��
�hޥ� T�CR����R�HV��A��(u��� e��7򒺙w���޳w�����p��HJ���%�R�Iц���O��U�P]�x[�d����p�E�m�v��nT��6��m��D�ܐ��j�wǛ_�x�an����3�\I�TNˡJff��&ʼ�y�Ă��^B$c�$���D9�I�܂�SRMIg����ʞ�|�4^��W�Iؒ=�+J�(��(2�&`]�C������A�-��];�S������DaW����#��b*�v3@Z)�/=��\D��+mI���g~Y{! ~�����wϼ5�LE� 5"�%�4�C��0����I[���9�\�����
��qݏoҴ,�s�)w<��P\�)"E�xb�D[�'5PB˲YR����Vy2YM`Ja�t_�L.�S����T��t�����M�=����JHL+J�euH��]�e)yCG}�L�
�<����ٳ�s����lh˧���_C$������
�r�O�Gf"[��$ơ�W�X�K�����eg��$ x��� h��`߫K��{���ٞ]7]�:�J�����~�L��~_����gr�U�s�=F�i%�s�k�Vq��S�B��m�����!���/*�3�+�x�f*?�ܟ~�ѓɯ��7��t�uUX��5��Ɍ�8u 	�O�z3h	���U�ةHA����������T�pm:-|c|n'w�[��Pڪ%뺲��1wo�&��8{�툐u׮=矖Oõ�s����V�y�%L��eCL_=����%���HLw���7��݆�d������b:���EK���J�X��7A�v���]H��g��eD84����wi��5t\�+�`	���c��a�G�&k������3� �4���0)ҧ׸�A:�y\��1?��ʋ�A�c ��+�}��{�ܱX������"N�N;���k3}/S��Ħ��l�|(�xC��m�^�+W��UG�����HO4��'p�ax�K}Mn�}	e+!C:��ba�T����~���d,��X�u[��5
�/Z��hs.���0�-@R��	n�JP�;��?'�s�oOM~'I����[���2�W˴��-��Q���14b���1	�RI�g�o|�c����]�8�>g��<MAr`�u�f]�j��'�WG���^�-��0����3�"[�ưbu;�q�	��w�٣0�t��ȭ�	�n,�i~���֢����Vq�#,s$�A^Bur�(M���BSH''�C9SF���CIZx߰e�Wu  u%G��HG���~�le(U�;����Ǻ��8vf)�Xj�4ǾK�a��,����+��A�=��Og��B>tَB7D/�8���Wj��$[����b�;����2��t���������N�7����A:���ZGlC��}��LYv�s��R���h[�6�5�'��liL��q��S.�Ub^zG��������'e�ļѸ�c�r�>|�Z(��78��N���7E�s�j-�YU���ہ������3z]�T.�W!�3�T43�
bU���B*���@���bK��C�8�9�A�w/�.� 흒mo����C�xm�2�g�}��rA������~�� �&j�qǷ�,]�%�Ԯ�R}�"ɖ!J�`L)�׀t	�4@f�zD?�j�-�*Ir�)sA��2��
,���n'�Zl^"9�W� zTE
n��祹[����t�=m;��ߦ�GM�8G�ӆ�)����d�ɂJV��%�<��(��.��p��Ւ�X��ҤO��o���,t��m�OJ_����"���&�Hf��$.U���h�y����z�)l?���G�$��P��d���̟��6ԛ�4q�ۢ?�E��Iqo��b�,��0�e8�u�̜���X�g��9����RZ?-9�O�(��z��g��V���sɪ���q���u����y�Ϗ�|{�rsDa2���P�r�2�y��ق��@գ���Ӏ?\������8���������_�&�nX�;?�
�����b�a�BK�B�GU9�:�L[��٧���i=��+����}�T��#"�iy5�;D�#PJ=~�St���q�[d!��cӒx<�<�6/��.rVRj��_wTY����f���1Bz�BVxh�ޠ���VL�D�c�5�� x}B&M�1�z�M��<��ˮ�A�X�@��_������1fg~rNZ�_��t?!��$a�Ce6��2^�2H�2"���^������<t�u({�i�t����`�|�Cʹj:U��1���bEl���>�<��{j�_UW(`�� 7L��*ǁAǊ;0 �����#�����'��˸xA(vC���m�VD�2��i�q�MC��;Nv��d��LTnA���f�ӱ�?�������s���kz�&�S��b36 ӐQ���,R��Tb���]�9���\v�'5і�R}&���Tm��1j�"
t����t_�Og	�9O.궙���#�3�?�l/�Uo�_2lZ�q�P�i��0!w_n�x��c4�����2��Eh�]Q�"2=�{��u��ۗ�{6X��x��á�9��Sd.^�r	W]R�m�F+b����ȣb�aiE��sDw*k��ֆ�G���A�z�e{���I#z�(����W�g-�d�؆��:Xu�C��%���V�
�UJ��Q�싩�.+��(2��*��Io�YI̓�P��L��'w�s<�:���6.��f2���ղƫ��?}�� }�I���Q��#��(��@jDJ��V��S�l��A���q�b����m�ť��ѓH�[յw�( $8�<�CZ�
8khO�r:t�Fk�JoT;�t�j�m�B����C��r��-�w�C�Nf�o��[e��`��	k��=n/��/<���8�4)���5���eQ��:{W)�4sh�f*�	�7�"��!%�T�E���{�v+�N�|dR4i��c�M�]e��k6�q��/P?!�Y<\�|>�]���U.Q[�pH�$�l�1�U`�}���L�K̸��c�W��������gi
@� 3>ġ���0K���a��Ov狔"�v�X5����'��5����,��yXQ+�
%[x��$[Z��:��Fl��0d�e�t��)� ÿ�v��~7a=��׾��̟�
j�g�s*� �z>�y(�D�'��2�4mkG3b��A�"O1�d��'-�s�����-����,pkT�tm9���B	%�`F�U�'����/��z�'���g���$Y���on��^�I3CI��z�����L� �׎>����a��_sV�d��r!�K�՚��z����u�Lc�k�5ZdS�y6넴c&F�̱oL0����x�l�r�d���CSv���@�⹮@���L3���΄<s4un�%��:ݘ��q��_W����D����t��Gi��)Z�Zɶ�n�'���XM�N��	9-���?T-u�)K��w�3"N��h��e����O����ݗ����pKJ�-�8Z���:��P7/��@�jWoˡa����~�v�\z�ךI��A�(�Xͧtߝ���UZ+77Θ�JG����y�� x��zZ
���?�����U;M�cb�H9���F,�r�z�,�k1}5W�
r��"tdm��:qDBޱY^��.}�7���� ������d8�'����H�.ww
W0D�T2i�|Ժ����\ڋ�.���6a�fTg�����J��*�9�I��ݾ1戢�-���A�A��T����K8�r�����*�y����R��W��Qw��Tڣ�e90�x�t�?�u��K�O<��Q�������Hg�J,�9��v�# �N�'�5��/d�L03�}�Dx.�b��Ղ���G��LuF���I3�Q�،�7Z$*���6l#g�3�Z�o��MQ�|��G�R�y\�v���^������P셂��ޟ�E����Pw"�&�)1"r���i��
�Ձv3�K�����r�;�%���R���&]��)?T�%��yx�l4���x��{�����\Ci���d�D���AV-�D
٣���kx[J����+m.�(�� S����y��f5��3MWc��ι�a�^�;K���,���7,�����,X����԰C+�����iwE �s���i�{�J_�W�˲�!�,)��l,�.���R�����F��\h�W1~��?�x'�M�9�Dm���:9�����$PR�?U���b�����җ��1�L7�ܞ:�j�A�dRk��tO�f#hi-I1�UE+�n��?͍3�2���m�j��ۢ,�_(��H�$�|4)��2�I`_x`�Z�8�tY3@O�_e��������8�_���$��������%���Q��
|_z�{�`%ƱƋ���/T��� ����2��9%����+�$�X���~j��R�7c|l�O?���?ɱ1vw�����tX,��kCTc63Gr7z"6D�|�oq�8Z�S�BEaw����ca�x1E�4�y�c[d�<Zs��Zg���m�5=q��i�Q������OC��U����r\J���q�m������-�a��u> WL;����lrN���&��5�dm���65�&��k��"��Aѧڎ������=���OQb<U2�P��=��'n�rhXL`���
8͍)5���9&��bZāL'��Jр�i�hL
�O�>�����&_�+�����ܒ`�����=�"Y~E
��U.Lb���˒�����aq�?m��r�AxЫʅ�ͻ+m!nt����	q���y
���H^��=�byz����@�fj[�G�{��j��*{�x�u�O�-ބQc�	7�o��VڥOV��^��z^Ӗh�:��'��J��b�O���K�78��?]������-���n-�k��p5X�"��D� ��Bt�wzv9͎<$}~�U�R>ꆶ�S�`y)(��$p8=r�1�|���7�/�=7�o�&q�\'���C�P;�}ѩA��ڎ�D�n��!l ���ߖ��Q��eTWis0M�SJ+�p�*d���,�z����r��YU�PZ'5�������H�w5i���z�ᗟg�-��0�嶋0��;0�1�u��xC��^���8�.-9�Y���n]=��=��ͫ@V5>~�X93//�zLg�WIIb�[�н��-v+�s��s�POYڂ���y�qT���;�K8���wp.�şUO���[Kc�
y<�;� O�����S���6Lݚ��;�.�}o�(�X��(��<�\L@ӂ���YŁ詛+�^m�F%� ���2�Pv\�e�A�y���9��FRR���T��!s�q����d��8��mM�6]�2����r�F�j�d`����J�䅟%����\���lQr��|�j�� ��#���wJ��A���S�i\!2�g����g��H�5��h٘I�e���,��].HW-� ޔn�_��\��Dt��a�%�(`
��(�'��Ӵyk���<v�-�cU�}�d��a4�p�_Tf0!����	w�65%��3��J�!6���:������VP7��$�-}cr�2�vM�ve�'ݰ��-����^��d�v+1�n�;!�.<��O9���s���x����� �B,�r@�mS���J}X�ظ�#�~Nv�I��h��oi�eUFS�t�4+~�ם�VR��%�]��<�&JKH���!��d ���p��F�a��c���x(�ᴡS6�̃����(�B�y��<�?Z-s� /�q1yr1���
�LSR�ӡs�Y�ҡDP�~o�ڕP��U\}��gr"����Q���_;��,�7#W�n�l�)����0��uL&���8���JA�u��)�Ȕ�$�˧<�aPi���iZsv2��
,�8�/��ysظ]k�gF��~��ó��υ�Gċ����v��CsA�q	:�5��%�$��7�)�2�C�o0!��&U�Q69w���C 0��VQ$�ރ#(]Z�����S��>���V�����A�%k:�1[��97G�)������?�-!}��Q�K�<�*OVI1>�&�E2��V��P,/ڽ��\h�'� C#6�o�n��?ι��M�@I��S]4���肀P�#�G������v�`����;�~����~)�R���塰�:�&�<�Ռ���"����O�p֟���tv���/�b2�ϛw\5�������r'Ǻ�2�&��4M� �[y	�H$ŋ.������_����]��̔t�?�� GzAR�{��')��I��&P��I9q��}�)�?m���zjA0�P.т.���V�D{�$�)�;��'�/����-�J4��o&w�L�k�--�3ȉ0Xꍍ������SOD�g�v��A��+�[Ϟa2p7h1n�,��U,�x���)�C��'@��jW_tl3��9��z+��L7@p��ɤܥ���5�P�2p���f�)Dm�@��ŋ{�#�GG��br^�Q3���9g u�x��i-��C�/V�f� 2�݅�[�ue܂��-�G.ir烁2&l�/8EF��=���w�fI�)���
�xlv���1'�Ƥ
$�JM��\B
��̛�����X"[����L����
�;2l7�� �U�[̒(S��hzD�B��<5�J�8C�H���;cE�0�UY�7�Xb�"�K�����:j��&`3.ܜ�~w� ��X����_=�DW�W?�p#����w�h������2�<�3G�#��c�B���~l@�2t��J{�Է����9x�W�/��g:)9OH�^�[��݈ RN�ޅ�y惽��׮Z�pW��
ueqL_��e�ݍ �_5z'�&j�N�`�LD�^����^=
�دP�ߏ]�+�lˡh�m��%��v�sb]N�װXmD��e��Lҷ�C���|�aD3M�l�v�i>Sȁ�7(Q�eNr���u�d��4�?�:ax���| �c� 5�u.]��T̽��>n ���Ɂ��
Cg�9Ag�e����gG���'�K/ގAo�@H���?������q�oM���v�n)�q�ʴ1U���LX�%�?t����\��sG�����<IK�z���2�T��$��̲��kt��,-�R��V[���Z�_��9j��w $�qrd����}'J� �w�|*2v��x�����<Gk�$3��8HgP�Pz����^����YF�yɀT�������`3F
�����3�:Hw�'���Y�5�{.Y�v&l��%U?s�%+��`�2ѷ�����m����]�o�=2�5	߶5?�'j�ڋl)�<�a��ńVx�V�b��3V���ͯ��W��7���.�=E4,	�TO�ba]�m��Sn٧���&�����8sp����n��N��]�!,(Y:�h�D�3�'�2����O��/�:<��˘F������E�d{8L{*%�f�B ��{����.�"w�G�넚�P�z��h�+�Р�OWl�X��s50
_�(�����*�gR��DA��lz�Vl0�K�j��ֽ7Z���7F	i-n��N*���C%[Ny"��?�.��D�@c1���pC��G��*�u;5jܳ��D���=��|[���w�gt%� ��t�yc�~�_�e���A�(mUjp?$T~���M�V�}U����qc�#c����).J�ƙ'��-��RfZ�*��A��Qj�Ee)p?qj�����<h���������tH�QU�;�K2�✾aQ��N�}�ba�A�e�yi�D�S�0�+SS򲮋���ۤ�)O�'��}�1�%1��!$5�N��4�5��w72)i0W#�D.��5�![�0~�	�`w�/%��]G�3�u��165L)���EƉ��G�B��p!�������˫�͓�>9_"�AZ�U�j�=�
Pk�e�N���y#�#<zK?������p;�Z��|��3a8Dl԰_[b�A����ؖ$mym��u�u�����m��L�Y�����|�($x�_}t#���0���j�������P6�,'�8��[t��_�܀���Y���d�,�=�����ˌ�֏eW[�{2ĕf|H��Id�2��%%^��UZ�b�2�ؽ��m�[�<���� �9T�Z��8�S�<F�p��Vb���U����Y��O��b�h�'j[���"K���x&|����oբ����^���;�`ˤ�����f��" ^��Ȋ%���F*��r�t���W������&��]Sο��	�W��//6m���D���:���4�jwn*%����Cj��w�1�~��$)�ikr������⪎�j�ۓs�9Arﰋ�u��E�o��E��	��
�T�f2v��>�'<t�T�G��}�sR��@i͉����jJD�+��0�$9��5�q�0_B�`��+�QW�-�`o���Z��V���%5�9fb���Q�.���ْI��	~*�2�a7���o�����u�n�%�c-kah ��y苧b�65h�2+��v�=f+�<�/��X�H��i�ˊg�&���`���wq�Q�/�`�C=0��h$�Jv_(l-l�!e����~=�_�A��juq
K8�ķ�*��-�&P�SR[��w�q;��#}*��~���cc �0Z�2O�]d*�%D҈�Z嶅ʎ����D�#yG0�8e#�]<9���T�L�1fA�u'C�.5,R,x�.ωN�Ar*�s���$�XT�v�C*ݤ+���ǰ�,�u�9/-&��ü5�@w
��]f���*E�D<Z�/���r�"�T���K��yw���;k6��N��P(J'�jJ�|3���q��y��2��uSx;�~.Q{�5�>��c�*������p|L�.@�+;�CC���M�>�֋% 5ю����<}�|D�Մ�����г��gDڬaN��A���[�ʮ5�Il
��9����9=��j_jd�͝ �A��3�F��	ű�N&���s�p%����]1�ۗ:SȋxJ^ ���ta[��c��ϓ}V	��=h��>������t��~�E<d}��t-tBKd��{�'�+.�PN4}/�����b�%5�Q@¤����-a�BIb�3Q�%Z��@Aܱ��I`ŵ`���_�#CPƙ���o�U��/}�Itӛ�D"�~�eL��o���S2�ym��� {�`Ƕ:	��/�Z�1 �ʪs@u�-R^���<��Rd�d�S�~~��@OS�Ӣ��J$��I\n�wђ���J�pӵ!�g5��)$��Z)����:�K8d�F�o��� lhd����Or�~�M���	�bӴCdy��n���M;�%�̓��fշ1�p���0+{�U��h�P8wh$��u^5" ���讛��Fy*Q{��H�u�R���sQ�_�e���b�-g[�d�Q!DK�e�fSK�~��^�6ڂ�Y��Ȯ��ux�q�Ӫ�p�S�o�`MIg��8��^�'��ߤ Q$�s(�_���o�^�	jdG��b�g	���?y���Q�N�ā](?S��@�W��A��x�MJ���Nm���[ &��觳.��b��>0awh��L���%�5�ۋ�n�'���=�)t(��\����������^70�����t�y��+� Kh�ʻ�st��;$X/�e	�以��l���p�ݼ{�zm�r�O�Q$/��`
u�
��I�T�v\p<�Z#�!�-5Dj{���;싽xBդ����[Bj1h�q羉'^}�7�/���t��z�g
�:���q�O0�)�L�ǩ
�8��\��~��J�<��߷�O�SqE!�|ɮB��qt�:{b�C�|"��ȝ(~*S�nO��?R����`�o}V�b;��`�p��O�����1��.��ph��\F�|x��|JU���m&}3�9�7��-0$��dZ� >bb�{��$��}N�iA+ �W�pJB�Q�]CZ��u�8����d4����oM�4��Mk�ϔXU-�®�2܇/�>��L�W����>��I�4˨U�t�^u��n���[��N��j/�ӯ>K��Э�]��{��\�h=~�Db��3Yܹ��6CM��VX����M���%o�Fft�i��a�:�l��ﱣ�a��gM�V��*�"�N%tP�7���\w(��P&���-ä�R�'�1y�������=ץ��
�q&��Nn�yI���+�2M�yk�kq�"���[�nZ�g���+��(��`Rǃ�R�����kKX�L�<3�S��Z��>���jU�(���VU�T�;Rb�P�;j����&��)c����+��+���g��0�p�U< ���Q�s�H�Q#�ղ$>��P Vb
Ԕ�g�WwT���u>����0�e��%�Ǳ�:غ��&,���(�����ԧ������E�a�5F$�i�����|,%��!�P{:��6N���7&j̕'LM�Y��a���ԥ�����?Ck�
@W�3��Ɗ+�և1^�xe�\���Z������<�Bg$�x�}&�
;��W��V�}�((�A�Nc��'����cvA�!��ҳ���q��ZW]�1�tr������.���'�iUk�oTi�/��fy�,.���S>�6ݷ�|{��"s��׆W�a;��OaJ?3���qj�� M�sy�m�!ҥ�z؀ג��P��:h�3�&�]}b���I�����	/p@�Qd%n���`^m��7�gN���|��1}��(��}����zb.��N	c?�1����	�q4�zZ؏��Gd�mԏ�r5�}hq	�LR+jƒ��R�m��Э�����a&��j�/�9%�!6��^�V�V�|{��=���3�xl�67�kv)��$Mk?�
Z;j����JNf�W͌�B������PSLA�3��(�� �����=�"�c!��K
<W	 �hY�%"�!�w�����T��Y�L|n�H&��^��q.Q�9|�&F���ǩ�Vp���1,��ɟ��ܶ��|��s�pD��@��Oϗ	#V��I�rs�\h�j�&��H���~§����)��
{ԙY��.�}� ��$
U�/%*&����ѥˠ'��C�o.���IV�v���﫾�"0��F�P�3-��߫�ܖ���G�}����i��]��}�;E!h�U�V�1.!z��b�G��~eX2�_��N��S����m��Rm�o�s��w��:x�N�&���f�GW4��n�s�B��՗C����#չ��"�2��6�E�8�Yn��F2\���E��DdoyS���8�Q�3k���G���P�(p�6ߐ�����=A�3�w4��X+����F0�3�ø	��ڬ�؛�\���n���tU�jG�8���Τ�P���ǀ�f(<���	/(��u�Nw;�-�x~�
��g��x�%sQ����މ�V�Izl��C+S~j����/5�Ĭ8�}%��
	M���\�`�p���Dlr�x��DSm���o����ڥɁ��v�	$��=m��$Z)*4��T(�Juw{T���0�	x-@hi�0B�r�M�M���R�/ wEx�sޢ��F�vY�1��CS g`+�߆��6�Ҷ��v~%�23�LjP�b0f�������2pJ��<W�u�;��e틘��u�Za8Q�_õ���G���k�S_0�5���i��������%
��BE�^2h�?`���9N=*�i��_�oAߺ�[lrU@]���.J)+�8X��=��c%h]L�ţ�*��;'����3��_{��%3�c�>���ĺ�I'�lZ<�>UM����yշ2���B�*S_�M2�6uU�nu�y���qF�B6��.�R�οZN �b	�	������|�F��9�7a
��Eؗ��x��ꀘS�k#�V��/Rd*n��g`P��P�y�6N�@ �[���R塰������jZ�:qn?��;N�Fw���ziu~:���땚x'����/��`e��q�ZC9���rQ&5�H�1�-���!�VS��$��&vX�wnJ,�!�Z�A_����h<�^7U&�&ii��	jg��"�ę�S� �LK���>�`�.�a��Rv0A� �gq6|,�7��:zd��_řv��xY^���V�Dؔ7��b�^
6�o���J:)N� 	U����/h�JH+k����p��S`!����P	���|�e�Okv��>����I����r�n���4��G`�ߋl2�m|�ڧ�$�q��q�Q�����PRؠ��H#}�n���94�^`���,>���S̱<�D��͒�4�M��x���S� ���a��.o�1���4����3N��rˢև]'�\_)�⼛���ި�re�z��~��tZ�a����a���ڝȊШI����Y}�~/O�&�n�M�2{�������}Y {V�sLC&x���ö́R�i<�v)��c��|F|n��û�퓭�'�09ӪH�I6>l���	�~Ng��!�3OPȔ�����U�g�f� H bg8O�P6N���׎>vFg�7�̜��@�y����Ҩ
�]{_E��md*��1�*���3%�����d¼���О�$�Vl��@�&���ڜ�!i�i�_��[�/Q�
U���!Kʻ�R��!}��玆��	p���K��`N�������}�jw�����_GQWH;���lHO8�R%X�f�'�Kc��Vb�f�{�s1)� �o�����&�G��Ұ�k�����������_����Sn��@���Pǌ���2rN%Q�E�lFĖ
�zr�)Z�[=w{��w��f�a�ˢ.N�9��C�����-�9hot��y�
 �>��� ��v�0mAV�/e'�M��q	دE�b�F�B՚�:,kʁ������g�3�|0u1�^�5�����]�cL�Wb�c@dOɍl�����x/�+Fߠ��\DP1BW��j���������/������)_R���μ�K�d���7��"?ØY�u	��� =~X!�kџ�/&�
Z;��f|\pSACA^��W�]ʔc(�YP��ذf���jB��x�b�)�%��2I0���1M�s��xg�<����V��s�Y���Z��G/#�!J?���Vͼ��8U`auE���V]O{��B�R�x,��Ābf����<E$�<��R���\���Z��\_��B��	=���kv�-�ǟ�z�R{/��j�g��]
��8��C�ґ���~g�LY�o��td��6-@���4x�xOSV=#�
�%�x�
��̴�.sDf%�x~Y����}�E���t1:�(�^���(<2�$���E�̥��G�@�2I�� �S0q~����oZ��C���;�:�Hml �$��f|쀕�w��k��'��h���*����^^�괟s��}gEaV������c���6J�����,Ҝ�"�T#���v�kƷgH���F��$��3�x�I���Y�_���Y��O�c�R�>�}`��$�4�������P���n(��~�%�.��$hU�� �0��
P�g(��O�?�Y\9\����S5;�zh�����
�cX��������U��-���w��Exa�.�`5�u!-�wа0�$e�I(�b�a=��M�T?���:�`K��e��H	hɖ��W�<Ч`Ъ�����c�B�Jm����I� �ٚ6�;��0�� 3� �^ �v�Piڇ��7�M�F�F�=��K[�b-ŀ$a��\�p�.�wZ^Pʌ�eS�#l�
�$^�7���g��Bq�O.�	Ncl|ث���Fq}�R���A��+��E�:�NЮf����$q��hx���`�tB1ݽ0r�����dV@nP��ݥ"����]�-���<����/��T��K��}�(��"S�~N �K��"!T>ˤ@_��w��0�+<vwu�Y���YF!��lF���cJ?&�C�f׋���&�n;
2�7~�Q���iנR���Z�UU<[ׅ�ګ���t=�OЄC��T,�-ye7(�!;{" M�8F�ME�c=J���H���ȍ:�������I���<nψ�9���[��,ٞ�(_�V���@B���t�"`cqT$�"��$�	\��o����y�lg�5�o��݉
����m���^O�	+�,�k�I� ѡt?Y�&g4�)>��#ݶ6κ�~>e�N���G����GA90��O�z���uR�3V�.<��P���ӶXd����IuזWԤ��M�M�K�'���0~���*^���{�,��莀�􈿑��r��7KO�j&0����+��#�n�4�FeC3����|�ӱP����#�*|�߈�Y�|>袝�0�d�Q���w3�= ���V�SP�Gl	����A{��N��o����o'^�˒c ��v�X��:��}�iUN�1�uru쉅&�'}�c��f\ )�
t�_���?��Y5�T¾׫r�Y菧���S��w�Tt�N@
��y!��Ҍ�]��qU�R%��p���?m�ezc������Tԝ���?<����K���|�eO�=�8���l6��P�x�?�a�tR����3�Ԡ:�����t��N1K�&Z/9·�g��B?ޞ3P!>��9���́c���Q�Gp[�u��؄��k
�I����KDkx���8�I}n�pd�HQ9��z+�=��t�S����hR��^(T����%�#4��G�Y��7������B�����\pro�����wH�2d��»�G�[k�%�N�^Mu�I����]{'���FŰf�>Kx��p �[l��}��-O1!�^�|_r��u�"/x�b��si�G{�Յs��E���`�u��bQ9ɷas��l6Ί+]��u0�l�K���~'L���J1��zr ���>�����L�*�!�?[�ڊo'^Y�w��Nr�������@��ŀ�����-��|�5��VmV�t�������1��g:�-)b�Q,0"�C���[��+8�~	�J���[޷�b���#��1����� �z=�dy�$�v 8<�C�+���@�h,�*�HU	V*�g�b��Ley�<�K��N��b�ϟM�ڭ��Ġ*��÷��_'���ؚ���;�!�n��M��Q�69����P��}�3�ه(c�![�t�f�e3��A�����	�bM�5=���f�����G�xh�J�$���������	{��& L�=��܄iĄ�f�
��@3�v[}�\.=�҃Ճ �?�"t�����R�42�_SW��U�G��3����E��/���+��׎-x��¹mSr/m�%6����~}��*�J-mGn~�	#�����`�V��3��o�!��z�r���Ы(E�R�@�$}{�hx 	��a7*̟�XJ<?��/w�o���Mɴ�q'������Ӓ^A�ۙ�37I'�-�����<|db#���lYw"m��tziS5�o9�.�����N�o\ ��p��Q`0N��z�~ye�.�C	["Ϭ�;4q�>�����y�B�*�m��c���l�H�E�|�����_ �O�k<�'�X��]`~�fK�t��i��������Ǜc�Ew����J~2I��˯-q�ޭ�4�Vk=�:���������cuL�h	z�&aS\M�%4�YB%?,�r*����>ޤ�*NG@	|N�6�eZwWd�-�v$����>�Ka�"C���gW)YS�UIĪ\���Ҡ�U��/�O��q8-���A��q�r&��̝U�aQL(J�h?p3���Nvv���P"�u�]<Pu�K��}mQ-�������Q�;�6yp',t�9�K���F��rG,��?��]��ԭ����o�h ���������N�f�I/�?��"�5���Z=����Tog�[]�c�4�\����|�8�W���Ja�O��~��)��jBpýD�n�hiĄ���D�8�u��U�JG�qM`2z��$7�Ff���:��w��L����G���'գ3������C[8<*�N��a����׷��}7�:ڼs�X���ɹʩ�C�-�a���f�s��a�����.��20/��+^97�C�`����O^`D�h�Pt����;���@
ޓ�P�AX�C�n�3��]�F�Qy���7>��tݠYo�����"�`�xiD���g�i���~�F�tRSN<sW}��GG;2ݸu�{J�F1����69��G�}��8B���W:^d�l���������a�	�%w�\~4����r��T���4/$���T����*���h+]�AyY�㤥�7�{��R�Q���׷����Î�8�����p���kNY%�+Ic�`�����o?\��2�!�.M>3���UU�{�9~��C��%$�cSV,உ�d���9����$�ço9������!o��0�
�2X��9��l�����Z�H�.���dϭ��~&H�W�[�|N�d����\'x�lIȦ��%��+m�0%�2O�����'ҡv���́7�Tza��&5��o�=+ �g9�,6C���!qY�9A��o�O|�EaB q7ذ�xe��h���!k`�|�̊�ruxҹ��AL�n���=.��vO��31W��-l�D,m<
��'����/V�+����� ~9�$�bW�4����@[����w��ر��n��S�ƚ�L����	V�_
x�	��\��U���΅����8�{�9�	����T�?G<�����b�[44�'SQ��X��RR��r@|*�J��<��Y��n��W_�cR�2�2�-�է�v�ں�aH_āk�%���,�2qa���Ö�M���Ç��|����`^@�ߙ��j��Ek�8t�t��q2�nW=/�4�3�1.T %��+
L2�?xc^���	��Ra�+�e��ȗ���H&r�&���G�%j�n�� }wj�]�}R[d~N���'>,o_���]��[��A3��3��	�� Y.n�]�1����q봯6��(��C��CJ�}����t�|�i�sZT�d�ar��y'�yr9x{�OĔ��/V����b/�m!��?����uxW�>	_DۓA/��B[,� r��'g�ҕ��m�̣�@ٽ %���D̲�ѿ�,&�*��W�\BL���Y��c�ȭ�� >�:a�����+r��GwfN큅��V��w��(�N����^@׆�?w�S�<��[s�\1:1@�ͱ�-�2�m"�/���l���/8��KMpTuX����	*&w�|�ݨ�d��ľ��
���o�,��SW�㩺�	N�v�����)OkO�|��g�3��������+�PhY�Ea�� ���}�s(���.��q�_��8հ!����l��!�O=89�]�Y�����(=!ڰ��ɬ֕'�L������O�͛�d�����e��C#�`��"?#���}7��z�\�\�f��$
7�66�`x�T��A��t����v����N$�8JAVm8�˂�Ȳ f��ց��z��f/m�vR�
�*)kB����^@�\���[�p��I��\$�y�[���,�/p���LP�)�{l�.�$�(�����<\��Z��ܐ4q���Oi�c9�+V�?"�@E�hOQ_�$ <b֢hu�}Ԥ����O�k���i���Z��:~�DǍ7n%�u5l]����%�	��\�'W^0�R5I&tI����½���'?�8?C(#�吪\'�Yk>y6FC���&�gD~Ҭ�]��������
����ԟ���1���.$~�_����>P�ϥt��I�>����Z���f�mC�B�H8���T<��2K�ԫ�l����x���)���@l*��bhbӍ�vZ����f[��.���,e������lO�P��7��%]IJv��%#�$��ѧ:�W� KEW�7 �� >�X�L����[`蟵 � �`W���%�d��26
�����M�VK��q�Fe��#���+�ӶQ�0�E�4��_��LC��]�� tw�z�޸m-��'t5�IX�%�Xw]���1[ ��Gy��������\1L?g���ml���&�J�a���WL��wQ��<�k �a�Ѓ5�ɫ����f���ë\&e�|`����©U�>��"�60��"��S�Um���<�n�w�_m��n��(q���E�g��dueL�J���Z���~?�.[vh�fP�)C7����V�� ��*s	B��O�n��AͶ��q˹��a�k0;K^���Y���N��`�\"����y�����R�)�1��djl�����`cr�y�p�`l�?7�0�\�C�e�_����\0�,��:,�32r-���3�����vjɓ���	�Ū�O:�K��W�D��z�4^�R�P�XS��;�_&ꮳ��',�T8�b��4]���y'�4��%b�˿q��2x�t�e�;���Q����� ��$jmb��2���X�d�Ik�8�2&�mtI���_f���\>��xT�� �������V�Q�#iyr������[H G���(|�[����K��W9��A��IW}G�+봎m�c��Zzf4�1��
��M�Ɨ��K��� "�LZ��x����^��%Ua��I���H��W�'m7;P՚Y����F_!���;���I�!7�,A]��������s����*���鮁t�J�\�Z������x�[/����ZX�t��8�I{Ǯ/V��h���9Q]���9w�ةc7A���'�R����H�<&FG���j�S8�C�6mA�����E,�"��Q�'zʂ���#[������;�%��u#r4*J��^��l��(yۋ;�u�)���g��������Yy��Ep�J}Mu�k��l�{$��U���T�qH)Ƚ)֐MȒu�:0:8�^�?4� =`�f7&2��Rt�-I�2��(՛�Ҹb�42c�hC��.'h��b�؅%��HĻXH�'i�K��?���R�?���|�i&4Kť"N�"޺m%�A���>�I�/��e߼�V��E�$�A�N�o�y�9]��%Y]z^�<�}�Bo)K�P+qR���Ό�>4�5=T�kE(]�\"���&ݎJp��f;h� �����ӧ�&*��D �y�`+���c����d��ҳ��#b��UK֥Ƨ�]���O���q����A�5�Wx��{ǿ��4g�H�j��1!����NN���M# �T]�3�KS�(�.�$�2ӟx��%e�'�W�u<�	y���Y�8�|mR����=�E�����B�Y�"�f��f!�h����$t�B����0C����oeP!ن^[��wD�����=�� � �FqvcT�\�@Y�Y/��m�����|���f�-�&>;�.�&ͭ�f:QOzeB��Y�<��Q�HP]�8	�c�l&3|�A�j����؈yJX]B+X���{β{��\&�
>�~�Yw�1'v����/	�`�:�2�������ڿ�o��K�1y�z�v�}M0�FAz����A�][���X��>���VZj�� x3ޤKȨ9gf�"���G�p���O���;��#�|j�pͬ����6#�h���X��餮�� u��1.0�!}̍ap�w|n��p��l�<��3�1ߊ[X9[����|w�.&_!>4��� ��g�����c ��r�M��ˌ�l�W��E`7�����<��?��+���;�'�.�%>��E��sH��81��Rw��� ?;4�ęiy]�x��ܤ�u�;�x��h�h}ФX�r�m8����R�rH��Ǉw��g�WcpB���ݲo��<�����N5k�ٓ��3 �p|�'K��+���l]ߜYi�o`4��*Z��<k�	�8�-G�⌃.%[�/v��M�4������ԟ��諕�Ttf>�P1�}O��Wh�P����om��ho�td�б�0dX |)
w��oc�F� �[���o���\�pe�}��o@���v3aYS=IXc)��E��(���;�{�ȴu�r���[�_c' M�ح�X[;�l�N�0(S�A�β�b�i�M�γ1��2CQ^�~�S�6�TξJ��r|D�E[(�R��D�1����!}#��Y������yp�`Nw�ߴ?��FT.�U�9b9���o�~Hz�S�<��s���f�`��K݊��6�8�<��ͷ��h�� |��
V��'�oZ������}����˰. ��՝t009EPs�����C�.�h��
g�����v��P�}�,�ѓv"���DQ�ˋ���A���?;���4�{"�fN��"�?{R�q��"�2�dY>��L�ɋ�W�r��o�˟V) �ΕR��Uy��`|t&�-����./̟n �q�`�O�}�І�$G�W谷�e�}�4'����y��+e;�z"�3^�jt� ��!�z��+]K�Fu ~��dB�y����/B���?�?�x`Q���<тx��B�1c����7�Df���;!�u�J�M�ӥ��R�	T9������婨�Θ�ؖ>���Mx�jAc����O���,��ozT�z�"z$ �9-����;_4�*��p�,�q���L�ǉ�r��Q����`=���>z���l�]K,jFI�T����5(v�&��g�(6e�H�0�C�YR3�ᒮuw �:-CC����׶��;�^��ȬjBu�i��j����Ԟ���`����S�����hڸ���F˸Q/�#`�}YՋ^��H:�'���җ���J�>�����ɁԃJɇo��&��H3ղ��n�{a��mv�f��J�;'�#�u�h�F}��>�`8�q��n�R��o�w�MA㧏�L�9+lmUɻ�.�Xf����Hϗ��'K\���y�+���31~PS�*:5���(ف��Md ��eɎ���`���{΍���l��yz���3=l�P�_�z�zu��7�oVL.����l�x2���7��le�N#��M��R`� {�'�|,]�>R�Ĵ``����35\2�b��NV�^hHǗ7u�M��&0B��k�/����4�SW�v���ݾ���[�F���e�:���>�X�ϑrd%����:uF�HkF�f:��QwC?��5��\+� j)�8�z�
�������Q�ʞ|:
B�)�p��x�S_���ր��j�>�0�+�ւ��j�+�������/z���A�pik뉇�x@�]��uX��W$�T,��-}2#sC������(+�]����8@�[����݋����T��G����cBuRj$�a���(��R���Z!�Qv�}#b���rR>>�P͖*�P��C.XoǬm��ֳ��@��(WG�B)�q??	[;Lh���fS�h���Pﶭ�'/�D��+��x{�m��u����*�=Y����
k7p|#'�zl$Uq~�S#����_�b.ϥm�4|�C�a�0:/�N7�0���h'ݟ��b���As���%Oq�(���,�Q��%�u��1e���`]>/#�s=R�>��<�,nߕqs%�	��Y��\�UW���[��]�N�`�]�.�qV�P�\K�w��4G_
b��d�� �X&x����['U����ڥ�/��_rѳeP��S �6��>s{u��}ĕ$^�����O�P)�}�k�bwPVHN?���y[�;�J=P���^�>$�[@�� ��d�*Q��w�a��I�³ ���fT�U1�}g�b���T��lR��kk3։���'2eD�����ңp���P��#7-�on�`�;[�G�{\� ^=��`�R��r���4�..��85#&〈H�GY �C�z���s�5�J�� <e>����U��ӡ"Ǫ������6k��HL�V��H+3`ƺy ����i��;�� ��
M%�9]6�<3��f.��ۚ��GV�9i�0h�^�ϥ82�l�<�\8|�Du���8�,�Xr�w�6�} �F���{��Y�,������%��{ Vp[�23�lo4尋CϚQ>���[~1�E�!L;�s�nR��c��X�QC�VD�J��|ǩ<��Xy�Xˍ�߬D�.Q���L]��	G@���\�C��\L|�Sf`F+Q���m)3�T��ދ���;�q^���YQ�F���(6����_h��ɯ֒%T~#�ϛ������+������	�p�=@Ex�Di��)��h�����t�]�Yم�}ե�bT`�̯i�Өݔ��C��C�*�g���gK��G��՝��L2m���l�gR���@v��8�����ǳ��$Rz�Y��f�"ˋ��[�K8|0B����dg�Ah7�� ��?���Ό�A��a��h-X ���1��
E;F�g4(�x�\sé��̳� ʖV�̤I�LRC��Hn�����2�}���s T�!����J]M�_�.�h9��[��f�C)��L&J!N&����Yr�� ��.c����)e�h�ޖ��@e'w����匊J��6��,uO��2�3uԱ��^��2��&К�4��uiǪ�����0�YO|������G� �ܨ��yG�/U���R/l�"�s�����8R	�P������>Ȓ·�wd'�
�q5���x�]��������P9B���������Rhj�f��eՃ�7��g�u\ַ<K6�+�Y¡$ȫ�s)<6F��oV�_���c6����ji9��(��%�6d�6,g�(���A��#�a�1+8�\϶��^Ch�R�.��� ��|a����U���(�xHTG#q1�Ɂ�
��z�ϙ;��~��q�r8���"Z��2��(��zP�IC:>�9�κ �́��'���G�MH���k��rn�t�Z,�B,����V���c����U�Xu�ķ��b9M��I.�>�3]�0P��BOl�{lhx�{;ξ�7r���7Î�O/�.qR6��5>���D�ae&��7 ��t>��!_ȦOĲ���NY�Y��y\�YB}�W�ܹ�8.z��Σ�0���$+�3�!y��L^q��m��Qrm���]b���,b#�3�0��&L����j�'���s}�(�X@��JQw�+������%��U&+?�9A,��|fє�h��\�<�,O�!�.��ʲ
����7dhg\5H"m8�m:3�Ԕy�L�����?����*�y��z����+-��;����bX�U�x(�g#=� �I�(3BJ�x�k�Ѿ~�j��(��`�pw1��I��� �����+�x�q	��g�<�T�_�V0��D�t��vͬC�gx�M*k�.
vn�lj
és2y��|c�׳z�r����ߑ��.�����sm֑,s�QR]�[���ފ����g�kT3��%%vX'�i�2~#�ls"V����f��d`>�e���,��͊ۦ��L�c�zru����UۥJ��SF�C�+�:%Q�c���q{6z�����f�Gce�9�A���@Jd�L7z�����ii�(����׹�Q�x�E�㺠 �/��\\F���N�A�o�w򀾼'�<��ۛ�id�V�|j�HWϜU:��}v'����a�Jɉ�a�� aҔr���w�ʇ��"\%��.��ж:Ϊb�!��S�W�K~w;l��'�=rRJ�$�^๤�9�,�+ۙW-r1UJSC�zt�~G
��p��S�{�~^���$$|���+mB�l�l��u�����+�y�Ca��ǀ�O3��uk}��S���%����'��᭙�� ��/�ZG4:?]B�{��\��b�S�M�o.=�T��倜Ӟ�3k�
��Y�����4���'�T�5f�@M��Iq4_�<כr\��nw2yp��!j���(A�+�b�������)��u9] wq�]�K���ݛ]�����,�3����uv�62�R<U�6�W�F�By���ki�|X\��:ԞH�ԛ�"K�W�W�'�+�$�&y���^ݼ�O���Yk?/_�&I���v�ɓc���'��WPN&��ge�Z�<�1�]�BI��'� ����[�'E|�����QJ;p���D[�ƞ����B�>S 	=o/S�:N{��9y�9l��K�e����u'8��/c�U?l�X�[:����{y�: 4�2-��X��w�`��g~%�vj�N%�(8- ��&��MY�Kh�u���:I��S�lg�ӣl[[I[���D(�g&��r�t�q�-� H�9���:���T6\	?][U�vr21��h%�k�RF:_b�ʍ���J��0v���7Hur����c�h!۾W0g�BI�����[[(�FL��L��d��)�M���8���L?�I���4�|��;�x�^D���A���z�'9���^�q�$S$a�iׯ��z/ӴN��@����n�r�V���C����j9��J��;
GX��"���@��Q����o����=F��)����$��{�`��Sǹ�)�s/%ʲ%�_27��/�#[�Շ�.w�=�K?��=��'�@&��^�-@�� �����y��/��2˔���4�s֕?��w��ٻ�ԛ��O��4��Z(��ӄN�S�����6�m�#N��1�}j�������h����:(^�uWB�+���^��^��97�^{5���"zMz��Ԙ�!xu��0`���GE"��g�S	QH�\�eC��n�5�r�������?��'�T_@��,,k�D6,�����D�.Q���)k��+hWB���1��c�����PI�&���"�M�r~���ܾܷm�E�bH(w��XbQ_�u�5b%#nfv�����U�Z��t��yIi���t��xP�5����|n���9�ڕ !qP�j߃�<��m���-��UT@�,X�3�����&v�H�Hu s�ה������)�#��cM�6�ɋ�i�R:�&$s��N���0�H&�dȨ#�9���ע��6H�J�B�_��M�d���5��D,ݲ�;%3��*�JL��Mڀ�8�K��u�-b/���U�Ҷ�z3@r��a�:���K�1c�2EI����p����t��/'�?nq�3��~�I|G�c�ݫ�'��U�˞�(4���R?�?2T��g���=��X^�+˙Fmp��R?$��-o�(�kx��4�wS�u,������!�.����m��'��'�ql�sE��ڧ���E�L��ӯ����D��Q���6�ۂ�Dt�ן�ө�Б<~ÄI1��G�Ǘ��k���hR���������s�i�Ol��g�A�8�T�r	U���a8ZJ.��"t��>�uČۼ՜��s׊�2��s�7��������|�WWn��'�F]���u�pG���YK���T��Fbik�6-��K0�g��"��k��
��U~�,[	%��s0��w�!}����G2��-'����(��DP�ѧ��f���e���`�&ڗ�G.D����X��h�Q!1�7�}��+�0����U#K��*:���ZMɦ���/��G��l7��=n��zܟ&.����UxӒ��}	��R � �J��o��������i��I�;ǟ:�:��D+)&1+<V8�\9�w̮��h�xD����1��!ҹ���俽���> ���Ձvv�0+�5���Em{�|�\^ ��N˄׫d�e�,��.�JCxN�ˣyL�"Z�IN �owuf�I)��!�C����t�-s�D�/}�7~?n�?`w�4p'���?��y��u4��8���㵸u��"�	]��o�|t���d����5�Rs��cd�E�9����FM����*#Y۰����%�!�\��u1ޣq�ɵ�h���{~�-�(ucd'ZI�;W0���p/�i�v������\\o����T.;��?���Ψz���f+�
�sߕ����E$��T E.�@o� |澽����>P��O�P�S̀v$�:�C��,��JN�E!e,&�c9'��{0�ݖ>�0�oF_Γ��:(޲l����m��R׀���5 ���X� g/R�F}8����\4��~�Ԅ������]J�H��<r�ví��A�k:�X<=�6�����x�B��>Hd��KД�Z�\���u�D�a�m<��R�ٜsS�.�D��&��q܎���;����)��!_��۷��~���ب�����`�G�
l��^V*x.��D�
�B<yLw�j/�!����(�� �ne�2��8�dk4d���Z�j�e�'I��(sn!�������ӳ�z1԰���˅���l��x�q\/@��^/�����$O:L�Z�A�j�H,�}�	�U9�j !��0�>05�1D���I�(r�w냴�J��X��	��/���wQ�9]F;PʅsD�= �je�b�_1H�6*��T߹��0�ALOI��j~p���4�d��ѥ��$x�V�Ic��DR��-�u�c��Y�m�r�ZGF�����;��T�pHl�R �Y�5�_�!>G��Ϡa���J����G�Z�� qO�C��h��M%��=(������@�<�v��i�����b�^C_���'�p���:?���)�gD�_��橆���y1E���c%I�w�_��E�6�:h�\���6~�V����D�3MQ�����o	��]c�n�Wl�0��� ?�C^=�l����5���`�R�}��Qp!O�ƃ�g\��#�v��jo\s�Yz'�,zB Zd�OC�\~_<��Z�Tt�e�F��N3z�b�X>|;�h/}�B8^O�%���+E�?t��Z'E`�k{�(��%;o��ӣ�w�0}q��j}oa�}�zmoS����$�1v��(@l3�\����טk��`X�}I$8���3��P�x^�'�
���b���!9W!C�pw�B����3D��4��3��=�$| ]n.�������*x'� ���s��G��|�j<�H�bE������J%�O��o��(C˃(��ap}�}����(H�J�[0<h��<Z�n^��]E�T��lo��p��N���'����С�T��Cf58�!CB�����6���t���)�#�UȈݚ��ʆ�
��/�"�!W�A(x�y��Ƥ�%)��Mh���������,a��&��P���\���0�?����Z�Q�����D�KǁHy!�-@R�:YtdW���
BJ#l�<R��+���J�֑m�=^���ن4"�c�z�m_�����>S H���ぃ�J:��I����~{T���ɸU�ރj�l1f��nʭ�:�]�bW��3rm��/h�df�EJ=櫮L�~a�|i��Pp����Ӳ=�,�C��h�M���y�t��.vl�
���!��f	�{���m��0E>k�깷���@3s~���
ރ1w�>����� �ø죡�`ڦ��c��x��S�QVC����T��������;�C�A�:���沟�7庹�0:���}J�.)]�k���h\��A�`�rGz@��j�������X��
�X�GFt��J�-k����
1zX��#���pǅ�J�P�!��7Mv5��R�"������f�-�e ����Z����=�y�Dj%���S\���~i3u<��Ap���Z�j:��&������s;}}皥ΰk�Ո����5����\�^�C�ڡ��^�JV��K)Q�&�@7�G��62�b�el`.�*��0���U�)8�f��ŕ6ފ�E��A5ī �YѦ�# �!��|a��+�a��4%1C����:�����1pi��:��b�j� �^1�k�Ϙ�R�-�;8�D�!�Ծ�b��>�9�������!�C�Eʂ��x�N\��޺=�)��o�h1F��Xp���	�TJi�"3�����↢�1#�2�v^w�����`7�@R�a�	�W $@�)4��'l9G�S#p�H���r�c5λQ��"0O�l�`�ҞG�XĉRգ�͐�������Mߒ#k\*�i�[K�rV`H�tR
m:ܖ?;8���u�>�jlԺ�2Z�6Xf��`k ���B�݂0(N@I�����D��C�n�<����DԴ?O-^­�f��C/Y^J�ӎ�,V��<;`�_�!��ro��ǻ$V�D������,x%��|�>'�G�8��_�A.9B[&B%�IV��Kw���;=�,�ظ�����:�0i$Ρ-I�=�,������p]a��Ͱ���{(���T�f�ɀ*׵{f\���#��-6C��5���!y{�d|�_*�ЉjI���"��qyp��{d0��L���G���츝���J��uGT��'Ԟ�i�qҀ~/�Z��>`!&�F���D���!�p����Xe���1�`�ٓ�+V}�oQ��N���hMÂa�W�~�2��*�4��CH�S����ǹ���2'��������_�63Ç��MF+����M��z7��7e��JM#;>$�H�b��a�����%x��oͺ�=_h>;K'�L#/{���	6�H�<�%b�S�����gmt�7�	z��ݧb���x���;In�Y{���{�i�"���&^�
势�������̳W�?t�v�k�t�k����2�����bA~���Y�?Q�F8��s%�n�e���v�0GrS���~p������1j��</H����H�6K/ O�^ׅF@���a�#9=h��݇�t�e�]�j�G89G�����³�ԮI�F�U�c1 Yg�y��NI	��|5|��/� (�S6#45�1��x�C&�ü~�\�" U�3+)@PӴ�x��b�����S��z�ӗ��(�A��ΤK�Ȝ��D̰��n]�Ts�@d���3D��Y)��j>�CA�D�i�x*%���K��~=К�Ds������a�΃�'���0%ߝ�/�Ѻ�
��π��>����Z5�X�j�Oh�ۜ[)k��2���j�8Q���Sg��`O�R��2�����79�A0B���yV��po�P�.z�|:�d<���Rj=9>#{"�_�>cF�&���)s���&%qX�?�߶�B����Z��)���s^W�*4�m��M2y^��G�"83�ge��)��9b��WmO��G���ܖs=�����Q��%iE&d.��f��_�ֳJ������WY@�Po�r=�p[���[o�p��8�BIc���{� ��p��˨�9�<�������]��t@1|NZ�X<�*������*�+w����<�o����y��p4�灥U[ǤmV�l��P�i�1G����y�K_��;*w{�6�O����Rί�a{�#1;+��dh$�L�!v_@Xby~s��n>����`�:+�$���A)7nزue�
�աϳ��s�;C���gǭ�����z����7��:X�ޘ|oS�͊��t�jbW�~f4�Y�Ѡ{A�c���J��aiR�h�"�g�q�~�P7(,���c)q�6J�{7/PX=���B^�uǉ�����s'\|�s��-P��ȟm��Ɯj�?Rƈe��s��mT�+�K�*�,�)W���r�J��ew0m�ۀ��Z�B�P��CC�8"*������h�^p�K��˂"�BR�y?�[��wW�:�,e��j;z{1ٲ|�Y�
��z�caQ��>￪��*}��J8�t����9����������.�?w� s��C�C�ӔT�t\�~����qZ]��XǦ�*�ѐF/�A��) ov��s�����9���4]�������^��ܵtXL��4�����(��4�A�#cu�/��p�#����v�1Bl��1��݂�[&0r����k�}���pt!a�R���&���oK�sy2#�3��5�n�Z$�(�5D};�U9S�$k�����!��!���.o��B�m�����>)i�>ĶS�S�mz.�φK�YS(��,R�
�o*��q�8�����
�����ض�&A*�)��\��Z�8�����|d��3�������~�y<[�K��I���֐:�F�a)�A�l�� �����u��.��8�����
�Z��7/W]�������{P�����,�R9��
�Qcdxq>�E��l�r���֩���%@����~��Xi�=m�׌)�0e��1��(��sa����[k�����f9�Q��98d\�sԡJ�G��)�9V��ƞI��_�7DO�nHh����7x�[.6c��4Lv�Ј����ꋻ\�0���Ӭ�_��]G���=y���@>J���J�As�B{봇�,_0ƥKQ�}���U,�m�8��H�{=�?�_�"�F�E�+)����|�h��f�W�}�х��������;U�\O05�	����b�`6Cu�	j��4�R��g>�3�T��8�GGY������n��8͞3�hyW�|� [���"`�zR�C�u��$3�g�k/FP�y�:�I᪨Fk��F�&5�,͒���Z��},��Ʉ�+��]�c��x=Z�쨝������4_�Yk����F��0jv��Zΰ�β��4�DRUC}NO�v�n���^�Z���;J��rB# ���t��~�fa�p@��p�좿���SF��I���u��SH��x���/��F���Lɽ<(�E���S��"6C�4H����m�����؛$8�'�O�oP��"Xt+��`K�E�F�!����v�����"j̰SuY9�}2�V�dӰD�y��}�rM�����z��d7@��5��	C�w�KB�w��\�m�T�!�H�c��l�4W�RVXd�)�'ϧU;���t=C�Q�V_�������)��@�UubUqB��!�)χ��R�:�B�B����	� :S"g��b�p�����ࠊO������J����J��N���Q�T�]��\pm���N'�)�Z<�xȒ���:$�oVOMr2G�>���ףЪ��q�/����0��UY�X�_S8sO����B*��)�^��As��y8�\[ �P����8/�x��Hg�k�������6����I���� =��W'�K0�	ޛ[�h�D�%'�E���6�bu�QW�P,���r�I���) ԧ룾g��bY��t��b�����X)���k0�hAq����R���DEl�j����o����@�l����P�N3V�䬪��F�	�c��Y��>��W m���s���i+��s��r#���d�k�*~�u���������y�}{��	��Gk�yaZf��Ln=�GOL�)�	��`}R�.�؉��=M�����t�HK���K�CM$�Y�rq?W�B2�n6�H��Q|w�o�`NH� ��݉$��P�G�L������/�� [�ʸ���uS�~M�*��3B�]=�Խ�+��Ţ-�����/���v�e嫦Ҟ!���t�	,BYo�j�w��Y�a����5��[�x�\��w_�ɺ#3��R���d^�@��=*�S�CZ�40��w����Q�i�[�ಅRE�TOb�~���Hd5�������t>�D�@!q�ӐJM��]�G�V��0H�AD�x%طv=A}W��Y����M�8� p�$����I�u����>��o�!���ї�-�s�b2'�.��Қ}��)�5��N��\�f玐|�,����\�r�%8��:U</�ĥ���h�5�y�dM��6��E��:V��}����nBw����v^L��v��P�_o�2<�ީysX�-�jo�Q�?�$�dE�m���H��P(�E�V�a���hL����6ꌾ�O�X4P�{�ǣ�'P��v��cC�=��>�ϻO�]�B�����-]��਄��m��������ւ[�@�v����D����T�@&����/ 4,n�s��9���኷_��TL��wfrM��>s�&.�9/��+��BP���x�a��G�Gs`N�A�y�X�`!�<;ܞf�'ߏ$�k��q���4ط���n�f� ��8�:��h�����X.�;q8�a���4\��Jy����P{XL���x��L�>]!{���``��,DE��ķ�� �E�/C�^��=��G_f��qu7/�D�qd�ߚ����S�㎮��6��I%^�����܋W��X�]\ϋ���l�M{�,��w�J�5���IN�Q�@���ӳ�*9f�H
$ρCo;,C
���\b�;͛�j��6��~l;����Y�S6]�^pS2��ps�9��)�y`�e�6�N鐁�"��!�D�_��-�\��;���^���{2�H��B!��������U�u��iǈCfv�b\,n�&M�}�v�����e�|��m���&���༛�,_T�r_OZ,��:6��e��I�9H��jXG������x��F��v?����\��r#��yB�(N�8��ѵ1��Fl9I��FV/��������\vJv�b֨�qk���D1/%��	�5*��\��	�q�0Y?���q�����h��S����}~��t@ҷ������%�m���yٻ��3m�- '3 \:��xȢF8�;-!I���sY�ݎ�z�)��>�#�2�z�,ttJ��"?<��/�WmT�w�YJ��a����l�h!���8�0���JVU�U�'���DAj���G��:Y�V����_�W��������&��ggȭ�����f��`I���{9U֭��ج�LJD���.,g#EQ�4!���P�ktmm�k��&�"3H�*`^�S�i�6�>ok$���j+��������@֚J(����Ƽ7�^�`��4�f��ʮUhb	���4*��ȷ��;vf'��5�@Z(��}9z�[b�q�aT�"um+��}������|t��׀��ʅ�J��<�#�?R�e.#B wp��Uiܡ�Qݙ`wA�#�A����-lv 1WK��RQ�8�����j�tCd���\w����Ui6-�� �GV��_r9ܾ1�gy:Lü�X梞wb���lL(�����w��H=N����`�&@a�6��F��W�>!l���*���#N�psDL�S
��g�Rȿ��� �)[��&�	/�ߣ��`fٻ��+~�7K[A9�׮N�dO�3����B~����7����t��z�$r�ﮩaV�άK�#_�9�<5A�\�ƀ|h�C����uzOF ��sޮ�<�Zp�, �s���Q�U�X �m
��"��\"O}9��}���k�u������%r��)�-���TD��:�~&��@1M31���i�X�Ya��,��Z���,�W.��Xb���J�d�|�aA��^pߦ�m�7ь��F[�R��~���(�d��s3OH|Ո�/�e�e�e���<1kd\��|o�E�\G}^u�_�M��l�M N�p}�+�W������ݣ�(K�ۦI�9ž�w�x��:x J�^��f?�:�q{���g'�؂4Ē��-�˂��Y 4�b�RB=��ߑBy�����x�с�{��J���h2ず��o�P@�}|J&T2e&�xs]��e��U\�b��'�ȧ�n.h��x��Z9L]$i�	a�\�w��8���G>Q�CMb���1\�pړ�@�AWyI��Y��c�܆��gC�]�]���JRݫyjG]�_�jcq�W���Xt�Ile��ayl�T������L��|A��*8�{��F8��Қ��|+m[ME���R� e�
����4E7�X�_G����b�t8���V��nm�귰$e��\ów�eb?�Qr����E�Ʈ����F�s8c����5�	Y�6M3�!�;�H�틣~'����E��94h�Nț��HE�Ň=X մE�'Q���,��o����{���й�@G�bs�M���^��lՏ��WHv��5_m�M��;��&>�z��RI�۶wB��v��`[�_�����5�S�~zb��Q���	1M��s'I�qd��oA�W�o�0��-,,-f���	��l��o��/�#�����g��٥y�kԗ$Q�
�Z��bB���$Lt�M�U�2@��q�N%�{��"q��[��$xL�[]�1�s�����6k�3�Qi"�y�Π�3eM���&L��R�|�6��$"�N��7��9=�e��!��w8%���K�Hd�+���v�eI���Gb��V�Ӧk�?�N7��5sA'��o�q�z�^y��>%SJ~�*y�z�k�cF5]�C%#��0��$�]�輽�����s^A~^�~��#,�?��rpIȴ<6,�6�C$ۿl�����?�g�\Z}̹S�+Z�K�l�0������	I�����/':�FY�\�9a�1���9P��iK�7�f^�<��g�,��:w.�td�h��0��m�uKa�!Ų���nحȴ��2v_<	T�����p��#�aL��� �:D#��'&���(FYy��\}������@D�S�TSQ��-ͩ?��ȩ��µ���.�-5����2�h.�4�ej�bK� 90 ��8���3GO-��װ��5�[��4��s=�~r1�˛���:L��TLV�j�-N�VE�	^F����ؓ���DI�^�>���7�ۡ�w�t#3���!����A��i����8���������$�M�{�A
�ؼ]}����1�+[SL
�l=;��4�#,z)jD��!�ū���0&�*&���D)�^�"�H��a�v�r�r0�����%%�9�ci�^vU ��RZC_����
w���m����IO��6�.�-�J�O�l~Fv��/j�e�tm�/�
>���Y�qd�\��B�Af� M��&vi;�8I
��*�p�䃂QV���P]5�)T��
vϠ�Y�����5�=jEģ�p���~>6u6,������4ы{WVń��^2��b�/Aa�2�3�+�ӝ��g.��3G"���:�6���HLR����=��j_k���}>��<��)e8�(�}����ʶ,&����E8�9��+"�:��{>咪�bLa���|�̱���#��}P����T�F^�5[ �!��j>=�/�`�/�~@��}�G���݅�R�ɦ7��s>"2J�S�\Yآf�!P���_��[�8Z���wT^Bj�/Z��4.��7#o�0�e���;��X�X��՛��D��r�
vM.��#�l��8�Vi��[|�t4$� ʒ�ܚ ��7��׌�,�.v�vU]�p�^����Z�H���O2|m�s��7j���	�c�#��c9���o���b�7�F��0��D�kR����z��1� C�R�����ȹr��,"p���eyAGj�'�8W�'��[�6'�������=ގ�h?�yQ}���)A��K5S� Q��%Bf�m�o���2>&d�2���"�8J�y�qo�#�b���栅ڤ}���=��,�p�Tl��5Sdo��fvB`�j.2�G�p�\�v��@����m(�<��^%�,{��p����h�V!���(a�|�a��2R��
�׶�K
;?"h���?����RJE�s�a�+
v�>`6�k��ᯣ���n��=�摁�s����37��R���H���6@G�b�b4H�m��G'�5ȶG��h��5(��8��\F �`�l2QP��[��'�՘�I;ʂ�a�=A!��^��YN��i
��nĔ���p�V�<���9B
�bl��B�1͉D��ᚔ�K^s�`��K�Ww
w\��軕���l�H���6���W�w�DgP��rSO�{����F~t�]�ްD��b�/	w]����]���.���`J3ڥ�80�tK��4�'"�c����`O��YH�wA����A���=��c%����n����b�0���R��4���{AMum� �q�đE�B[I��4�˟�!�����͈���{�U����.A�W�6��GL� �v�;�ւT�T(.��u�-s����q<wC�^j�$F"D�f�I-Q��4��(�ç�{U�W<sMI.L�?A<o��Dp�яx���ɾ�&���wޣ��0�s�ƕDJH'}�0״�gI�J
�ES��^��c�\��p��?���_�6c�tL�4�K�\m��k��P���7j�5c}k���9S}��q�>����H3��N_����N֘����5�����l��1� p�i���'G��΍�q�̬k�����_3�"F�4&�gS��!CYG�BiȾح,�ce��Lʱ��#%���C�H)�h��m�σrCr�Ĵ��K��y��@t%wL�z�8���9�u_�gO�'�'?���X���OY�58�9��a�G�;��E$��-��q^�6���c�����U[>�Q�ڏ�F��c��4�#��aqW@���i]��8����dϼ����%W������s�R4Tg����?.�(�����*\4q�����"\�]�Db�u��>vf� ���p�LzP��1���pO��LAV�IVw�R�a$Ϭ�9�> e7�^>����d%�
#�e6D�OLhML�P��dq�{<c�F%�f���z�'^EU ZWe�hg;�¦Kۚ����'��,j0�"�cS
7�Lr�m�Q�5D����M���v�0�L���VK�r�ǫ�aq�8x�9��`9K�Ӆݙ��5� H�#g��`�����?��zs��L�ˣ4�>�A�?��Q�8N�Wk���a
���*�)�����{F�Z�]�ī�	O�"����?Tl���� ��:w,C��m,Ga�һ/T�֐{r,Dx)����y�|��� ��叡O�m�[%=7NlK�%9tc�u)��Z�?�XqP��Z�)�1z.C_��uB����Hl�\�.��q&������.+� �f�"���
�K�bh�mVB(�ߓB
�����=�xc�_�#�'��D�T���>�Of3 �AS��z}�_.�q��u�����b������h��n�T�`r�|�)P*�ŷ����i�G�PGnʪ�H5�"m���������t(v޵���Fx�+���� u�\��ө
��ط����=�Sn��w�#x���iJpr�?y�U�ܪ��L.�-�	
��b�������އɪ��31��!���N�~`G�9}����c�]�
:Y�e���s��X������L$�(r��׸"�}{����0]=�\�갣n�(����B�F&��>�7�ʗ��Ge�D��]�4�.F��`�PZ��@��&k�t CL7�s0�l_3+0���0#��/���$e�7�S�[�rfy�|i�L�Yw��F��Е��z���pK\z����o�Q,*�[t	MF�QO��ޚVX�����4pe-��S)�]�;?�ݐ�\	�><�Io�<��:D�Qu�8l��p��$�w�kS10���XW�J���asѧ�s����J��f��]�Md�$۪GD�0!	�(}dٮGC&� :�%z$F��DJI9�q@`mxQ���wy<�ۧ|��BO�MT�{�%��$���O��Ě>����u��|?%ɬ]N@j�F.[���0>,*B�����Z��}jw�)��w�W������	@��!�8L�p�hl�ҫ3d����R�̬�荇j8�ްi�G��P3L
?d�
����������m�������U-��ɗh�_d��1���Xd(=�B˗еj�娞�X�!�+��ߘ�U�o�yL�V�bq��T�=O_M������Q-�d�ղۺ}"�u�IA�i��~|�:�رW5�s�.�i����Qy�S��;�1H:�.p���b%F�9<[���^PY(|��@�*�X����$�iG
\5���8{�Bȴ��.wT�����Մ�� ����/Z�<;�m�"����N/���b�7�gu�/�����G���X��z��\G�ܣ�Z�'ȝ]K�-�����^}���ITm�d��k�)\J���}�]�s�FTu�(�5V֒�QlCL&�k�+�����<k�ԇ�]��FÄj��L?��X�m�L����@��Xk ���j�T\C��G��6us7C�Ӛ��ͣF�1r�>9A�wmF2�u�9
l,
d+^a���ƶ/��*�X��`3�$��k� ��4���B�d�����kh�����Ա?�\�9��z
P����4!e�|tP;�\�H�j�d��+�Pٴ��Z�d!��Ŏ{��X��眊^:��0�-�ΣuP�˛b��z�Y�4v>�by4y���'̫��t�V�����A��n���i��t���5��7~7z�mh��<�f�����N��2ξV�x ,eL`�v�G��X)1?�a���8[�ը����5�ȁ.垗M9��k��v�l�z�n�m�䎲�:�F�~��Oَ�YG�L���Vr���ߍ�W����t܂���Y�v��;$[��2K`���w��e�5���oshnw]�O��G�4NS����T�l��9J
%�5(�c����?�f��c�&���-<-����g68����~)-`���-�Ai�đ��ah��-Ǔ����8�P�� �t�3�=gq�E�;a���l�tf�K��W!�;����V!�(�f����8�6X7C�P�.	��RahwShૣ-��H���Q�}��|Biv�����OV�7�x[����K3�0>ym�Ϫ���jT�Yo1��!��f��Y�YYB���M�KM�+`��
G4m_8�"�z�/��@C"��~���;z�y��b��`�z6����(p�al��u�����J��I�h&q�U�u�65+d-��u�gxG%&2".��WQ?�^�!�#�e�1"l �E���6�+H�j��Sc��jr�f�>N��ߊ�,k� Mv�&_�f+��v嘾(b�bṡ#�,%/t>7ڣ��h�8��s"�n���_���yFE��_nUA�Z�F-b��6�R���i�P�p> 3���b�ӳI�.��<��?�r�G��2��� )1PFO���1'����wPֳF�+�%�y�ױ��Fm+5�|�2x�=��,Z�N��c�c<�
Vu���$ɶ0���J�QI�;��M�f�����t}r2 N�2^P�`j�I�S���in�W��r�5L�J������s��=�W�"Cs�ag b�~������#�c_�'�O"B�Mٕ 6Y'~P�LQ���C���=�O���p@p��N,`�"e)C�=�,�js��CcU"��~	F�F�����y�iʑ�`�s����"h�^��W�m`�Ω}�K0XI�Ě[0.��_
D�oχ��2A��P�(LGx��-�r��E=�t���z�7l�i6^��?.��=Vn�Y�Hj�O���cS�`��~P2I������/��_���:c�]�.��w�q�]D"�}t�КD� l��Q��n(�*�ѸG�� ��F�s����O���

�N��h�<�)�m�w��-zh�T�����r'^Ғ�&��N��F(�\�}�aB�>��AO
�`��n��h�eV�G��/����|)iTz�Q���7����!,�_�z\�5����e�ғ@�Z �$A�^BB�6�L*�򱌚�	��D��#t5Z�B��f�%�G�r�0�Q�/<�HB���t(r��~36'`b�2I���&�君����_!��j��uc���Q�,��
�<���ʀ��>�`��Nl�
����\ ��7���B�v�s�mΈ����	�4�[��q������Bf����Y}KZ�ppLê��%u�{�5�Jc-<I�ܻ����8)��|h2�(i�)�K�Of$9d��Ҡd᷷�r�?]q8��ҙTډu��Bz�z����S���dJ:��_͋�}�d�SL���4T�!�����*�>��c��{��C(Y���1ʣ���5!ǝ�K�. Ў�,s|Z���z6����ŵ� ՞��[KIl�b#S�겆���b�$BY+f��<j����%����2a84�q��nV6��e�㿝�������BUx���9�Z�lC\��I��t}%=�	꾫�����9�p+����5C��<��_��_ )mVI��<ƪNueqO�΅H�.��i�W� �7�sY�zx�􄱹���>s.�����+!��6�|\�n{�EQ����������">���	���l��ӅQ���Q~X�J=�r����=�裍E=��D��6`��*cל'/�O��A��N�Z_F��\��%�Bd��4��`�0]���M��~QW�
���E�����]y�Lo����\pQ�T9PLC��T�͎���f��V�Cn
I��eJ4m��>��թǱ�F���6
�4	�ަ�L.�蚬�}�	��9_7�ś�qfdp����������`IZ{w��G�{�7�}Rcx[%0$ܼL������c����*J�&L����BAz����r1�9@C
�f�_<� ɢ��ļ��z0K��xF<��	�rb|�h���y�=ŉE��j�NV�˼rGlz�,�Uiz�R*#�#c�M��N�*� �6s܈���><��:�!
Y5�[Fq�~��@c;�y �
g���['J��i����h�䊗��~Fk�	B��X]P<���fK�M� d׸ew�~T|�s!����HCjH�C�_�Øj� h2��|!��^��r�>��m�x8ȉ/�����3d�j�-���l�� ��r4Ʒ>z�C`Z�c��.}S� �)%�$��?�#H;|b�T��8�-L����ҧxY��Y߷����I�
�XאҽQ�^d2'6��4ׁ��K�L�(=j�o��Ƕ�6�Y.2:� � �-"*�0Lj[3Fu�����Gd��z0���* �*�R��� ��Re�*76H�̺~�����]�!�T5L|I1����:1���~���YՑ�" )P�~L��@�@�2�AE�r.��B|-jWi@���y��������`Z��	�2���x�h�����Ŧg����A!�%�B��v-h����P�eB�4{oć�;X"�����������?��//�|?ܬp�����E��F6��G�[Vޥ�;ޢ� ,	B̈�����>�h����I��Q�n�D�
�#�pMORh��{����5�~��q�L�L�[� P.�fr����b� lf��	�4����UC!����Mc�_T��R�ͦLL��W���4Ϛ�;C4�v�QM6<#/A�� _{_e��6�k��#�c���,�鄜��g�63�x �l�y?B������̊p�,h�u���%���u >z��ʖ"-.g�q�[$�_�e
���oy܆dT��ZH�h2�� ��}��^-�9���#	V�а	xO�������}�������ǥ�q���dly<���P���:u�����$�.-kF�G{tG��k������vx�*�e~zC��,�y�#7Ov+�M��ה�Kj�!�� � M�^��1���c8��:�
�g�4��:�k���o����`�K#J��0��E"����U,���R�[�?�E�ʃ!�m���^k�Ȋ��fq������^�%���<��t#��FLī���2#�s���3`&�iF�v1���t�����.O��t���֕VZ-�~��c̗���P��T�ƍ��i������x���,��"��~�)����s���Q�Q]�������G���>V�R��*S�*u٬xȻ_�Ƣ�w䆅���$%O�1<Ã�ˁ=��
&K���`�|M��y5Y�[3���-x1_rv���+����>�ڌ?�5��V_t��A	>mU��ĭ(�c��E�{�bj� �F�9���ߨ��/2o�9����<�,J~>O�?��K�/��@F��/���h�'���,��j�qID��ƫ�r�|7(�Xۂ��f��%F����q>��q�\�b�)4x$��g�aQvY��H-q��7�-di�_z�T��o��=c�,��6�:!���ڿ�Z1|#v/�#ώ0���ޏ>���P��ZS~�g�m�b�C��vy﬍�'�+�c_��p��B�]QOd�>�K�Z��R��?�L'Kr�[�ZrBȆ�%	�i^���2�r�-<�)P������{\�$���$�+��\�������Q�*����-�1��W�Ǩ&���h&s@�ԁ���"5��:?�o�����0����ݮ�ܐ2�c�`��+�u���,�0 ��F7[�9in91��*=��Ka��Y���僨�xS��9�&o:�~�D��i��`����h3 v�����]qSI�g[�S4a�ŨkD=�6��VC����N���������z` r�<�T�d$R��Ǭ�}tw�}/����6m�O�'����zv�F�R0ݠ.������%�@���^
s�ș��W�O�Z���(��H����t��0&=m�����B3��}�V�M�b,�H�]�Sn�=��-^���n�I�g��r�[��)��rs�%���X���V���+i�TH�~P ;�k�!���W]�>�j�o��o��":Y�;Nu���)��GH2,�u�j����������x��Vsh??���Ő��WF��8����ؼӡ"4�����7�'�s�D,���;���Z�B��;�l� ,��V�n�d�KԥO��<�}O�#���]��KJ�u�Eih����N�%e'{��	.���]`�R��)IqP>��%��@<]��$�����6��Z��&��ڌDghk��7����} .c-"�[��q�����Ӈ�ZRs�e�y�����ڴ6���휳8����Y�PO��>�_�j|}P:�ft�L
è��D��	�W�j�Q�p�|N4�_�_�� ���Vz�0C&��d1¸��!�4���].����b�y�u��v���s��i��N��X�L�C��9���N��e�L�O7��K�y�����ؕT'�pB..�=a�s�_��&4��w/xI�G�_���r8ɶ�ᠲ*BͲ�8�
p�e�2�m�ظS+}���0���^��Jr�WZ�5T��k�6@����4������9|"�Z]^�.)zlk�[!.>]8�}�'�o}vcvD�:���Θ��:n?
�@���	�4�)+MybE��MF�0V� :��d`�#�3�� `�`�Wj�ڦ ���C:��4��W�9��ǽ޹x4~.}}�(kb�]�)�
�~��V�� xH��<NKW���g'j!�^�{�?(��w�X��=��/$����D5&>(���h����	�-)� �:Ɛo�g��h	�kdofo&�$jcŦ����U�F����D��ԧS�^�� $��q����\����+%�=��V�zߑ��X��ͽ���j�5�l��&>s����T<���y~ŝ�p������=X#��x $�#qT'��)=)�5�!�2L��Ƈ&kg���/�_��"YZE����s�(�%�P��x.J�b	3ꨨ�S�@  �r����/J���M�Im�_'*2�I�7��fȇXNR8�P����NQdj�V��gK��G ��r�WT���Q*�	Ydj@�.���� ���Sw�wK� �+a������|?]�	��KX�(�E3C�$,����tI oA��ٴK�Kd��8>y����gS�QE�9�u�:rn���i�VH*��/�Q͍Lm=��l!M�S�v�M=��ή6�lx�y��	Ui:�Ɩ�����ف-�erM�'��srE�(ְ/��,���Z���f������@	�������j����ex�X%����T�Ar�,I��ܒ��Vx�W��L����a�/�,��Z��^���"����H�'m!v��i��{V�C�r����}�i�\���D�ω/k��&KUkP@��K(	�wN�Ν�$�M�[ם����N�k��g9�C?�Ӽ9<�ed - �-�jƙw�N�ȹ�{�(�p,����+�s �3�i�>��y���� ,�B'���:~���n$�<�� �NG��%U�KK��(��1�S�@	���>C�$G�Т�t�O NN!5oG���9���J�����Ö!{������/,ӯ�����q~Cy�)���n�=g�d�P��UI27MZ�4��C�Fn�B��"�ͰÊ۫��e��p�l:P`�[D��dU���ZP����@��=�IP�j"�Y���-cF[�ͽ1�k}r����A� �ſ����,骙����+U�eu?٣/��t�ͯy?��	C�����Ւ%���z09T_wױ4$ϛߐ�GF�7���g��*��ƀ�5�h_��;b�կ��ܼ觓,ʧ��\�ÇG0S��`B���_w=�JƏ�M�Չ��+�^<H�d^�<��|�����U5�,�|���H����F����7տ��j��.�^�N�
n��[2�JWs`��Y�qD����"��f�V��h�����X^^�PS��l�������;k��(�j�J�q°�xd�_n�/3~Zet|����׃���tLB+d8&/�u @������Aw��>(�ʉ�3(<����}�#�`�F��p9q�cd��+?X�,�$B-8�6B8���p��I��Y��+A5ID	��T�Reİ�}Su|�i���W�*���b�i�*�"0T�%�{�((�f&\y���8C�rTx�� �!�$�*:`h^�#��KMf��	�	���Z�hO�1<�P�3AI��޳��U9rOz���C?���)|���dEM�2�Ȇ�ųfS�8#���=�>N�DM���,
(�E6*j��J�z�/8��Z1V��&�|7�&��>��ڀyp�|g���`���b%���P(���y��q�)��j��\W` ����d���F�;���G����l�VB^��}g]t�鵬�M�����N�½�.Ж,��z?`�yD��nn=�o9��`8���&�	���6}L�_�1��3�F�>�Z�+�J��P�TKs�ݾ��`�[z�o�	+����`�����F����{oWNx��P}%!�u�Y�W����YU�UpN�Tz������D�΄�6c���-y+�2��l[uZ'�&��}�z��U�Ȳ(\�L��24��Yˇ�8���B^���F"��ʟ�jf�Q���P��{� Q���?�س���q��_�FB9�\M[Me?�@���Q=d�-��P"4iV�T6���j���0+�y,^VW-�km+�����F�]��$EI/�!4�|Ov}ZQS�*b�" - �R�#!��0keo�d&�S��ش���3�l�l��Bq�@]"��Ǡ�
�b{�dgW��1)c(m�Z\�����pF�-@������fg�$@�+S�4kb��S3nI��x��~�d�yT_j`������pER,��0 �����N솲��� ����>��h��go�T�nQ���4�\?�B��zq��^04UݫA��-?:)J�(Mi<"��
�殯j���D�A�X'ǁO]�ae_�5|V�ӆ�l�]S��$ֈlXaI�����nE�~O-K5���� �L��1&4ۆ��R�jއr���|�?.d��qO�ox}��&�A�\9e� �{U�/�����]F����@��|��I�?�<�5�&'�!�wOv-���`����B�46��s��:�D�*��(b��V�n���4c���!���Ϭ�@bS�L��2�I
�0��bfeg��o^�Iz9�;�b�.�F�J��M�{'�ނp{��9P��J)%��B����Xb�aߥ�S�:�q�	�"�Á�}L�h����lt�I30I<C��t4�1���b���]>���*Y-��b�8�0%jo/���}ӂ�9F�-<'���wM�B�i��1y �����r�ӳ��ؤu1�QN(U�8�=�˭�k���Z���EN�ǧ��k����6��ζ�7< ��b�������1Ӿ��]C2��5k���A�H��hԼw{vR�� ��T*�5�zx�PGƆ��Ӄ�X�7���RFİ?���s�5^���#�߻p��G�S}�[�$}��a%1J2�>'9N�ǳ�~Hnژ����0F��p#ëv���5m2��t�N ;��:=���).���������e2=�J��Zn�F������J'K�TAi2��[Ʊ���gapZUgφ����n��q�n1p�%�M�E\�$1��Z3��\�v��+`C��A������.�>J�~��F�:������c�]��hRM5Σ̋	uX@<�5�]��8���u(��E��4����M�h/�]��(��F�L'�@_�[�F��6�E�[BH�ݡ'E�;���wp�m�����3�h�C�U}���'�7=��"T�p��!4�uZ����xi:���A�A��ھ@)�A��~O�^H��R�m-�XI���y�MÓ�Y�<d�����#�q�T�3�y8[��4�M�kA3�6�*'+���V/���8��ȡXq�6R�}�(���ʴ��vGd&�(�~�M�X��_�h�}�0�vm~��&����!���z�BX@������e��?��VA>�Oh���_�b)Z^}��9e��&0�������I���'��a�o=�����"�|$epQ0�d������KӰtn���t���7�ߑ��GA��(;R��7+X���,	�U�iҮ��N��+.ԍJSc23k��d��I�kxq�/��/C�ۑ�& ���Qs��Pa��Fv[W�m1΁�J� ����P�j���E�ۡ�t���v��9�usڔ+��U�!:C�V�y#�?���T*끻�6$�4zWЦ�t�����N�j��G4�a�O?�-H)��
4n:�N����fP%��.g�*��X�r�ʌ�W�@V<�&�����=�_�ڱe������!gQs�\���Nvq6+��F:������d����+	_��x��=�P�;���P�an���� � t�!�8��$�O4Dʁq�g8�R+Y�j�ŗ�2��r>k� �bt\�k�s*\��|{�4��_�%=�A\�f��ؓ�
w�ȗ.32�������U5��w���c�5��hX?s1·>���@��
������l�V�>�&�����O5�	��yr؛)$#�5���R�9�V��URH��aCY�砮�Q�M*�~���B��؟j)�WݦVn��t���r�(Z��̋��wo���v�-ɖW�t͖(d���>���\Q"
a������KW!�p!�+�}౻�r�"���?�68Yq�sG�m;���~-�M��~�+A�گuۈR`��5��U����9,��@!�h��i�XՆ��N���n�R�~e��a���"��m���@���lצ~�5�T��H��X�[�����SA��d���9?zjBȶ�L�?T�HNz�00H����6�3ޑOt��N�hÞo��d�r	��1�g$%Ӝ�|@y�\���Hv��}��G���`�~��� �|�ޯr��-M�4Ԅ�IAH�k~m�]�H����;�Ŝin�:t�+l��9��ԹY�5/$�C:�)�s����pF<�M��$��ΈX�����2��h�֐~k3��"~r+��t�2ܨRc�'4b��H����,�Z�<��,��<��Hk�M6jn�j����*�)GN5�4�:+m�]"���5��RF���^@�A�ʺg�8�����x$���!.���7s/��14PU��[�5p+���|RX[��u7�6�;���Ѯ�� ��Ş�Y�����N��JR�B��2�ג;���}󽥇)6��vt��s{�?��]�d��(8�
�Y�Yӹ$ֳ'`�ˑV�2�"T��!cR�~Nݎ�qiVr��Y�8;J�.W.���țJ-^�5W�V>fҚ��c��8�=t�Z��ʄ�r�5T�����rP�B�*����z��n��tR�c���7���+(�,�#54j������� 47oW�0j���rcK�qY�h���y4(�G��2#��u4���L��7fyO�9^C���ܓ��%�:�f����UfmB=��J��}!�s��=�����a� |a�r������W8A��W2(@Z�ӝ(����4]AK�����}�0�����I�Ӫ+��+�k�w_�Q�ɒ���?#��>O�������dY�����*P�O�bd}��U���j7��r[�0d
[�3!��K�M��/�ā��
�D���K0A��K����5=JwE-�ߔ,��%t��Ѩ�g�f��=c�"�f|��|�~u�?\o�I�x&nơƙk�_�����xA_�B��znsy��k�{��f�ҋ�G�j����_ݬ��m�Z�S�9D]�@+� ?=���A�C��j�nQ��H#+wq>h{D���9���C>Izrx;��o,ˈK�����ѿ̸"�Zʙ��=h/����� �@%<�#���<VAMpi��7�$�@���WB���k]{������P}|��G���'*U��pY6����3�=!�� �m����h�s�T��)gZ��ٮ�$�2�hZd�Mi���Ԥ��-���L.>�%�3�χL��M	Ccc��$�k��}�R;����3I�?p�c,pK�G��X.�D�q�}��Ҡ�T/y|���A�9��"iZ$J��zV.��n�T��mߙ�a}�>��}�8���4�"�*��
.�A�8��r2�E`L���\���S�r�x����x�{��;閳�����6"r>���^�?jpn�xG�[PXB�Tԃ��$-l)W��9��1c��ԂJX	2:$����I����h�Λ^s�do�=֭��*�O+��@,m�&�P��I���7������H��� p���ВH�{ixt,:�B8�.�R����\�٥�A��.TX�:K,��D�3�W��� �T� ���dux�T��%�q������\�tw���k�#*����dh���u��zBy	w�gF�>�a���9@9�r!t���]Dm�ήl��W�AY��L0�w�?B���r\��QO���
ۚ����dң����D�����!q�Y*(9/��g�6�U�满UHD���lb���$�N�MK?�"kV��Ǯ��+��m(����
���O?��1D���j�CI���gϵ�w
#$ol��-(5��x�d'\�\k��W�qK���A��WMo���%����\��R��ԩ�l�ALkK�X/C^b��Rh��c�z0��χ�u����3Y�>�==�GYǱ��󾞉��;�LP�H�J$Nzt��]'!�b���Ǒ�NS���Q�	q*���S]��!�g$�~�^�ߌ�x����Iʖ�9		��G
��u�B?��dRN�]k+��E/��(/�����H Z3��k[�=s�wk�r-}zu�>�*�+e�	� �c��%)��c�<!����t�]~@^���3}sJ��]6�����.����:��1u�z�*�~�BAFk{���Q��+P����M�q(�#�-F;��-�4�1�~�w��C���o´��>m�l�?D}Ay�2�����jL=�r�_��V��霄���n����+{��H�ޱ2�l��y"j�I�vb�9(7D�7���A8 u._'o'Rn`�-oJ�D˼�X��55�`�ӆ/[�SL(gs���J���>��NE>�t�0��S.�d���2�[�,�|:em)�;o|4�G�K����������Yb�4�/�R�x�a�'���L����H��ɴ���K��ey�F2�����mR�R��X���8�m����=�H��[�Ԯ���I�It���G��5��ג�X��8��5Z�������X<G���?���Y�K��µ�ȑ��m�{�=�}�{��pl�� %P1�  6Na�#(	鬰�\�V*7�[�h����dT���)��I�*��p�����v���-W�}�Ҕe�:@u�6@H��Л�ʴV��������/��VqR���
��8Wǥ�$�������<1�P�f�Vj_��\��� &1�̓kA�C��_*ҺCh�OP�c7�	�����*'��5�ۤt�b�I���e�L�T���8�yrF����FȽP����dF�aͱ�8�D��};W�����5���7ˋZ���W��H�X$�0bPs��`��6ok���H� �����G��r�;H*6az �U� ��1O�.�nJ�F���1�cL҇���0d��.k�zuu�j{����8
o�2������A�.���f�"�Do)�ƈ.�H�-������Z���@�<�=�v
���+,����%����3bD�	,�-w�'h,o�Cb�tO��{a)��vr��7+�f��s�%�Β��"�Ru�Q`�=�����w3v&E����9h��'���B>��X���`R�DoA��'�)Yr�-,ˇ��17(�[��� g��v�XVN>��A<z��	ճ|aδ��o��6�N�=��m�<�=�u��A��kCsJ��W�D�-.DG��&��c<S$Ȍ�"�t-���G}��d_�N��G7Ө����||¤$��l	���3�h�b���,筷١�l���������j��
��?o'�k�&���'����T&�V�S��N����=��t�@���^{�m�c�m���w.O-��kKp�Ħ^rm'@���Le!0� �{���j��'�ݥƈ���&>[o#��+xj~� ��@Mb�4���6چ]���)gOp������i.�.��iyɮ9�&���Y��|�	ʇ��ʓ�m���w{7�PWC�m�)��U؂�I����zL�2c�2�dѫ/%l�Mۥ'_:/�qV��?MݠJ��H&����n���6d�8��հZ��Q��D�(��	E��i�/	%�����I��ӥp(�T1ۧy�FLS�T%�/p�T�Nuӥb�?��S���8ZW�8��؎y/O[C&��uȞs����+_�<��n=@As���*�᪵��s[d���?/� #�)�E�~.D��q�F���'�d�I�PRPvo���02ؿ�w/+r�Y����f��5�o�(+;d/�G$��m��';�B�����G�W�lI�I!���D��t�'�8����0�[.���ÏMv����D��U��0��3��c�<M���V7��|�-r��]����u&,U|�Z{^�0l�#ߎ���}����9�t1�
�vw.i�6bjO����N��ه�%]c��
�3�o5'�O���t~,�eֿ�"���� ��'P? �j�j��:�؊t]f9�)?�Q^%��Q:������b�b>G�:";�~IW��Pg���ka3+�sE�u����L��E(?$ �O���H�y#!@F��b����z4��P"�:2���]�N1e����r0*-%��9�L�w���>�>i�í�*�£�A�M��[����S���E�c��"��)A�7A,ޢ�ϝ��j���X�6��w�~����Ǯ�\��~s���.ɸ��B5P�]���8���$���c��
����B��Mm��?���n|O�Ew%�挑\b��L�!��7�8�^f_�9�?N�L���J����w�������S���qd�C���5|ܞ�.�C��	�AZ��nS@����5��XKf.{1�\o�(A����?��g�(��H4�Jp�g�92�"K��)3��IĞu(F�S1�����c-���-BQK��qz^��%�J��M*u�R����j�<��
D�VEJV�X�4�����j�jUu�B�ق&��ߞ6Si��R�0F
����}W+3}����y+��iÓ����C�äͼ�������C }A6
�bb�#�#]R�:�j�����=o��ݞ��4u,�L��� JX�*��u��	9�^���3����*^: ��	�?�մ#�i"P{���,oG�ƘP<�-�^ ��zS��M�Z[Z�����µ��)��**j3[�;�<V��p�>%�f��W�f$��U,�Hk�����D�$R�7C{:�FϺ��=���O{�㸜<��8g�8ZQ�6G��.�z8#��q��MS�F�M*4�IJ����.��
@+Tlh�����ʑ�<}Yx�[.��e�A�ŝY�-,m��˩!�H���	Z��xP���e���Ws,���$���`'�~����	�|�~����?~~_��9�s���a|&�˼>�E�aНzВC�7y���#�@��W��j��u�9����h�	jvG���x�$��r<}�/�ˀ�4�'K���U�j4���$z�a�FJF��̬��?U���G���.�P������&������em�;J@���"&��w��O,s���r��E[#�l<L�r߅1�AD���H�{�<��t9�>si�)yn-���x[���62����R�бB����?�W���K��B3���qK<������E����W��P>�j�B����)��T��gb���ba�G�A<�#�M@��ҡ�%����ju��`��Hk��;O�g;��T� ��Z�Cv�,C1=>(ΰ�ڀ1T��)^d��'��n�,|CP	���"&<ҕ����=+c��t��^k�Ds ��C����`84��;l��d�˿,ƺ���rщ��1w�Yȹ�2*�Q��������q���g�4���V���wy�el�+�2xT��I����.���Vj�e"�+��"�~=c����	��EN��F�}i��z# YnZ#o?��/���Xb�����,��ș_��<��$��G>W^������D�I�ظ�F����H� ��g��9x�x�W� ��W�J/7r{�u?O=Ժ�՟3��Xq|l┢����6�I��ef�*D�2*0sh�"��4-kT�v��YU���0xʨ�c�-�q�a�c�|[p�h��N]��6�3�DJr�ڜRI#�d��I�(NW���/P� %2[m�Q�D�ر�}t�帷bKa2(�pZWؒ��Cf�Jֽ�b�*�8}��#}�H�é��5"_�=E��^�����E���Sw�d��0呥��6���|ھ]Zo��יCW���p]i�?.�`�OB6:v��F�AS/�����;�3,'U�8Z{!�����+��M�c|�U�����x���jPA�޿�R��ن���B̞W��4���z�JFؼ��&j�)0aA��W��?�P���� �X��~��}ܤjMRK�Z~O��^��*��Rk��$g�T g
�]�=��v�fzP���6�"~�Rr��q���#�kW� �k7[�n��gCmS�]����rzԿ�v�����gP� ���-�^�|�a��򸰋� <��枵y����%�B������/�R��%���L��g�����_���b��~OK������X�vYll�4��>e���� U��V��iE�Ґ�8���YVH����X����L�Ħ��j9��%GB������n����ۀ����^�ūċ��9%��N>�_�tR`3
f�;u�Α�gT[o���\Z�W*��oVU��s��y���*��l��y���6ta.����_�m'/����xz5�Xc縷f����O[W5o���~�Y�K�f��,ga���،����<#�:\�.nwE)�$�*�/��
$L���������-ŧN��QL�� O����O��,HM_�mT!e+j���-�]���	�.�C�
_�k��l��	e��XZ-b2$2"�S��՘	��^F���͌Q�4�����Y�:�̰��\Á5)�aG�H�2�ލ��3�\�\t*ʚ�b����V��M�Y�8��8Eq�ֳ@D��P�u�)K�e���
/oj�\:a~�6B}?n��c��;|"c��V�ǀt�%G�Q�+�Q"Y��g����0�۲�T�D���EYaߤ�Q)>�۞-��R��	�W��cK"�L迓���̳+��Z��6c���8aF�<:���G):k��4;�R8nj�+ t� ���x6������ǖ��-���xNן��{'o���t���ʱk��i�U����A0l;
�cXĸhP�<d��dK-�* �GD���CITW�{����p5<���o�\�����7y% ��͓y4��<U�y�@.��U3�#s��K�%��	Mvt�X�BZ�.x4��C/q(��������J��~O�]ʦ��0�^l_V̜��g>-�@�ɦ�x�Ѥ�2�9\��;�?f��T�dy�������|�]^B[.��Z�ݾ�q Z�,�`��C�E ҁ�'�h�%�$����!�vo�<�����Ŋ��bX|X�
W��y��F����o��8��i�Z��0?^�v��(Z�c�����o	���F�U�ն�J�@�(�����"�*��m���%�x�ʌlG���˫@�]��T*�,�l�/5I)o��	w�'�t/�����������(a�,���a=#!�!yE�JC�A�n�D,P���	j4�
\���4T� �<ƛ;@�-�u���_h�|C�ӓ����Twn�ĥg���" �1����64�M%S��ItG������Y������ْw��l�S��1?�N9��L}�Y�+�^�����m�i1�,��:|Vy�r+�LP6��%�q��p��� �OB�P�9p�u���J_�\$w]*숙�f����x�eb�EZ'F����,Pw��id�A����k�BJT���ǰ�-k)E3b�)
rF@W�ҕݛ�ҋ�y�W2�`�-��w��|��3jzG����˅'�^�~�zSJn��5���in�8Ƹ�k�	*@������8�"����1&��� ���ح�}���T?���Sm�>��n�,�lVr���u���Lh�>�8T�p���l�.��B�u2�6���&���j�i�Y��:�\(�
��4&��R�a'����9���~���-�
��l������O,���XSv�@(�I�,:L�ݷ�6�2Z�w�p�R3(�\��~_��p�r-���tX�ߵ�T[�na�T7f�H��:����e	����mW��H�u��E&��  jj�,j�S�꘻�C�})j�*Wy.��Kψ�.�z�j�=/��l՝�<C�����"���)��uy-�����������Ɂ�幙X�j����@��]�#R���[�#���P�L�D
�/%|sؖӼ�h�y3gG�%yL��x��9>zpsc�Ҙ�B9+�gY�B��n��AV	���9�d�T��Ǣҳ�y%4��L��c��(%vS�k��x�>:�=S�6c	&��%��_I5�h�/��GiQ��:U���y|�>��r����[=1��}2����������&d7��&���:��=��9�&�<�Y��oψ51�7n�H��x��o�7m�����ޢk�T���"-c'�a�u��S���OŦ�apeP>��])���7�Yx����[���s�����e�ї��Q��$S?:�{-Mr�a��{6�JX��-+�Y�l$�V踬�Ԕsq*P���=�^���37����̂��l�.�lV�&<��7�Treo���e�He���`�2ج_!��
�Y̐kp��r����[��aj�ǢO�W�˾J�Z���=�Qv�Y��u6c�N"6�2ڐ���q��ڭ�)���b����긌������^x6�͜>tC
��q����)��9)�����ٜA=��U�;��y��i/��a{5*��^�r�R��,��qjٷ����� �^�g"���md� }�� v�6V�;Ox�"�7�����LO��sO
$C�}��V�"��]K�萋=��v\x�����-����2!W2	o~穔�jd�UD���&���dZ'�r���=��A��s�����蛤9�;Ý�9��p�,�+Xޜ�TsE��H�{����ܲ��@o#j��v6:���g��f�p.�.5,s��L�
���O��D��(��	������ F�h[`@4�rF]���os��2PY��;��yv8��3�X��*��U����O[K�/ZkFVq��j�PE��K[櫝�𗚸�k/.�R�(���x��8,��;1�7f���J����%8#�_��/��o�q�`��P�;��|a)�/�'�q���w�������G�����7#�Xp�y~Z�B- )�,���<�o
�i
}WB^.8�m��*�'�f5W�������P��f�y2�"t�qB��(�J}��Z\�&Nkq ��:��tnE��z���a{��~�(�/��Z��B2���;j�P�f����'s+������t�+����|D*��'p#\�H�� es���V���'�--ީs�V;�x��?D�Y?qR��}	$��ڎ�V���c���V�0�w��0�-�w�'<hY��,��t0�: t��	�F��-ac+��U�e6	��m���?3]�<��L���l�w�L!ejr�F�0�!�?�x���/VY��ٌ]l�wx�T��ts����]:ZtqŻ�W;驣`��;��z�a��4&�.�6
%�n�(������48)Wts�v �⯗�j��{P�L��i�{Vk9D>4���<��2�t(C���mO�	t�����+QUm3Kc#ټ���.�
��i�\YAy:I��}.�`�A�h��j��jC�Sj�!�<�m��oK�_���j��ډ�<7�҈ݭ9�{#�H&�������@�.X�C�՜�����<����v��K���胉�J����2Ua3�x���t���Z���A6���,) 5�\6-�����旨r���|�z�4xI<��5�h�]�H�ӏ�����n�s�_��7i��AS�[���}�jgZ�Et64��N�m���v���SN�̲�3�1H��I�_<\������*g*��U_@��k��*���D��k��j�|��>ۥR�������F\���.��M���LT��]3L��slK9�\�+�`�.�2n67MR� �e��FG�s9�'n���������FYI;]�e�s�[g�e���(ϲ�����H��kZ 2ݐ��ӽ��f��sq�^l�F^�=�9ʻ��K@�.��|]~Ioy!Ţ��O���,`��X�t�d����=7u�]_�wܶ�i���,�E4||�>�gݶ���&��X�ܸ2̺��d��3A5<�F<͑�h��$�M9���uS7.J]!��:����9�Ё�k�әxdӄ ����{d��E��^�2�j^A��\�>
�Q%�|.$*r�&}2{(���� .��9	eqxv�P�h�0ç�Q�"�t}��grI@[��$t#�K�
��Me:�W�q%7�էD�r�3 ��8��S��X��AY+}5�sk��"�63���:���w�˷'vy40�h��Z�*���H�T����[�2g6��Ea:M���J"r�а"h�(�z�'�L
���Q���V�Y������ܻB ����z�.}��"��,2�!'����|�MwrZG��̃��FE�Py3�����|I������{{��ix�lI'��j����7R�f��]�H��� Ej���)��ޠ�ǁ�:�8h�/�58b	F(al�NAy(�s�B=�_j�E�p�2hn�Z܀�wI�� s�0��M3;-�^�l\}�c�ܑ��	�q�TƖ�yXx�L�~��Z.�w�;��L��r��2?�r�_��c�����x+V�`�� �tb�>��=�d�ͤ[��I��F ��)�	�'�;��E#U��J���@b�z�E���P�+_�z&"��%�3��O����'';φ�?�<�"ˊ��h���H����x�K��̾�|N�9�D���<koY��R��r+m7�|1Eq�qTM�R%����;@*FY$�{ �xRж�qľw�UY���(�����,7e��9��9��لe~Eb���S5�f�)G<F
��D0K�+���[B�!Ѷ'U�I};X��h�P:�JS�ȀO���5�l�ɖ�c2��2/[j��9�l%CSM���j��|ߪ`��i#�p���V[��S�U�v�hc�Z��#����ް�o\��a��Su{̬2'P&�~$$���!����������K��x�p%G;̰���z�UN���Þ�'�����)1^��V���ph�XtB�C�$���k��}�"o�Ʋ(d�NT@gϕ3��������t����v;�|K��H�lJm�v�."H�c�0�I'��c[�ܨ��+��ӆuy�x���>|
���＆d�DTx��n�J�/����R�h\�c�Pvף��#n��+s:ݙC@V\�OI���<���S�&!�j�%�������]�[V>�3�޵D#󖖁K����#�"�w'~� �M:��Cq�k���E��~Q����P.e^�&[2f��Yj�(�Q�e��^v^7�jEu�3���ZEᴡ�h�E�`���}$��Y~)[g�ew�<��AL!GO�>#n�*�ރ�ъ
���Pi(w���s
�u��S�w#����N-���.r'޷a�q�|$����jl�W�
�
�^���V@ǵdȜr�����}��� E�q��6���!�D�����2#jGgfi:���z=��#˯���8^��蛴b�����Κx��n؁V���.n�ðηzoI�������xiW���%��5�Q|�K<A��4p��c�A'��m�/��$�ߕY�
�"��ŚcQ��9�B���+�q#-8�y4\�|#�ˣNKy�k����H�x0���i�ɢ9��c~k�\
DՍj���`�����T4���os�׿'/����㽤U���y�o�k��X���$��PT�@��G���F˨&����p$n��LUr��<�l�� ��EfVn*�yv\�x����brK���x�4�����V��6[�\Dg ��=��ƅ��q�ҧ|��jԥq۫փ�:!1�H7�Q�hK$����梣A�F�s��q�G�F�p���X2Թ�{U�v� �S��?ףe+nI's��7a��m�~����h�}�1v�h�O�W�kp��"�Ҿ
=a ���Q�7���Ԁëӷ3}9h�NV��f�m��}�c!p�5�j�?�w� ��0��a4�b?��wDb�v�Ȓ��M�sٗn֬{�+����z�S:�Iɡ�*q�
�,Rp�������)�=�J3eN������#�8�&��`�(����ʒlE����=v�yp���q��?���}�H'=K����:`�[��l]�p<�~��ē31D%����"���a�txl񒎴���x�J+�FP��_I#�����b/��5���Bİ���z; �_k�y�æ``hH6���h��z���`3<_5#�������Tc���GA�-�H��}�:Y>� �ԃ"�0xZ����
�y-���(��Z�֗�����0G��Q[�����E�tBN'�t2s��J}Մ�=�"BJωA8�U��������g�'<�]<Ay� OUY�M(`��`~K����@�p�"�u������EX�:!kvsa� �x<]-�Q��s84�JO9��\�6��̓Rr��32RXb�&ć��U�ώ�3��о��ۭr��dL��[vcY�v�_�|�ؤ�)��`��#˵@�T^��{�q���U�d&w�px=2���N\��j"<�U�"qZS��s���M�e�D�A���'νZ�up�"����gE�zuΰj�� ����.���I�J�����@Rb���pC����B�M1����9I8�m{q�j|�t��̤0�U������|@����a_�s�Mn:�D��,w�*ȋ�h�ɝ:����|��WYu2I����vq���jrF")��D ���(w�S�y�gdRި\�	�H �h:�p�W��QӁc��f5KJ���g;�KpL�Z��?E�>�{E�Y�osf�2>i��D<��40c�&�����@��I�q`��0V�T��~��Q��#�O������^��Ȝ��_©Ϣ_f�� L�<�R�ScM/û��[81f(/���,�YԂ�����@�*��Y��hј�~7�/5ok}�z n	-��߮����V��ݏ��0/�$D�Ć|2H�%�D_�M�<���6~Ϭv�?�>�C�4Axc��«�| �N 9[+��Y�#?��$�P,�6Tj̓]��k|4y��W#�x4tl��D&�����)vh�fiR�2T�f��ʞ"�i	bݿO�~7�.�Q(�H�BtG�S5�pN˭\c�,ƶ�BfS��؟G���o�y�8tv	sk���3h-}�.��c�*�	��L]sYg3J;Ԑ१�Ƅy�u�;���?G���6n?��y	����V��r�C7}v��(�ޙ��+��-҅�s� ��d"L�g��q~;�3��3]�|����6��~����.��z��]���o�-�����O#��C\Q�����-�$�����k=)�v���eusϛ`Y�,��9��SɄ������Z��4;��g���lо/r6\�a���� ��4�v
t@�$P�1$>g�sMy��=���Y�>�}�����Xvv�^*te?HEb!'�(���K�╌U�[yݙ���Ӷ�.�5^}*^E��t�|�"��\8-�ox��5�S��� ��3���6����,�%�|�W�a�N٦m+���s��#k������ �����SG�^,{�c�X�n�ӓG��]��?0�xb���E��_�]?�lW&c���ȽzUQ�޿�N�׌."�NC�C�"�ޅm���q��M0�(���X`b�fE�0� �yv~�"��;�#��1X�:S��9xhJybJ����~�� G���f,y���Я���]�9L'}�r�vADCocQ�&�?+	D�CD�3�����Z�zp,e�R� u,M[��f�5�>؁郯t0�
�RMu��2�"Me�<��	��8�U2��2"y��X��{�.w/�)�Č\����/��`y�q-�"r�L�DF��>��/�&D�'���\Sp"�����o�1��wӣ XKm�RjCgVP�"�t1��L�<d$/&p����X@v����`8{pJ0��F�T�����>��3/�nY!���:��,x$*F�A�@U�D!B	�:u�1���؁SJ�N�N��$�Smw���Dz��~��6j5�Ȯ�+>��N��8)�瘈�(��Kx��WL�o ��#MGi^(O�[���<�N�
��q6���5��Q�����ٍ;��� �:���kf�$k{R�y��o/ƃ�l�5s�q�y ��}�x�A��NI��g�ь�b��s�_�����-{�?G|������w�0Yϼoxk��������7��o�M|����KB&C*�j��m��z}����]E�ϋ�[��7?%��  <��z5�~y�hKȩ�!�q����Ĩ�`"O =&�*w{R���� X�v�l�TM)��d�KQg���G��X:ؤ|עJ��������I�_��P%��K�`S��D)x*F�Q¢����=g �m�YX�;������� koSad>�K�o���>�>OT�ʙR�욥t)���yl-~��+���l�(�N��H9w:�{!��d���<�ju�0��@>�� q�L즑�9lZb�%�+�D,���֘J�pEY�D��B�� 8�� Yjp]u$�B��-l8�}zܷd�k�ZEń��K<����s��S�����"����8J���Glߋ5ń�������C!���㶨���}���8B�r��`ғ�R�u�`JK:����~ӽxpʁd���t���R���<������C
�-�$F�>8#̂P��@s�R/j�pzR|�H�"(� ��>���e����p�4@<>}u;�a�7�M)Њ�;���N��!{]q�:�����|X<MYIm��Mx��s�Q��k���fII�?�/H�L�c>rv���Kg\���Zx	�����
f��Bi9%�m�op0KXǆU��C��O��[ �~�-��
Ô{K^s8"L�2-U��H�D�h:b\�/q���g޷���Ѱ���� �'������F�H�aΓ٧�@�u՞������ս�D<鿇�[�f��Z4�H��&>4�ط:���3+�	}�
��Җ^#~�E$�����]llk]��],4Y�dƐS�I&�z�n.;����8��5%.��C�3Xp5Ia�������1�p�*rF�D�BҜ���f����jq���L_H�+���o��p�����b;��u�O沮}J�!�r=T�rk1�f��syO�ܚ~��nw�¼�T�rҟ�}28�=�9�XA��G �2�DѬkO��0ƣQ.�Yw���j�TI��=oJ%�O_6-5y�ty�	�%�t�DҬ@r�0��R��+�p>�%���q&���T؍-s�8�+)�u�ϺtR��#f?*�ZӪ��|7�(�S�$��9J�?օ�q�ʨ�o��z����2qeE*��U����t1�M�V����R�z��oX��L�	=�)�Jv��6E�
������*_Р�2j�����8��m��FD�-� �4U�
���o Hu���5�k4�FĆ�!�T�~��C>έ,�2�v�TŽ��Z
��o�k�+��J�������p�����vsQ�g��h��;؇���C�0�f����:��PYJ��LK �s�?x��<@�"e�#)B��1�4��o�V����fV�����i�Ӫ��ǒ�9Dy�-�
Ȁ�>����<�����|���>���x���r��Ձ=�=�f�]!X;�R���ɟ4�FMh�Zi�B.��'���Y_e`�jk ��ր��3���$��%�#����6��L촒Q�;'@L�k�ꂌ�^��k3�^w�]k���!O��;M #���|��Ir�y,���
����m�%�U�����3_�2��v���tj*�;' 
������Od吇���������� 4����%�w���t��%�C�Z�b ��	�oJ7K���E�~�H�R?H�ka]��Lzz�_������}��Y�;z��@A���Ԩͥ��u��Mh(�����&U�bp,OK�4킿T<��7����Q ��-��%nѻ<{#P�k8j\�T�D*���,��łㇲ䃦�ϋ4����b6]�Kܻ<�xbZ�J�[v�yUm*C����:���<5Ar,�8�)�Bv�� �s���.�58�]^���=��I�V-�A��ߐ�K��u�V�����-�p�P�nJ,�?���S���$1�'M������R�����7'�Ϡ3��1����(?��&�'��%�!���P���7�9Q�[�D�hUWc������$ao�j���>�7S����ŉ��"R��X$���0��3�T��u���s��_�Jh9�;������͹�m����|T�X��[�����9��D�M��A�����ڧ��Q-	�b�q}�k��`�V��Husi�9�g|�j�s����4AR}���h�Z�u-��ӫѮ:ͺˑ����aH?��v��Y��|x���@����pA��H0�q����e��,��lm�k\d���������7����Y�|�W�h#����fh�O���.���װ��EAx7��5�)��u�[�7��!w��N�e9�g�^��d���m�+�0�=���\{��{՛��`mr��ʵ���V�����������1�u+ZδGˋ�V���ػI�Ĉ�6�?Ĕ���	-��O��Ѵ5��S���ѱ��g{�c�N_�M�#7�ըT���_���!��3��ּ`�<e��}�2��YS�����!��ǔn7��F��f�h�L���>��GP&�	T��L'U�*��Y����9ę��E`�`.�M]ѩO�X3$8皿j�#j�L�aT�B{4����w���0d�	#C����Tn�����k���iv�����ء����ă���6��b�Д�9} 6f�^��;���Vv&�[�\���g%�W;�>ײ5����M�������0k��Wn����Ÿ S���d�/���y d뵛�o�sJ��'�6�v�H�u6���TE��j�h��;�L�� ��9��Z�b!0i�z�u�;l{��3"|��*�z��b|�ǒKs����Y�DgNWt�#E#�Mء^��i���ʷ4E���0F�th�'�^p��\���TP����Q���J(�N+��k\�/���P���^WO�A,`g��>>|@`�4L5�//6a��ҋ{�y��%#&^-ã�A%�[�i-ւ���A��П�M��:EP�S(D��`���P@��\�Y�L����"b5�����G���9��q��#���$�>�̎�W�a�b3�u��x!H�U��Lq9�|�;s�+	�.Q�/81#��0Ќ���~V���B�	(��c�/2��ۥ����4x��nM���ʪU̔(=�~�X��qYr��JQݖ�ċ\�;+�M)4�涞�k��0~��]���h]l�n$�^;wa�w��Xtl�G	�,�"����oP
�]<�Du]~=�&�Ow���洴&�ܻ"d��lob��:��}a�7�^�^$.2�2���-	�6�.��~0���c�l6[�E;W��U���w��p���3���@T!���}Bx۩T�yaז�л?�M�֮ID�#�'��F=?:���gC0T3u�-�f\E�m�"G-t��l��o\.'>d�*Ƒ������ n��Et���A ��[�h��m+���<�fъ�(��@�eu��S���YI������{�$͈ƫ�I�g1�$h���'ВG���"z3)�*~��v�����	�K��=��J�i<Ń��.��1�k�C���)�=1�7]Ȱz���7�n��p�bi�Z<>�,���A�`=w�)�)���+�2�Y��:&�5GD06�8�5������| �S������%�R�o�+^kR�%�Vs0ۋz�ؕ,��P(��&��n��!/�|s]Ww�\O�ֱ]&w�,����F�z�a��ۣ[�ŮJ����ꔳ�0�\��y��e�~�	G��6t���v�]@sJ�K.��)<B�����^ď��AF���O����N�[L�|��e��,�κՇ��Jc>F�*wqٟ�Q�ζ]m��YBÏsƓBG.w��ث ?]�v���E�
��*}Qt_i��XTC���<!I���fp����1u�j�_�g�Hm�`h��I����u�"F����z`k����IZ�\���<ҧ>{�û7=��33�z�wY!X`Ǩ��X�/�w�oH�0��uų�Ec���Ӷ��s����j����ze�V��:�m2��ͭ��H�D��[z
���Y�{J�6YkԪ~�a�r\S�h���*
>b h�R����t/��B:}�k��&s�T�� {���%P��v&������1�T�)��r�t��l�Yޮ'�?��0���e���^[ۙ��r=�Rp���'͢��E���G�~ �(��{������Uڗ8�������*Z'f�g{*[��N�9�w|ly�̇�/��
?]��ד:�Pfk��Щ��2���Oy������tyf�Ů�1��ɳ�E�;�=)��n�Z��_.�I�n�YZ�J��
��W�m;=�)��)w|Z@��p=��^'��r��U�4�.=�����H�s>����9-�W�Z���0W\�|���x��.���Ӗc�h}���#���9+0Y�$����޵�U�6�cp�����;�R>�H
�v�G�8/gd��!���ҧ=X˼w+�pBf���i�T�<e�	Y���wF�Wf�6�bN�V��+�*����S+@yN�c?�L���T�R��)���=�Rh�ÄnȾ�10�47b���#|c�ES.��9����u3�ox���3#��I�T?���N����6�6ލ[5���-z�y�'J��O�v�1�����Ǭ}�#��/���A��v�p)��#yy���u'���5�lZ�����c��!Dz�9�a��e���z�8��T�O�����2�m�r�o�e����҈6����t�ň�ٚӄ��n����R�v1�A�jܺ�[�l�v��4�ǻbf�z5�J.��
�-��*�/�g�~�����0�i�o)R*����9ij�t<7V���7I%i��C� ��D��_�YZ�kg{t��\#�uM4Ha�\����\������]DƙQ�&���3 w�hX?0KD����64������>?��`3S���0�|�Hn+��b�.�N0~,%؀��lt�ޡ&���S���sS[���}D�0li,�t��'�������zz���Q��<+O������p��!ţ"s�| ����}*�@��bK�J^�΂ڊ�M&��>�/��ϥ�}I�����g)��/r�W"p�E�}ޤ��9��@CF�������RI_J�
7�t"��Yf��ҡ��G��	���޵��ۍ�@�4��C�G=scA��d�V-ڳ�Z��[�rT&��_]N0�׎�"����Z�[�R})_�ٔ+�Ha���;v/�&��٧f�#v��6j��XZ�}���R�>�$DR���_�x�Kww.~��8# �@v܂{
w�
#,�6Ͼ���]������?gřb�s����ڗ2^��5���q���,L9�8��:[���*��8��r���J�QĞ���1�w\���r�����k�gZ�N���x%wmNB*V-m��ԭ�S0pP�����S>绺{�&dCTσ@���<˒��׎�������re�ȧ�g��x�Б��4���ȫ�#~�_Q�97���a�F��+��Z��%���E��&�����#�,�hpi��h�����a"F�l��J�;���F��V�� ���YV�˰_\��(R!�o����SE��0�R�,h��7�������f��:��<�y�����>����ɴ���U�jiKl=��}�b���H��/�]p�",N�X7P\��U�H#FG�l'A�����Qi��[m){����]�c��M�ܳ�,4����<�x��Iy&^��U��!D�ߎ���Q�p�}p�t�t�V��i�r�Vgq`Nן�dC���6.OҴ ���c������ZFp�uD}�#F5�,,�ݟ��Iik���P%W���P"I-�C�����R��5^�Mt��Ҝ�P��p��?��JM�[WNSJ��C+��ov�P)	���]���(<�K�Є�e ���ϒ�@GGr< ��}���������X�x �I�/�D�{q��p���C��΃���F=#,�<3��ןo��{��G��BrǏ��k��h"����H����W���.�J9>jle��c�$���P�j�ZI�l�~Ɗ>�&�0�[��14yO�%�;��������I�8���'�U֠�V�Ǡ:;��ȓ͊�fn	�`c��Vl6�b*�V�v���v���� H�� 8��hOP�|U\tmj�[�`�_r�t�uT�14�%T@�*�7ʢD.����T�b�ĥ��ݦ�A�L�ZZ��_��z*ِ�+�B\t�*�0�.oc�L d��,��QMC��Ɣ%!�j��x ���UX�U6Lbid��x��3�̧�AA(+�s��*�.�E�%s]c��\�Zsw�y�����	��t'�N�9�*1����'a2��K�0kP�(�}g\Qbg�K���*"�5!kcm��O�d����x9_��D�/O~�tZ2�:��t���V���5|䬪�W��;��0O?��)��靛a���b��ҹtj���lwц��gy�=��4���(��[N���<}0�*MO����B���%���C�`[� Ύ6>Ql��\�G8��v��� Rc%H�Z������ZI"��y;$p�F襔C���	 GB���[�f0Z�LF�Z�j-����i�X	���*��zD 5��414��r���K�;��<��
�$�π�-�ijJs�ҁ-���V@���_OG@K�8UKJLb3�>�����x�|>p�����_2M�
� �+GC���h�+yV�;��)��),�5����ADoO�5S����l̙x��:��h��6��6���[Ja��T�'<�H��g9�ؐF�#*P���+~8u�i7\M�d�L~˴�wpWd_�@�[D�I���d��4�"�Z�C�TH�=(����/����c|�݁1+&�̍����y���gB�|g������0�b���k3�V|� ����s�_TgHWK/#�2�{��\�$l�Ϥ
m��Ǣ����}pCG�YQk!�G��7�7|.��h�Z�.�e�Uq�V��:�B<�|A%x����VM��)�Y*.������O�s���t� `��@*c$<0�)�x ���$3��)I�~$zk	��CU�@���q�ojj`�k���g�pىa����s� ��m�q/6I'��n���H_�S��ý�lk�����q����r)��#;0��$��9�i����5�p���6��������ե,����r�;=���N�H)��N�?s�|����5_a`�����c5.wu������f|$B\�>���!I�/��4
��w��á"�n�F��u�E[A^^Gp���������*-�;ɾ3�%xz��z�"�	VҲ�_�c'�dj����8�]iY,V�ހ
��D
"��s�>�$��QМ��a^,���ȮS����@�7�|�3����݅H�|l���:[|>MV�B#�谖o�5`�z��X��@�	����Nݜql$EOF������qV�炜��0J𐎯��҆.�nN���w	N����7�Ą��o�㼞Z�s���i�)�K\�')��r���Ӟ��{瓪A1w$���������ߎ��Dt
4݉�w����S�LC\�
_-[[��(�˔I5	9�
T��V���E���}����m���MavK����<�y��H�]Ǒ!j]��#�4�w_2q��j�]|0� �H�\�7�bH(n��T��w..�,��(�CC��`�:�JjZ��a�S ���q�����U�84��F��H�`~T|9��x͡?�B@Wzp�SV��u�]��a�)Iw��]}MU�L����/��$~Z�R�}�,���tK�t�]
t#L�
�p�0�����(�<��쌬�6uW�Ҙ&<"�#v{���b��Z��I2O���b�~�'���hf����]���»�6�RӨ������W/�-t��w���d�����}z��r^��20�/�9�pP�3��V"�,�r�����CF��!b�0�r�����^H3��zEG}uV�8w��a���V�O��t1�wuA�I�/lЧ�e׼;O���h����Y1��P)v�����F+9�/���E�>f�-���2�����_=�P�� �o�)��g���}�%���4��E��V����y�asy����Î3�\ �@����.sz.`�ܑ�w�Oу#�b��������:�F\N��w垝�k��Υ�*�j���E�,m���+�x�"���ƣ�K|G:j��&K��V\��'�:�_�	��K�l'�������?7��l�~E�W�F�_�,�������˙~�G�j�4@A�|�|����3b�S�j�6�<ԙQ�VX*��>���,_uB��$���qYz�Pk�)��l�\N_Ş�>��8F"���e$��ߛm�JD���ؒ͌�t��L��(��� ����U&�lb���L9E���L#D�����t�z���G8Tq�a�8T+�`.�nF��$~+?�4�O܃�킾�	�ܵp}�h����� �����8�r���g҉�H�
 �q�,�`���d8��T��Ux�h'����d�8�������s�@BV����ݱT$����M8o�U#"uGz�Dz�-���+�5�ʬxr�e�������:����o�Mn�3B /���yd�߯�$H�0��FPa��̅�6lB��PZ����p$����a�\�	���`�ǵ+�|&hP�=/@}��|ů��z��Q�]�em�|��y��G�3�|]Ӌ
�2���x�n�sGU
8q�k�u/W�Z�p��3ar*���e#w(В�MRT��?!�%M�&,^Ʊ�G
� �*��Ded�:�h~b��5'���D/��b�q���q�!�g6������:E��ڰ]I�D���t���&
�.Ə*^8	��M�9��E��Ei^��n��������Yݐ�u9;"��z'�V���	Qu�{�E^�������f���FW�Z4I;�jwֹ�T���zgƾQp+
��S���'W��ƹ�w[a?:���O�ފ M���̎�~T����]��B1���0}d|��`C�&�k�e�Dg�z�WZ�~�"�Hg��	����ýփ͓��-���-hݹyP&l����7�;�7o�L�{�SSI�1�ku)��҈D%��Dɕ޳���ځY�,t��;���u&.ߚ2sm���#��W��2~������h8.{'�t��հ�wR�O��"��[#i�n��!kN"Ċtf��L����,�k�ܥ���������eLr��Xb���ɪb�n�����:����
�X�� ���cKz>�.��V[�J�&�oa~����wt_{t�p["�fX�0���j�jäv�N!��*3Xɨ���W%h�,��&_B}#x+��yfk��:�{yD�������uR7[ɉ�
'�yxI� Ih�3!�X��Р��C`� ����6;=<Ȉ���/́� f�z����W�e�xm�/�ބ\�`ya��S���;���)B�ȥ�n���̼;w���D@S�\aIl�<C�:c�J"C^���gg���;O
�Д�{p����öIg�L���;���ߙ�����#_B]BvH�;B����D��C�,��p
�!���|8n�5��!���t�d�-�������A Q��X 3���âΡpQ������6�,6%��r�q�鍛pmˑz7�`��~b��F�w���>Hq�� Z�~Z����KEf�|���zI�8�q�Ix�z���u-�Hv��|�Q� ,�����tΪ��
��3�sV�661���,�ZI�-�'"��� ԝ[4;v��J��Ã�k�Q$����G�}eOY4����d�/���و���K��}��q�q�.����2��	RX>��I��fgJ��_ne9�>����j�.��ק[���sq��?1�L�
�U����M�.q��\u�N�mnF^�VU���ڱ�7�C�Ȫ%����>4�>y.�Cֺn�u�b�\+��I��}�x�	rqy�׮-���,�]'�h�����/��4d��ۉj&v��2�ŕlu�\�H���|S��Gn�6��jdx����w��w�*ُ.}�I��覧L.W�@�X��5�7�B��;@'?i��K+<-Ϳ�:�U���I���W���k��Yi-�'/c��u�m@����+��+0 Hv<���	�����5��X��.�t_��ZZm������Zs�k�.�G��{�~|5�M������H�2�����炭ݮ$�hNR� � �P_�y�V��iL��k����y.��!�/xvS��M�ӥ��˻u�� ��Ӽ�8���^E��q�4�Ȥ���8ί����x��[nW�ɰҼU��Ɓ�7�3ȅn����e8�+��Z�Wv�U���+���+6��%����Mj�U��*����A�^VRFHT��q��GZ��v8�7��`놙��Ɇ ��Jw�Ah �@��)��-9�Ŗw��oi�&ڢ=hy�����&�8�c�]�.��C�d�L�o�(�q���h�N���/qA��bmB/Z��佗{����=Z�V���'�i����hi�0*�>�Հ�']��7"��_�|��^�1�u���p̓s�s����@�Ñ�N"����SC��W G�q*���G�����R��2����^G[�-�����9p��Ţ}�K$	h����Zӟ�_�J� �[��A���]���OZ��3�i�H��jq��i�$�o"�O7��/���/� �\e�������$��5E>�v~���{��§��ml� ���J��r�fT�!|�M���}o�~�����b��c���Iȯ�j���7��2�NԦ�=<	p,�]Q`����_U?o�������J�686�][�奄��w�f^U<EC��d�h�l�l���x孥�`F����hb���!�D�䜧*�����I�JP���I`��N�xh�Q&E�v�B8;{H��KN����N�cmX�|̸��
�(w�i�˗�y�0�5�G�r�D��d"��p��#"�X{-B	����nA���(��z�W�K���.�)�1B]f�
�M��ͣo�0��u�NP�O���~���sxw��G�Uw�����o~�s0��d���J�ƚ�Q�E���.�6{�@V��q�:���+z���U�gup��}��m���l�{5Nk6�	f�+�晫k΍��%��+&R�š���EY����%�_M��M�*DZ����$��/�+�Xx�#��q�Z��D�30�m��Loߖ�Y��ۓ��l��P��ADĴ�S���:�c�N�y�]i�5T��d�,<p��uǓt�w�2R�M
��X��S8���2��}	���5��z��2)%�G�����\���b< r���a�m��M�ĸ3p.�^d���gȯ�Y�B�w�c�^�
=�X�U�)/�Q ��+(!��6��m���B�W�x!��f���P&��t�����v$������PҶ�8��QK>3V�oG�V2'�x
IS� 0c���.7�w��Y�|�����a�=/����V�i�P"j�Ғ�6� �ٌ,?R���i-2��kU� ���N�y���E+:ypmCKt)xbq�>�W�%�l!P�6GV]I��^&T�I���:�7nS$�ٓ_*nw8J�@P� ��G�/ە��IC|N����q���ISOb1�qҫ��Nq��}�18�S/��]i�xo:�z�_oR?�1+*<l�Eʝ«s��1��}�o抛8����k��.��g�1�nU�y��b1�=�(g�0265�����D��q�L�r �����_u�b#Y!=������ f0��5w��5>���e^2m>xQ�^���d� 3��$0������(kCv=�(�Q�h��kL�뵢=D!ET��=\�U}���_�qf~/R������w+�HV}��H��-r��ENҽ���T(����\\?LJb�NFr�4B��ς�(A��uw|�Ȅ&C~�&f��$���P?Bo����<N��"#?@r���\�������O�h*w��/V�V	�oܑ6"���	�mb�6Y'd�bo:6��w��Q��кZ��wMD�>3s����r.��td4~�
�hޢ@hY��LM�(�k��qx��s��k��?�Y�/��F��,��Ad�3/-��4��ip�z�S+����ݯ&s�TǸ�SZ��|rTv��N�|f$��h�o�m�!Co��&��}��rl��b�mg��:�ngKєJ5��ZE�_�t��G�i�?�zyT���'�GR,�	;PMq��ZǸ�nT������-���@�<h��n�!��28�i��o�L'���&�m2B-�YG���oDRsV��<*6����ur(ۺ*��чJ��hR���'�I���'���Ez}u�o]B�������ˏ�ʝ�W(�~�r,���ԝ����G�f��)y�I��|�{g�#|]�sk%�m"���5,x��i�~N��D���(�(b�yju�#�*�Tؗ��#�(:���G�,��o��aK��l�mw��;
R:<p��2kk�p��|��C>�55ь�w�^v�1�\i-�����Lދ~$�16g�\j|�\w,����S��2�5���O�)f�n~Q����������!�Q�p5�K�k�E��'z���D��\ �V ��^������*���!���ß7t
�RTQ��Jm�`��u�c��4�4�~r��ڽߚW�d��K�+)\��yAQWS񱜃�����:� v�*�o�=�e^�I������
R�/�K��F�:(���ş���i�d�OK��0�R�`\����-�nԆ��@�����)�����t r�Q�	ʛ�A\rX��9^wo���& ��Gב�Uw�^q�R���Mۙ�+���A�A��zjnr>����%��u�V�J�V���|~�XG�ٻ��ఏ��*��ێ'ha�t��y���AQ��$U{1�I����������]�΄ZT�P򜺓�x��N�FOTA�g�L���J���h���r �u򗥞_�m����f:�եn	�ߤ���&[z�b@�����Gw�8�����k1kqh!�K'�8���$�����4��Oz_(H�^��`C"�P�0wG�W[�S���t�('�𰭛c^�ws��C[�4H�}޿�����4��(������+?:��1�.�#��<�)�v�E#G*&k��]`_�n��%�B�� +�ӿ�h'���_�n���8r6�T�~%�\wX���ֲ]B2f����RR[^��fWUtŉ6):8���1��Ng�m�T��9�Sr�́õ�0�(�bcghE�@��6�W_��P؍qOOW��AY���O&\�ߎ��n�t�%�}��������VO�8{
O\��Qa���F�&v-`��� a��WH`�1o?)�mm4ʡ���D$�Q_�x J�䷕��cv\�g���T�����ܧ������V(���Ay�������
3�D�[]7���l��%��g�C#����Zc���zM�Sp4��	�F�u3Xpt(��swF��=�U����T-�5؂ ��ꩇ��0����p�Dn���a#��9���AG�TyI-�>�,MCNcjT��YGi�Gld���ܟ��hm��*,�/uS_Y_U�����8�֨jdN�<J����Ѥ�x���z�7/{tk�(o����������q?�%�ʈ�x�w���u�U�2�c�q������-z(�Cc?�dW\�n �8��|�A�k�C �2*�mK ��aR�+���h��_�@�O�q#`����	�z��5; ~�V�u�ĺ�Y���.�u{�齓�'p8�'��pu��Lv��i3@��e^c+dȨ��@�z�B]�l��Ӡ��Yc�o�(��*�*�j�,S �Y/�x&4EL|�ͬD�b�
��>�ܿ���� �>�D���=��(Fy��'5O�Ov���T،;��uێ��s�����R����rɦ���A�{\��3�l�����q!(*(�n;���)`z��q��fw4 �a��Ĳ3ЦH�>�������Y�t4"�Z�Cn|�-	b��@unm�[P� ��K��l�� |ћݟM@���m��,��������Ul�����7���N�����"�W�"�<&�`�^p�܊�N�}OTE���퇒���1R$y.A�g����
�洓��i5��
Z�54�՚���|rz{A��TS��!�,�Qz\*��������!����y��qz6h��<jO_a-#��:�;���٢^�L�c�'8<��m��<G��_D������yb��<�X�O�3	�=�b��][m��j2G�?`�h8�Q2P�i�`(�C���m���r��� ���H���Z�>yx{�$�aZXjXf��>!�c:'���ʬ�0+c�P�w�\��)�$��+V�����U�J<�q�̆�kɟ�����z� r-̓�(nb�J(GH�qE3