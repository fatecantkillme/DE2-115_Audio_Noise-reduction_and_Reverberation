��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|�L��58b�Y��u�m����RVu���?��6X^@��&(N.t���G�]
&Δ+w�Q%H�]�j�7a  y�2���c	�a�}�"�^��k�YY�P��C�}��Rp�Í�Y(��DR�k�4�ן�ΰ�;�X=�-rj�<�.��ϱ�_v�~�B��v�4��N��a:�����{���RfK�X��������r(H�}�݈Rmu��Y��^R��2�謙�{� �Fc���_�1��;'���\�8�*q��խ=<]-��A)�t�S�,%H�l���ܳ�Wz�$Eϊ�S�,Gq}�W�����=#��
�U�ٱ6C7s��l�k�Ę��I[�v|MUG�	l�.
=Yv����ߤd����[�辸:���:\�
f�̘ܽ0F)vb��Z�W�6^�_]������%o;0��=3����+&�%S^�JxC�˳U}Q�4�Ap����#k/�uEم�wmKb�|��'�ul]�%<^����H)���1b�����$<������� ������I�!�c�3�:k�
C��%�Z�'_	+���c��OL<��P�K�����]�(��V.��%�,%�&��|R^�m���Z�QQ�Z�DI���+{ ��/h�V�'���2� �W!�+���t�g�үՀ� �~�d�'���\�/�閹��q�>6��ѐ����q%J��|8��
����=}����>��x���E	`g8q!;����j2-�7N��>�$�#�%�t���t���x��/N�"��<Q	 m�-m����(�}��4�zD�J[�?� �I+��D{e�G����fD��G�&L����Ҿ9�݉<�Wp�]H��K�m1`�ʪ���O;��5��>��z�� Ᶎ��D}���U zb>S�sy8T��
���y&�̚��o*�P���T��>\�f��/mr��)
Q�̷E�^'�Q�S�	��,y�I������@���Ao�i�w2�\	(�cWI��M:k�k9�<A�3W`-��(6��ɐ%E�4h�h�>03�|9l��:���d!(��ϲ��b7[����昭iJ�������ӛ�+���O:1��U��.y�?��:A���qM���Ҩ�$jJ���1�{��$@�kʜ��C��.�=�:��t4A�t���]\��5�h�Y���w���'�$J�-����p�>,�:�?N�Q]��xk��?#|�?�˿�~��po��9�mD.=�H{`y�Y��:#�Ǌܳ"��6�B�k����|N�;+<:��x��<�٧u����F�x��%wq5����I1��Cڟ��ikb��!�L�P�Z�e0�(���)��_��nID��G�n�����R��'� �5��[2r%N8��d����Cn����(�t0�R��g��������iaa�Z_g^�4KDЗ�ƙ�Գ{<�}�����+��i� �JI!i��������?��(�;�3bZ���>n>Z��u�K�̿#�GÇy©�F�n>L�W�~��Sq���!�w�%��G���	{͘;��:��t �y�K�ȣ�N~+�{DZe����R]a��r�w�w|��0�yMYq�;��Y���#�G&�/�%_��9\��z��	�G(sP�g��gqgy^{�G!�?�����E�"Sľ�L�gr�Q��݊��h?ЄW8M��lů�w�􌿘�]p�����K��,L;��؉�:����ot#'����qwa��_�;s�
AI=D�@s��.�f}W%�x9�F.@x�j�ǉ�t�ݝk�a�E�2��n�� B�N�߆���T�����/<4-v*�狯7E��j��BW��^ .bht~Ɂ��,�xh!�!&]�o�p�(6�~����J�w6/�}�Mp(�1ϋMp0d{0� �	F 9���b����M��� k҇�ƉK9��9�@�ݰ��rX/U6*����M^Hs�"O�Y��+S�����2ߟ��Oh0�￷��dш�C�gPc
F�S��9ɲl݅��C\	l1O��!+7~�[����)bq?���h�ȴ��U���qO8r��Y��o�C�h5�}���F6�KNtɊSv|�ѼZN�������f� 5��#����������z���h�����:&���x�Ӓ\U�o�ι�� q��������X���F��k��U:�@�x|}6��4�3v�8m�X2�m�g���Q2Gj��5�ײ�uxFD��͸ښp9���3=�r��oni1����|��u��wp��R��
�a�c;�r=8ݬ��E���N�������,ZLR����T��8*�RB� �e���~�WH�J��
hP�x؏rA������4�k�	/�7�	ƼW�۟�:��2��#}p��e=[�E�����������D�g���^����=Q;X������9̠%�f����m|E`���Ag����+d����S�����54ߚ6�0ɧaN�H�l^�r^aW�ض���;ڥsR@%x��?�?� {Blh�e�T����:I��*Ƭh�4���!��s��?v������L���$�#&C�bF�qi���^��VA]Y�x�ᖺ��D��vJ�S{9�3�nY���-�p�RF���s����;_��q��u�ܞ�k�M�ݻ��G
�}Q�p��_�(�`\J�;ߤ �D	_?���ԥz1:�Lk�_J=o2$��~b*D���jL�����'����^�ZΏ�U��3�#,ό��.�U�:bL�e5��zN���<���������Aތ��Ly�`�,5Lc�2J%�B��zVnd����M�����e�8̜��+%"��H�d`�����C�����9Tj9��1��_sc��=Fp19}q��eFY����H(}Tm���G��LH]p��ݐ��hA���j빼r�&8�"�>�-`>�vɪ��
Q>���y�
UȐ~$5��[m��"��0��{�e��[]§����/�wG���Y�-q�e�R�c�0~��Ѷn�`4�)�w̻��T����Q���1H$��P[��E� ���BJ��7'6�W)[aV'��������/���|�>1��	1�Q���䄵]٩��t{4���g|7z��z[*L�Wk0�X�֘P2�r��ߘ<R��tY���P�_�4Ÿ�!�"-l���������x`�?�.���SƠ����k��vQ�O��!1�-�5�C�ir���v��vqZ'���%�"�4��#Usj����;�&��+L���
�(6��ls��D�U�7�C��D�N+��Z~-9fw��[��ö�4���Fu�k�m��Lt�^�������.Mſ?�[��g�}'#u�2hIڼ�h.\�%$tOB�oB�e� }��{^���