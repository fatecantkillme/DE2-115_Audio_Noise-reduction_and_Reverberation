��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<��&��aL�x/s{j��B�1n��IY}��'�������7�S}�(�9�]��N���_:�|�w��]�I��%N;���P��bA�t/SJl���
 �p�T�0��c���[���L�g��v8�<�������_ڃ�쯆*D
$��:�U�)��o@'��qM^�c!��to�հ��H��N�(<�4��ŋՈS�rџ�p�h��zH,�>9���� 7�t�}\�A���2�I=.S�z�	;��d������ygMN�%a �7��-I�Fi��}��~�������@$j�;��q��ߢ����=��WD�-�d|}Ab��^#P�������|�z�[7i�[jb�`�e,��F@��D�5��}�v�]z�N'-����HN��9�,k1� �3�Av����`�.=Z�)�ddӈ�5��G�����cqH�TAB?B�S�6!���ԟ���q'9䚷;)�	ul֢�Z8�;�؍7ÁN�+�����;�Q�V���O�6��葯�|z
qK2��� ����'��u��Sݜ,�҆����_@���XIņ눲�:rFE�&�[ե��nr������%�S�G���S�.��M��t4R��,ɘe��3���D���|,�ͮ0� �P�S�EM��N�(�g�k�[���A�M��
�6#
����Ż'�v6�g�x:�0�ڷ���N!e�������O	���r��G*��Xſ�/\�!LF9w��|�w!���u�D[�QЖt]����]J�A-�&��9F١G7_��ۊ�Y}��r�1�g��l8�găBɒ��7�bl��y����Z��`	�n�aX�\�P��E+���]��5#~���.�N(��?LDǹ;r�i�Z���ט 
���!���V�l�u��\������o��\<�y0��ѐ�Ԕ��Ӿn�����p)O�����2X���}$I�v������9��%�b�T��D��2�;W��m�í��e�`��}.D�|G/܋��oiN��sD 4�1 {mn���K���z��GY�~JE}5�����ԡ/W��k��'s���н�"�å����^���P)/�F�{� ��\B|�r�&O�G����M|��������������7�҃�\QF�j���V[�[*̤�;�����k��d���}��O��E��H�IC:��ڨ�`H��Y#��7!�hL��7Ӥ\�}�M��|����~5:���B*	Q�P�#s�o�
��� LV�ts�>��()�V��<�|���l,;W��߬�-f�����A.�8��P�퓒���BL\�xK`Q�s]����C�Љ���[�<��_�$<k�9�`Q,+;xl��B/�G���}��j.�%`��w������k�W8����*�P٭��N��!Į^�ގ[$w�Q�t�E��F��>�Y�oc�Y�q}[&y�\=��4�b0��g.!k5��2xoP�8L���PQ�l��R�+	�qkқIV~��}�r�?a�^��F@ӲPl���q��2��TamC��%jR��kG�%���K���7T�.��_{i���Ɛ)�)N�K���맚�1|7x��c��� ?�^	����:V���>)1�~�rwe��f���>�S�:%i*�; |Ī�y����=`���Vc5�ҋ>Zo��{��U��M�+��%��p�*+JC��מ�������yE͊��F�W�����
/m+}h�~D�(��l���b6�n+a�>~�)6�YezC�κA�9��!f��#:�3:` vȰ=�CB*���dJ�oP
�d1-��;�(�&����mjՍ?��&۲�Ts�W~��r]D7�;���S�C�S�>2'���j���1�(�"�|��n#�,ޮ�B�& � ��`.��ri�-IV̨F%�I��(�� t�D�D����� �&�FL�2�y�zn�p�� �l�f<��p�l��g�wV��p�	Ӝ���1g=�wR��� 6��5I��0̩�,��h�t���� ~���Ь�}%0�`8�	*����r߸~�a�L�����g�1�al�Ӈ�9���gBW}�[��/�����:]]"yw9_N<���4Y/ 1a��s����g@ter�&swיt��cNY��F��D�g�c��X��Cy
+�up������r���c��rF�T|��Da�VzݝaFE���@P����y�:;�*��M�$�"M��Z1�`���.�+��Di��j�L��_f�5���k��g����ƅ5q�H���b���k1�������/V�Nڤ�69�h����Ʃu3rQ�ۊ˗��z:5F���J5��_7�e�:�3��;#�7�uԮ-��J�C��r��B�t��b���UZ4�J���}�O��o`�[r����=�}�2�3_e}�c/<�\E�D
8�>ƹ&B�����)���o���������������*n��n�_t.Oz�3c���4����6�A1���P�F�yD��6Ly&U�8��l"�UH�a^b��Ƅ��O��!���Ŕ��;�J�v���&��t��kZL���E������<�s�-��o0�zT��T+�_�K?3�N�M��x�!���9Uժ�gx哒���!�0�n��MaJA+�)\���K�~m!�^e�Q1�1oz;��@4�B��:��X��� l`D�4[��d3�Ұ�lr:S2�LY�a*�R�8�˃�я���&u>���:��U��|<zj��x��G�o2�NC�|B������S��餵�`dRf7�4THiu�����N �$��.8��4N��/e���*}�X�!�̙�%$;���E2������AVo�ou���Z~�����%<!?^o��: ;�1��4�*�a7a��W�{d\���"HL��[��RT>����`�6��S��z�(�{�vm�˘:P�Rg`�ߚ�����7��� *�J�?�No�|�6U_�>���)����~a��Z��i;�;��"mQz_)$�X3��7�m�"��.C�$J�o��m ���s5e�I��(����P���"{�,۹���N��xB�A0@���W_����U-i��v�c+��Ձ~p5s�������@a����� �/���O��ɖ;SV�� c��MZf���Kv��Q�<e-�D�
���#�esU;ڙ^��%�'[���*���-�L��dA���u�ϮJ�r��W�S��#���h�w�oJ����F������I��n��
Mgy~adT�[2dz�C��فR*��5����Cv���<�S�ҵ��]�ȪWy��=�@��{TJVS�j5r��~�+��N~?��X#�L��(�O�g��弐HH��&R��3�q5�"��'3-��R��UrmϪ�<Q��_���,�-zy��bDx�u��������8"I}9�y)��3-�κ	�_�r|g�|A1�a�sS���^�ƎPL�|�K��c�I��Q� �4ѯ{?���8"����/���9��7Cx�	?$]p��q�4nqq�}Nێ<%�=��/��A�mU�2}��j��D?e��\���M*k����3v�m��0t{V��3Z�K;X����Q~6XM6'�
6��6��� ���|Η2m�hXU[�kǋ�WZ��r�8��s�`�f���#B}~ܺ"@��N��`���C��Ǌ�W �\ Ѹ�d)��mD9Hz�4�[�$����xύ�[����,�1P�>0E6L�3}�?��BG��=�m2��M4r��Q>�=P��N�[5�W����� -i�'�M�V�Bc���Tm��d_�T�2��uj�`�	H4�Gܝ�v��妽=3_Qs�����������*i�}�w�ʥ��ٹ����u�K���kmf\D�5ʏ�1]�+F�|�x���E��<M^�@��	Bb���n��R�}���"�Zwn�q���X��L��_���n9E�d�Rtޓ�ņ$뢋��e���ŷ�Ӓ'n��ۃ����w{8.
C'�F����n�@�v�{/K��xPÎ	�'��QՔ�/5E��]@�����2�JS��j����0��Rݹ��[�D60�o^��2k��|n�R�ǭ���MD���&�q)6����°���=���Ն�\�@>X����P=PS���Ǝ�uС؞�HZ����a�_���|�+"��_1t���2M���i��;�R�ѸfM�{N")�y��,�{��p0��m�>ܹ#_�����Q��8<�N�v*��ю]����TcfUħ!bPrA,ֈ�I�M^E�|�Ӛ:1)�R���������w�vy��,V��R�Qڋ���^FA�4d� m0�+)�|Ez��1Iу����	*�[���A��3��2q�\]�g��W��R\��H��۔�s�)����H���l�����]r��k�ɬ�)f ���ݍ�\nk@�ۊ��rs3�>�3!��C�i�\��JG��b�~��ql�1ϳ�����T�\�]v�N�p����&@9��C��myhb3��_;�^�; KZ��p��Zl̑+�BPrH*p�B;�K�5eJ�{2mP>�}�J���%��OEox��d�"�;�uݐ�Q���"�eYձi��Cz��~�($�(�}�o �(AYp�RU�
K��Ot?�!�[�Mݻ|�:�S�̳w���j2��5Q%cXӐ�X%
R'�R��-�+&=�[-Z(ǰ��c̇ᱬ����ҐZpsI��Q6��I��T������$����=��1tE��o�gz
�w^r~Ӛ���^u��[����g�7,��?	���.�u��W�-��U��u���!%'z��h��~�K�V�hƲ�{/�r5>�l����ߏ�Q�㚸���
֟wAs�C4,T�_y[c�h�!:�p=�Z�
IK0j��Fغ������f~�*e^i)[h�0��O"�dX
�'��j���|�[V��p���kZ��V7V��Ir�#�ٮ7�����#?�G�/���(T1�}\�gR駣��ܘ�J��P��jc�n3��p�X�k�I�.�J��+��8]���oN=�k�><|N]�W�+wr�l1�?�r�]h����u��D�9�P��g���w�[��$�$+��
�o�t�\-����6���:>�x�Š����J`�9�EvdVƙV�r�|�9��r_9��[��h�*��kh�n����U�����;��}�Ɉ�����g!�Hkx� �����no
K���<W��m�w�O|��A}��H2���xd�`fΓ�e,���:Q�=�ƫ�ӳ�B�o7�3�m#gA�H��ɐ�+������&�X���(�5U��^���㇤C^�%`��҈β�[�w�H$��^��[��]�v�.17$�н��Z�.{� ������u���ҦS��#�Q��7��yh��F] ����0��.c�5��ܺ7�>OR�������wJ�)Si�g�h�I�#B63Z%j8�LϬ�έާ^��I�,ëN���G5�Ԇotq	��P���R!�@�%3��G�L��1zЇ��#$��Q޳�#|��C>z�'��=�nf�F,��qz�91 .��w�m\���(sf��:�d�E�~�|��u��^61u��'næ����^%�t����d�}b����<c���C*�n��T1Yvp@.
�~��f�uI��Δ4#9�c�1��?���#�9\X^-r�OZz7S"	C7C��}2���A�-�_�.o�4?����C� G�T���R���KVo�R�Rp��+�EX�7c��X��P�K����64��T�K�v����Wi�eM@�P��F�v;�a�X���2�	j�衤Rq|� ���޸{t�]���7�{���F78Οk�T� �J�-��jj�z,T�F� ;��AA<�\c�s�����/RX܇i���P�]ǂ��(��4&�
m�u�\���s�і�̙���b�����F�B_Y���M����*q��6z������,��pl���왡C�ߦ��Z/7qjk8��w��P�:KSw[��t��.ƚ�Ep�1���YJ��FɅ�����m�z�b����N��8D�@�M~z�:>j#����EA�"i��4�;�:�r�F>��ό�ߣ�r�F�_`c䍜@��}��0�A���8O�Cu����^��m�6m,#�#�B�ubQ�}b��cS��������.�:_�[�H�q�n�M�^��E"��K����ߞ�
�����q����tC���V2�]b⁺�#HWojE�9
��	.���弐b~����i��y}C����J�����tvx�@P���^C�i(ޕ����p��5a��� �SC3�C�D�ϭ�y�
E5|]�A�n��,�d�&͒����g�|�F%�g厀����]3Iҹ?P�m��'Ԗ`#�m-���5��9�W����Rr��K�	0�8��d���=�z۸jba��c����3���<,Xj���ߴ�!�Kj��NT��-
t�a���:��3Ҏ̨k�#��Dw�H�;�����B�j�?�?F���G�P�`��>L���j{
4���гo��m��u�Q���[e _vA[���ј��Z��4���1:����E���HC�/��8c �s��*��+�pLP�큶�Т�뉬�ۈ�긿�l ��6�2I��^��H�z'�gh+Vy��/�0d�:R�����Hىho���|�PF�G�ʬ�2?W��3U ��g�Uwêcz[?�^9�{�R{�}�S��t
�O[�$Mm����?��ځ�;�C� tDn��-F�$bV?�ŵ�#f�>n� �̉�ǆ����p|f��#������=w���!����|�J��L�F�Ұ�	�^_R!�Xwi�'sq��!�� C�}�g�62���T"�+����0�����1ҟƚ��'9x���ҥm����t�'#�	֒�>��Ϗ�Т�%���yo�;�P@n?av!��x���6���� �����0�m�#x6u�H '������B(�����t���ߙw4^��2��W!��W��h)��¢.}s��͐��E���՛��XQ[����jG��a�7<�/F%��vFZ��<i��^5i�f@�Pâ-��BJMeΫH���P0<�3J��2��Oh���k�P}z���ܨȉ]��#�(o�����7����w[�5��X��Lt'��n�yFDU� ��Լ�4/[b�����}A�3^$S`�&5�^ h�!E5A`)M�i��yd�Q�>�sx�Z�^ۿ�;�PK��+�4o8yz@�F
=���a���&��RC�=�.�����b�z����l6n��Q�&:r�T6�_6�I���3W���>b����Xأk(�T�M�Ao��'F���T��f��Op�P�
]������D	��_�-���p�t��.>?"ED���E����v
_=�հ�/�Gr�@�/�
F�� �eF>B�*�+"{�:|���#z��o�"�v�#/�UP���[W���j��3*��(�|�f�`��WdF�o���8PިQ7�J����N���a�(�nɜ<vح8��8����
��d�v�ű��8�3<��ʻk>Z��_8%vWRG�w��[�̯��}b�`�Oe�(���:7af����	Q8E�R�5��9�c�y9j�]��~�e kݐ
�o-��Q��_���M����X�K���}c�f�T�X�a��%q�ܑ��)�bb�3|����S����*V�S�t��j �Էj����)ldb�[v{d�o���c��D4%R8��� ����\��A�yAc0z�Y�IQO�����O��C|���XxX)��onc����л��3�hs'��MI!����Ԓ�8�CPm�b���q��US�}z���M��$l*c�ۚ�t��Bw�qL�ԡw���E����1l�lX��e1����&Xfe9!lI�5ݥ�p0�V��xZ��z��V� ��Y�X����\Yf����="\5)+|��^����:ڑK8ཧ�A������Q����%W�a�p��}�N܊�h���~��Ek�Q5��VK-���p�E)%�^�k��sfP�)%2� �
+c[b�S�ݡ~��ɉ37�b��A����$M4Y��n�F%?Y�S�.bM;`-����L?Dk�F,g}/	yT)���6�d+��!z�0u�@ Wg�[W�t�mˇk���F�����iC��ª*�p��߿�)������w�.ù�s���5�|Xlf�<��Nw:� =�@����?�<���rt�Ak�s8yE�L�k��᫅#3j�`zz�-9����+!X?W.�B��mE�ADQj�<��W��$��c�$�n4���~M���J�,y�P	���:#2�<��Ή��<�����7~�"t΀k�۶�Tn��r��mxY��U"�O@Q��"o��$��2=#K��$��� ���|�\p�C��qU���#@V=�:�ujҩ)��
�����j���Fk68��ppک�b��;d�>p�&"sp�r&00&��#X�K�Y7�!�k<�:J��z�����	Ūi� �_�`�G���K�5cQT����tP1C��ZJ1W�[�ho��k�N(Dm��a����q��~M[�S�4Ӈe&����Z��y��8���0ơ*���^���5�l�X8_޳�h�!�����L��bΜ���ٳ�㪥Rkvjp���9TX+�v���:B��K��,=���'�����w?�y��8����� h~���z,h��K";d_��`������4�m{?#H�ҖRg49\��U#Ǥ�nVfQ�`�V�	�g�)�p2KU�xQǴ���p�v�V��|�Of��mSD�#��O�a�V�`�M���%�g��I�};c�z�\Q�!W�aQXdm�+��Vr�{͗�%j�;�R���8� �u �UE�ChD�	��̇Ҟ�����Fw�V����}�`���6��*�K��Ι���F/Q�1W=,=�l<��3VFIr��&�c�g���tB�u_�"�:JC|�s��ƧA`���$+��XNT�
5~���:H}�'Ѫ��
&OzJ	�A�����>�`���R0�Y����!�'VL������'7���|��cFa�����j��:6lX��)���U�@ e�(���˒�@ �.�j������w@&�m�T�P���+��7'��FX�(�{B��q�� ���_;�0n8�����^G@כ�2����3T�XR��P�'M�5��1'��a�/A��;�x۷D�Q�������ƥ�����r�u�cP��h,�)~%�=֤���U��H�����?\dD�l��Jn~8�����vǜ&����yZXX�οCL7�U�f�%Up�[K�R�R��в�b5�����鴕��c��6i�9����h��c/`�<�eA�2���	�-9�܅�mҖ��\�*r�yF�x|���G�W+��b�Q�a�c�4��gk�)Z�!��ir;�z�Ħǎ�RZ���ϖ,��H��Ԍ}'�j7i-~7����|qRTT���!�m�J��)9���#F[Y˳��vV��O|՜��gJ���|�\u�}ط�o�Ļ�;TU�5���Q��s���C��s��8�sm	|3���_]�������9E] �)ݧY%-�A|^���ӥ���k��q�xt%�w�@3�Uq�NVm�.��m��9��\ҍ��Ko�@�s��<��2�T��Vp0�)�t�ޥnkW��;�>�5η��|<��e^�= ��c�G�����_K�1��n֮��6�z�|��}����o����V���2�3��J�
'M��5�K�?�|�Qi��1�y����!IhQ +�p9te1�Ջ�R�%��q�M�{23��=`�f$�6�v�EbLj^] �T��cˏ�� wy�p���Q&z�3���F��S�|��A:0�3��+B�wB�d��ӌ������y��b�t��n�Ys9��H\�!��_,'*s��e'Xc6�0A��>xe�!��u��i�M3N�5F�G�mxbh�N�p����f>)�1�K�g���-A#x#��f愬YO$>�W(�e��E~���P#䡈�H�^����G��ě�LA@��������9+�F��z���t�������:�]J�w�!@���9\m���ԙI.<�`]��3m�@�~^�\Z�NT3���Ą�'b��@�AS��3Z?��Ș�e�+��'��Q�d��Z��ђ	iF��=y�%��FKT������ګ=xky�))wQZ~�#MV�ò����g�v�[8������C`�b�;mln ���$���V�"4Q�	�8�SPO�v��.�i���
<T?)OZ�"�O��O&�јL�4G�]6�Us�a�H���,Pޛ����w�����Y�L�Mj��^���F�z'}�c o-.�{ښn�y ��C�2�׻v%HN�(cn�y��="Y�|��6X����?5�U��/ZfPE�=X YX�szV���1*�[(�'��+c�e�%��G��� ��(!Ͻ#�k��-S�߉�gP��3.�ߦE^�ȇ������`$��s��n�����8��4C�e��H�}�?�6[Dλ�����yEZ������l����4v��4���2��%}��L�3&�[=�P�}b�c�JӢO�fR7}Q԰|�T��c�����<o`%Tr��Dѐ'��+��l��jd��:�4�G�)`|=�}���:O�y�H"�L%������iUuڍ�x5U���!��&4�է\���e����2ƥ�|���q��HiY���sk�MԿZ�Sᨷe���gXt+I�0 ���Q;#�Pkb��Ȫ"�l͋�[�勷��Н�k�e��] S����h_T E	j\n��a�.S�U����gf{V�ތO����o�侵������[�;��c8�
��[ ut�,��̒�]��+�cY�e�'�QI荩V��Ђ2:�vw�߶�mr5�7Z�d�(�����q	��䯂a�?�%��g�"��ʵ�g�����#nUw�Ku�����C��ńW"݈�m�.}�F9�.-o�g���G;��	�Wm'0�ƽ�1h��F˼�Lg��6��A�� ]�ZU�K�e(�����ϔC����3zx��.���^���<���Œ��ѣ��R0��~��ƕ;�9�<�/>I˝����|��=]����>ԟ�DST�f�Z[+��Q'� ���'#y�\^t����z�ꨇ�x�{2d�:�JE�ܻz��45nR��\ap:�4N߰~�P�_�������?.!.:�X?s�~�W���k�����tH�m-��ǟsp�۷pNP��4�^:�S�/���7�]3c���\7J���;���=h�<~�cR�	v��Th��p<��a�#8�;�bU l2�-,^)�I��\!rF�����h��i	���Fp(<OR�?�&3$^z���WQ��9�f��1���e_�0i2A9��~�6G�/ξ2Y<R4"TM�ؤs�|*�!�OUR�$K���`L�ͯ�?��z�mjZ��}rr�_���G�,�����f���Fe�����¡��'�W�Kh4��Z�f�&�,�O;���'EsR��;c�#�P9��G�D<39|+,ФM$�{�Z��Y�V	F�ִy�~��xK��.m�l��s�+.I�G02����&���=�a����l�a&ڟ	k��j��� �U�h�kAԌ�S�r��e��8��$4��]!(��\H�|����^1Q��Fģ�g�x��&�l�6�n^���nt�~wj>/2a+=u�qm��iLǯ��Z�R#F_�iEr� ����9D�Y���\i.(��^�]��B�M�<�B��l%�4����|�m�ٳy��(�>��\��8H���#D~��!�_A�����R�@SF�Raclc�S(Q���I��p;�+���s���4dJv��1>pT-$P��Z@�\�.��w�AB�sU�R�ԇ��ҦS;W�fo��ґE�H�>ے1�+�47>�㨸�-����d��7�g��'gf�)���ev^�ȳ	{�� n�㝂kd�_k��AL���"��b��<��d*���tq�&o���=&M�6�O��m�'���#He`6S���ܠ��,�s+���m)Z_�H�֙��ұe�hw�0�Hgud]�:Z����$%��u>uk��S*XQAۈ���c�߹v9�y�����;���F0�j���h��
-���q����``g�Pc��x�t�/RdR���ʃ�j`�*�����g���5/SB-;�F__A/����2~�Z�/L�c)Z�S �Z�$�ZW�j�[���kd���oX�$���Yd�89�SMQ�p$�웅�K�)�����#�@.|j��C:�V��^8�OvY}#R�^��[R��֟'�A��Qr϶f+�Fƙ9��]{x:7��rxT�d�d/���2��' �DZ�����gɎA�Ə5�v<���%b�N�+J��+2Ƶ�R}�@d����S�2n�2
�;f�P�}YZ��^�1,Im���F����V~�N��V���f?��	�;#�
�u�u��s���燺oa��*~����H|�D���U�1�@I�~���)�G�H��%0�,��k�(q�Ƴ���ԙr�����5~�}��S{�n�t�{���м=��� ��e�����<�\���*]��uծ΁��x���[%�x�*�����׋�9Kes��}�5�c���8#\��9�Poz���Js��r���,���t}U�J=��̹i�y+)>����-�X��G2C�r�J�$M�o��,9�.�՟�^��T��t�[��i(.�������Ѥf7���g���$�*���+��O��ץ$���x2�!Oy�!�uP�C�޿̓�d1����a���[:�����#�o�_�z��S��t/̀p�� a�ŗ֢�@�f$4Dl��3�����5�E�3��\��5����7]�'\R�~�߰��H�0�t�C���5��˓p�К�䱜_�|��8w�w���4�N�J�l?�����J��U2^Զ��{�3T&t�`%X-<�(n�m�iV�3�S�j!�Ե�t4&}��*;���D�:����S���.�l*��	7�k�mTV��(�@l�� ���~_�9���Rx� ���`�7)� �krN�V�r��a?�v�aw�I<�Eƍ!��D�Cy��>�UD/����1y�*�~m�,͗_�V�'�#� �u41�A�sP�U	R����\h��optpE���@ȋ��9��|��փ���9�D�1P��1kD���}�y\�~���*���(N�e�T:]��)b��8�<�n�W}W��]B1���R�\L�Ɠ�5��V���ah ��#K���@��[���g���y��`'����8D��^C�χ����ߚ��Xu,˃k4��[�߆@x,#?B�-��4��������V�=<*�������kj���qx�w#�g2�a�ُ���^�f���=�
��l/n�����5�,���8�{�*�����Zm�N�Wj
_I[���?dYt'>"�/|t���bD�^~*��7J���X/��3��'FFɲj�t���um)��kG�=,p��H=]Y�bǃ��[`*T6��5!�I����	���̜��X}!�i�n/h�m�����-�bTF�w�^��Y�}Kn�
qK���VC~�xFZ�V��A����xm2r[h0B|K�Vv#��F��w�����#%��

��V&� ���|����&C"�A3\��Ƣy+̳��FyN"Z��g,b*�0<����Po��sP<�dV �Q`|#)S��x����>ވ�����������O� ?&�����sO���e!`�,qW���+^���u�h�xA?@h.'��v6��j�n��#�|�\l���,�0�J�P��VB�"�?, :����J��;��k��_8�7��|�jE�[U���F����;�;�奼N���v��5��o����c�*~`ѣ�جA�b7�Q�&O�0�G��`ӷӑ��H�
oY�ݨOF�Z�r�rBt��z)����POt�S3{W�P7'��F�����3�,���S	|��Yg�h�t����Z��vm�����cH���v4H��ۏ�c~�u9@�q��W�*q�IktG۬�ֆ~kzIjI�@|�.��Q�!�<*1~˞�x��6�:-�?�#��T�+.��c�2"��ΦE�O�E��M�F��
wU�ˌ:d�m�C)/�?�z������G��ښN�_�����_M�Qe��
��=��k� ��|���Q� ��o[և/�L��gf�s��E�N]2����b-����ͧ�����m����z��n���}X*1�3|�ܿ^�ߎC��
x�Z�}铺q�*�Y�����*��X/B�% ���6��1�uP�R��c5�ATBɦ�T�aQ?L�=f^d�խ��4��]����X��05Ѽ҄NR9~�#A���KDjYŇt��pz}Ǔݛ��&�c2�᎝�t��l?����!�l.S�k���4$t�װo��Ar�Լ���P�Wt�ϩT���E+0ʏz$�	�D[}f�� �LH'!�߲�FX���v��+���yheA@6}��N�Z�}Y��I�Kkȁ��%V�VXm��{+#Sn'v�6E���,R�[.�Wj��U����Rւ������w����<����L���G�kpC�xI�{Ci�a���XHm�=G���]��>��0	�m��|m{!P��a~�