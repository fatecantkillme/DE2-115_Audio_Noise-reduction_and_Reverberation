��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�8k�)9�k���J�f ۘEN�R��>�Ug:�&�1�q��N�Q�Η������[��;}��ܸ���Jb?]
ۘ�>" ����_5�hky�=�ݐ]L��Y�$VxQ���19\�۴�q5��K����ͩ�?��A)���Qt���QL;(��	`P�<0�D[��P��#p�؈LV���_����3�S{�v�Cr������䡄jC[[����	�X�Vk'ܚ����bI9�mi�zE��3���i�w|	� ��I
�;_N�O%}���z	�\��pA�&\��b�F�n��^��K1F����P/�������d����1#�����(1��`��� NҞ[����j����&`���p�gr��ӗe��۰G���O�@���`Y��=a"�,�����[�L��ڼЄh�}:��}+�`�>˧5a�R�@�}��YSx��E�z���"h��!v�������__�Ny��i�n����D�#E(:�}��И��t�%�O��3�^�4�������a<�i��7a��b>�����+KK.�S�م�;�q�Ǉl��u�{zt��p�ZܜQs�y��l��=Ҟ�aH�E���ѥ1�K����k6�{B����G���T�oO���!�&)��b!���i�	���,*�B��/��~�=��\d%*�%�HJ�	>�)��r�k��ؐ3��:X�b#_��c��k'L��p񜿊��e�$4l'O?+S���`���g�_�OER�⻗}w9����4 I�]���"��l�wi-�Y�Q�oEVIKЉ�Biq#T%`|��h�� E��e�C��"I�ciHm+d#Q(=Tc{��.�Ch!�9��m:tm���D'~E荭�~8�}�����k�c��aϨ��I�b]1mi��Q%�woh���Y�v���$<�}/�rYf����ޮ4qD~8�U �^�e}���cB�{M�R��H2E�k�L(^Z�Cc/\z��	�[1�T��d��o��{!]
����C[�>`N'&�\Q0z�.�����3�)�g��H,�Fz�e���C�	���9�2GIH�b"�~�x^�EF_�[���s��8�3V����TaX� ���Γ�̃*�&Ü����e�'Ρ��W����I���)�$�f�p�4A��މ�)4^P�WL&�Sq����V�4ݢ����oF��e����S?�G�WQ�]�K�q�1{1�$|����U��ދ��w�ԈW7IG`j67�l��\���Ֆ��Na��
uPP�ȣ�����[��S�y�@`���_H>$��	O`%�|�v2��D���A/����TpCZ�$M��e�o�\�LE˶�ِ\-�����6�m�k�蕒Ln]2��ɛ�HC֊�e�Ĺ��o�o�1!���������c�@7,�!���2�T�3�����AQ�~_,G=�(���c.ʀ�/��;���w+����w�
�A�D�/5�1&�Y�(�������W���H�_��4M�j�A>-
v˝4�X��q$���@�����&R�W�-*6�x _�}�)�D��O8�{r�ab��r63��Z���ï�	o����� ��9�
�!�?1\y-�s_��\Ŏ��sI�a
�So�
&��|��=Kwl� ���4�S9�$�'�
�Q�F�\���vU)k�,��1{ko�~�k���y��/;�;�'[�
��nrfK�ٜ�7ڿ���F�V�֧�ц�)��W�M+´��l�6�pZ?ܓCxP5��	"���=��}X�����f�|= p�:+�i�hi@�T��Z4�R��4" ����v?�,��C4������Ұ@&k]�>�v]nMǅ2z��,k��R a5�
:W]��~�K��2�8�Oo�!J �3H ��0Z$�=�|��\|���O|�y׋��턓tTD�l�'�Q�~���æ/���K�kqW����ʹ�#ׅS�(;���L��!ꤦl2���ю)r<p�P������)-v��?���U�KCQ铿�~��
�Ρ��eS��mu��s������l���	���%������#{��f�H���C���<���LȺ�=������r�R��}a��)�; 
ءĲ�z9=�cj1�O�,�G���iK����P��%t�(k�H�>�R9H�z���E����fsgh:�0���
�_��V����ޠR~� �����3���2����?��&��� ����|���0:��dp��d��ۺ��ޮ�e�;�d�) �W��J1���H�>����>7
��
�����X"�Wvm����>D:�':�PD=��J{��
$�'I�~q�=Y��6<F�nt����:Rb�E�1��%��S��lm��*��N�D�q��� ԡV���U-In�Y�s�I�-��%�fI䂱�)��� ��I�r��<=���+G��f֌���FNl���'��s�d��FZ����;dsz�}�]����1�5�;.�Š`�)\O4͆ү�r9x���oW��9�&�m����Ұ�c8�&�(�X����D�Es�;=qӭ���l�S[���q��Cz�@R��?�Aᚱ��#ìiXBIlm�W�U���蹧_����VkWB�0�_�	�@�w�x'���,��ˠ.�9_�1";�b��+��z�A��uo����'��'D�w�5�[ԣ-<dp�TEb؛�U8��/�ę�<�\h�>�8�e��A�[�4`�F&J��ty��\�6�oԱ��0"�����=�+��LZh (R��5�p3(*x&���>o�����:�;}�dA�M�BdAn�h���"a�&�#��6�1�Wq�_��'�`Z!F�@L���Oy�T|&��Pnn##��'�tj����h�`X��PML�eI7"k��2��b ��v��+�| ��)+י��8O��5���D�r��P�c�9&���<�}4}s���|��pP
(����j�C(���^�.1w����I����Z?r��a{f��*ǈ��Ba��m���|�=,�s޺�.%f
��tws������ԍ�w�f4�$쇐�� ���њt�)��h� ��A��J1X�)?��%�qb{d_v6�Ñ�m�7���-gC��qW�;~�w��G �4����v�zHړg0�Ǽ�o��
��T�![�bY2ٶ��ǖT65%_���}N%��M�*��K=���$��(�oQ��5.u+���k������й�
�#�vh�;̹x�1��C�X���_ ��8�NRp��-�&����ϯE��ļO[u����@���j� �証�}	���]����P�P>x����q ��U�u�<�<J�V? hd���mE<w�E0 꺙u�X�bY doc~]~�v`��;�-��"A��F_���n��oY�ng�e\���L�I�QRX��s��n�ȧ������@ʅ���#��u�)�e��@x��P�J������D$���D�J�_��^�{�@��V��g@��ka���Z)S�.3Z|���+e.껇4�0x31$ �P^d�"zヰ�L=�>��"��7���d�
4�U����]g����:�p:U'��j9m2��EL`b��Pz�|=���,���+_f���cF�6��S�*ja?��=:X�IE��0䫘�{�9�h6�'�0�[ �e; �9�����w�a����L3�G��2�	�#5w�iy
؂qx�\���8<=L��Jw8Y�֣L�~5�NƜQ��R/D�|�m.��O+�w3 v�9����́��a�C!+Z�ey�+�\�*c|�-z?�w��b�-o��c}�rTU�����"���|V��-Gv+h3/� �Xt��i	kc���������TL�X�TMc!5��fcۤ�-�ǧr��l��
��+Bx~��wi��\�I��^���עy��\5�<G��q�yչ&�H~�1��D����ⷩ݌m�C7�{D��X�!�Ч�8���L��,��e~˞�\��&��L�L'm��bt����nYa��Z����(���R�W��i���OA�vƕ�б<��"j�LX<�	�Q��?�]��G�����㸇/��
������ �?ٽ=/2���Ծ��O���)�n\K} tQ�����_�$b���$��OL�]-�,���9[n&��דp�)�l%�r���njT�����"h�%���rl��?}TQ_��<��@����9T�h�����,Ƥʗ�m�k���R<>�r���-c�Y�9�v��\08� r�,�MȰ�Ǭ�I0hJ4��y>'CA�,1��<�����x�k��1$����Ǝ�z�' �Q�*�G����(]0��=��H�>���JR�tC��[is�����*�=�G�+k��	-���&�x[,�q>���K,������QFb�Q�C7S��W߽��?ߦ5�4�JҮ͛nzH]��,�z!]�k^+H�C�����:��:�u"@���r3����׭Oђ��'���g�8p�;'|S�ߚ���S�}�nY2?�Se`�uY7�9��?��Kݖ*����Z�*k���]%R����&1��5Z=�8����[���'�S��<���E������s&Sʞ��Qg ��d8jVL��a�P͒5�>��pH�����i^�8�����/���/�92Y4�`�$Y��Ֆ�X���=�"��Y���@�B$��\�����-6ÏY��z9�lR�;dL�V�O��I���?-� 8F���q�z��W�QPШ��!Z7tN���R>3�XC��!Z���ϡ~e������G+׮现=NJr�W"(�4���.�x|����YQ��~ &��`[���kW�VE`����U��()�.����C#�O5x{��_Y�Ma���%O�� ^�'�i��(r�l�� =0�P;B(�!jm�ꐃ:�,�h��T�劼�`�ۿ)���1�Tӭ�m�5i����GC�_�0p��4��0��,�ll�d��<=��6~�w:�lf���^  }!9
���:ت@9%fz�t�ҙ�m�g�����=?�i�d����8kM���l��`�"�^���1�F�s
T�Ҍ�O*�{~_�����Dc��4��I0DJ�b���]o������t�Z���~�HJk�ו�La�M�&":6����@�J��k�}�s�]]Ǻ�3�ߢ�I�$v꠮���p����(T� %,�~zл�س6J�`� 7e6N�s�de�'Z5��J��l�e��e������C�o?.������5�4&�B+V;3��8��6���ޯ�Z��Z�h�N�E��G�9r��`�c�����2|,�h0Lb��I��e��<ƪq�0l_�������*�����!3<r$PG�-�v��y|)�H����ő*f���	\�˕�w�Q7[^�����HaE�5�z*7.�ty�^ۥ�a%P�C��ox'����Ca����'j�̝�m�Xl.�U��T�0���Y؉�M��D
3�4=����d�z\�eYxSF�t�~%̺�V��V��q�6r<R|�.&O��?�5oH��t��]]7�� ���4R<��ɱ��ђZ8Wc�/���qR}����b�M4,Fj��<�Ox+���҆" 1�T���k(
Z��~�q^�ib�%�������L��m��MV�I#���kߑ�`��&=��bZ�Iԋ�9��\�O�@b�}�TQ�Re/N��A��lf�`��O5�~�cal��˷a�C���e�>���5���c6%�:��#r&]A�����6ǌ#ŢdX5?q�����~�X����?$�te��4��~�5u����x�2+����o~��q���/�����6A�`W Q���y����C*�T�o�O�R�ؓEDua��3!:�7<ĸ�$�7��&.Gՙ������������S��ΪJ �VE�zU˄qBtgG�S�U���&���F�rC����jt�%��V���S�ͫ}��7��i�V�����g��t� L�D-�5�r���_	�9>޿l�� �\��U��/&�kz����e����`������Ψ˾��'��r!��q&��.���#�@�#�++a�<J��c�q/���j'# �a&
���*�0�@�bs�x��{�Q���/Ĝӥ���a�ryrܮ���w�{�Z�!��[�#��g4ỨcS6F�W�o �Lq���2XNt;��8����&&���F��F+jS����	��+�S��̜�5K�aPS8�!�b�p;rEu�f�1�=3���-"�t��<+�M�rpa���SŨ[?"�d��nyDm��r�����Տ�Ӣ|�^�C�m�/�?�ǻe4��M���ʨ����V����3Ϳ�^�^�2؅���A�̋Q7�d�5\m�䔡���a��M����@�f$1���K®@�v��Z��� ����e+]�c�
�H�@A0v��Y��u�Y���G�]�+-�a�v�i�o�mN��1�K�P��{+�!y��7��_3�_`�^�#{���v�dLl�4MF={C rކ��R��-�-��U��д�x;`��Y�r�Z	@�0�{R\'��6����v;�������6���$j�#��+IXps\�_:�r����r-���`��<��E�������U��w�wY�����/oģyi��,^�5#�Q�F���#w����ci�*����$++�z��W^�U��L���7.W����"Є�D{�e���Ba�fȿ�h�K��9 G��1�H��91S�?�`P���0j�X3tr�����!��x��O�(
�B��ԭ�-o3c�!�W�����׀���S�#&�(�l�Y��`6~6X��TԲ��ޥ��ૡ!�lcCE̫f���'�;�ӌ����r��$������WZ���P�S7�n����]���[�L4?�Sx����g�6)Ip0�K
�cǭlgZ�]�]�Pfr���k���<7��N(��e���޶������(�	_����vʱ{*z�ӺMVe􆁃}5sܿ�\{p�������8���\(�<)�'���jb��S6��c�i%�\�>�G��74`ej'h��ǑZd�hH��
=�M���h{��I�4�^@�X �ρH"�H�[�Y"�$����B=�+l���L]1Q�f����+��z
^�W�QD��G�L���f�I�n�O�i�8�U�M����Sz�Z����y��-�(.w46υL�����4� /m�߀�Bj6�P+EQjpoD�J��D���X�@��B��N1��&_`X����ʖ4[�Ǘ9+���ZG�;w�*��*�G����^�j�Jx$��&)*gI�l{��JѦe"����\R/ �!�&01�߾_S1� sf�Z#N|N�c
�	������h�(��^ג)�	P�U�-�T����d���Y	z%�~���ߪ���$S���!k�!��%K�&M勺�ڝ_��B��2Et���jB�@F������.MiI�r�ꗤc "I(l�A!�p��{ֽ�{���g��>�B����#-G�Q�H�>��^�^����@�xRt4SZ�Y���չ��@���lI���]7�<�֠���RM��Ƌ||4N�u?�Y>��f@j���b�ZG���x�hk&�P<�<�[ԣ[L�����ܐ1Gճ�Yj�����T��	 =k}oE���(�3~�;�R=�����rh��0�F2�1<M��Gt,�^���Y� ��S\��2����븨�qP���Z�KzT�h����,��\��Mʏ��p��@��Q�)��Z��|mZ��������r �HEm�ƽΧml�e`�kD���X�F]e.�C2�2+��g��������b�����YC!�|����yV�4uq����\82�J>�Q���c��2��p�ӑ=��16��Ө⹀g�3u�7��� ���%�Y�3.8[w!�y��҄����׹iJ���T[�t�>K�ظ y�Ah��j��)��S)Q�
���S��i�GJ�GkJf�8"��O���B�_����	E(a隟s��9t��1�D2V�%��20��spx5A�yn��'HH�\��+�
� �7���~SO�B�$��B�f�H��^L� _���U��@�쥩Y���b{�K~�)^r3��!�s�lZS�Q�VEx�^�;2�k�Lx�就^):Ա�T��5b�!hG�i�b����9�"�����f�RhūW}J/KxU�S�,Բ���?&H��b�U}�{$�9��<�%�Y)g��_0�y�=i1��[����� 
�5�X`[.�[�C��ت��&�Q�Ր�^f~Vg�4\d­@4�ᬹ8�N�`�DK�]�v�~��k��z�w�@ڀ�z;��lf��6�E *%�B��L���L� ��=ZCX��n�]�f̜�;W�Lk�ڛQ�|Ą� �?����W�+�0]=
��7�7׌��b!�1���׷;�����HL`(2��ƢweG�qY00g�$������K���HL����;6}��<�D�)$�u.(a���e����Z�W�G��I�5���~�E8^9Ź��n��r��T	Z'v竌����9eEGA+D�Koc��<��.��f�P�� �g-)P��Ч�QȝYpφA݌wBږ������4�R�tDBJ��J������v?}��b����k�?q��wɸ�}:�F�����{��v�z!���Gip�����ΜxU��~����������
Ԡ�0�t�)���	$��p[J�y����j�Nc���Y(?4�Do�bX��ھGVl�K@�8�Jy�(i|��®��8=�놿���$�������9��	a��$�l��e��������L@��~#���ԅư���D[̠����ˢ�,_z1�\�����B���'����(i`�f�pu�v�<�}+`���2g׀??/&8�H��L����r�8LaR�9J)��>& ��B��������嚼�r;��;��f��$l��6���̀��ǻ���i
�/�K�9J��)�Ѐ�$�wi&p��%���r�����qXd���:����fb�B�(nGy�y4R�>�N�<���� �E�T�����Z�G%0~"�C�����
E��)�Ҋ���yJ��ҙ�2R
���l,GݢL�K�4@�dH�/G�e�HL�HLzn]+1�L���Z�&A��=����oE��������	��
�$Az�/rԽ �"R����
�:�2`)��vyv�ljv�a�^Ca�y��-�	��n�������j9�B�m�Q�cl	ڗ��]��G���LI�+ͳ!��$���H��jR��B )�48����?]i ��A�v?YG��'� ��ʓ�OT���I�B���8��j��]���g���S�Lk�	���dΰV�����Œ[�kV�.lOVz��/�Po�>�4Ϲ-0�;�Ը�Bu��O����~Þ���!�}��_�xcA㹴6P(��I��K����r (LW�艽�p�I}�-ں���
LLya�a>�~��J$�E��u��#<�a���Y�&r���7j��0��(�#�h������خªV: �tr�Fe0�l���[���b!R�]�����"��WH�f��?J�|�a�pV����?�f�O,��lf{g7�(���m�ы����-f���]��d�r�+#1���c8>�Ot���Ѭ�Z�)�BzjN�� �7Em�փO7am�>���2�^������ ����[�����t�pN�?�u5&�8�oJ%v���×�ulc����8�c]>��wݮdذ�i�j��C�:M0�����+�i5t�J��&����sc�6O<��j^���rٮ�^�
]֭���(�g5��0w7r��4`��П�K��(��[F,�����I��%�B�_���+���\��i~����땹h&._���~�?_dj�(�c-�B��4��䤥aa����6ݪc��%gUd�� �^�ȍG��x����,�@ m�a�����1�r��&;P�٘n�hoO�p+��@��;%@��T�(��{�J�_�%[���-�M���\����%�5����~�(+t�iVE�Exn�9y����VhC���j����|�p�ҕ%I)Jȑ��l�pd�H�������!�@r���X	M�kD�� G���+�O7�k��)���2�n&���@Ӊ�F�.���*g��FI>���M'vB��&��j��H���b	3|���Z{�\	������z�rrIq��-���'[0>
=�[�A�s��6P=�Ϲ�����ib-&�9�hP��,}'�������/Ճ)R�f�Q���mX��%ʞ���F����鍣��HMP��CNk���yz����r��洯��I�n�7��v@�<�K�7��bz�%��*���P���?�ﹿc��U恌 �N(��t�s�U���JánSN��;b���sp\�8�m"�|�ڰ&��	�⢤��� yT4���TXK���v��k6��
��?�a�	�E��IUuL?mqCK�:����M����-��}����ي�FΆj��р���a�Q�!a%b+*~��)A� �4�ǂ�w���jI��3udG�R�F����6���������ޭ0��w�]���$iQ}b�:�$�h�ot/�����D�Ȥt���H4�V�����G���Uj9����[��s1� ��I>���K ��(
��y����M���W<T�=z�ܥ'��z���!B�x+;���m/���;#��vP�J��v[
��rb��� (����̹H�`ƽʍ;��� �t�I#�מ�p_�RA�!#sѽX�Ϸ��(Vd+��2��+i�e���͛��QP��b��>HCgm:.��yK��s�|�I\d���Й�/@3�1T��Von�n��6\�ѻ��X��_y<��t�eM����J��a��3S����بZ��ҋ��k����n�MR"u5���$_���h���m	?�=;�O�_bH��[���M_F��ͬ�J�w��D���[w�`�Dܓ�Z�|�@E�bn�
����&�o�"�ƕ�����D��9�3(˺?�Q��Q�;Nc�˵����5%}�v���/�T9f]Jg~�z�.+ɯT�G����F����,O��Zm���'���FٓF���f<�=�^���}�*�
���LI��{����˪��S{���� ^�*@��VbJC�y�3]���	��pCc�Ǿ��l�f��������1��
���Wj��;�K�-�4����_��]��- 0D(�x9�4���u+K��(R(?�\G���^�c�3ox�=p���7��)�`�R������9�M�W�ˬ��5�P�2���r'\�t�ş�X{I~��M�z�ɨ�^ʔ�oG"a�l����i��@�fWut~3�/����#��!7��o:�M��l/��egs'�Ϡg����\��Bc�[Øk� ��������#�4]��Ȓ	A�>�!���S4ї��&�:ώ��;�;��,�P/o�#$��^��B���J� �Ą�'e:hv���n�Pfoq���.#�:��>6�Z���,&�%n�]�����1!�MOKu��D讀�~�x���/�)Dkq,��8'��0��lx	���S7�%�Z�r�of�"s�����A�c�x`�.�}ɜ���p}�F�Oo؁y���
`D)Hq�Wz���J����Ik@��0yh0���F�7^��>��-����v�V�˽DF�V��a���ƧP��q.��%�5�`Ē�eČ�F2P�v%�����j]��҉�%��T��/`��Z��cq����K�@���1��G��Lnl|@X#�<q�����!���:���ϭ�zO���T���13���cj�=#��a�W�2=Ԛ)z�ޱM���1����d��Q�y�w�oҥ�n8ɜ�-zѵ���6�t������%�����:�P��x�m��Ob-���Ԍ��t�x�b%��<K�iW�+��k���8^Ӯ�Ҭ���)�Oѯ�j�}b� b�w�<�Ϭ����M�������|����}��n�ꗜD��d�S�.�Fu�a�Ӷ	@f�'�@���k�7H),]"]q{`���C��ɖ�P�]`W�Mj!>E�q���|[a⸢t,�I�0�	Slj�V
}@Q鱫w���eue��_"��+�fpS}4���z�1r#�k\�ZTF|��ds��G��� A��Y�n�yc6��p��"�!����3�N�-�F���YÏ��m�q�T�6U�\�M�"�U,���SJ%�Dx&��T	�W��9�Ozag�zt&��p��uX��j���t����;���L���R��Rh��s8�Z�K��L����ˇ{�̱?� 5�>����#���i\k3C��F��u�zl�����L��v������/߲�������x�b�;�?����'Y
��uOTG�d!�ڸ�U��� u��&�џP�k&�����n����(���KR��>�{�������5w��`����-�p�vvT�*��>��S�ߺ��-�	����K�s#$ȱz"bJ��rNr�m�m�b��XV7�c$�؜��,ݯ�O�a�y���k���q��u,�]�]�L0�ߎp�Ё*y;��v8t:��fEN��
iJ�,���kQpM�V��(sb\���aOS��k�;����3N�m4/�p�'���n����R�tyU%�I���X�v5�U>�Ӡ�*=v�s�",;��B6ЧQ�UB��I�v�U�<3[��H"6@P��&U�*�+�'�	gb��[��0�B��k�(e�����%�_O��kӜ��*^%�z��O���K��;-Id*_�S3��$��	�x�����y&�F�0�_X�8we�W�S�=�4�SM���$b� Xu.�~�@�B�CW+V��k�R��P��Ë��p/Y���	�
��0�fHr�{ц(׽�)��]���mW�AM�s'��� ���xػ3�w����.}�i0������~�e��0FxQV�����q��[�C��3�\��SЖ6L��H��ꛣ9�*k$���7�Q�j�*���Xb��ay��1��_�B�(�"mE�e�����瀍�F���f9ܮ�Zsbg���.n3��:�����∈�y~ow���j]ƪ7�擩_����7�{��Vԃ:����w~�|�q{(*b�u����b:'(bE�:�ƛ�t�8�`Q��on��	 ��-y �H�7��XT�
�o.rWu�δD~�Ԉdp���v����$�|Q�-;�F5�ueq��8��AJ�� ����;�Z[��RUX�
bz�7+XFr)c3 ��v��?��U��tܦ=�@�
�(ٜ�����.]������N�y����=��=�V`)�x���l1�������bʣ��׮)�\��ż���G�����p�="`��(|l4��jO'ya���?�t���d|yM�l��@�����0�IHD��,r��xEMs�Õ `�ܒF�U��	VJ�VL5e��ka.��RL6-E?+y���5A�Bt�P=�����S��8�H��>�'� �ފ|O�8��o�,\@��L�|��@�)8�����K\�*��&����(~����s��Rx��34�*ѲJb��2�"�)\���!@������S�|Q��2Ey��P��B�Fh���2��A�/.w�J�M��*���O��X�++�wY,$1������;�1�c�����pru�c����˷R�}AZY���MK`�i���ȿ̟
�>%�|�jr���}�{9��{]�sw^��ȟ�7�lWH@Fz�%�ƊP��v�+��kC�_��
�Q���)px
 ��U�-�R!�㬟���Q^�j��,��b;Q�7�Opq�lg��ߒ꼾L'�=ek������8�تxr��}�Ӧ\�Kd%н����3�!��^C��u�(m�:��s��陇U/�us*��j����v��#SNw:�u�uOY�4[��p�t����F53W��?	G��� (� #��jE13���O42z�`�]����������Ȑ� �g�RprL
h�	��Pn�Ɔ��ZŶa薄�4bU�����{�@��B��lh�f��Z ���qf>����V|���b\kb<��{_�A����\��\�c�@Q�"ā-�\r�N�8��NL)�%�b{�z\��@����M�-�A����3P����ُ�1�9�m�(�w�8h}���2�����uw�2���ǌh��
� b%z/�;S�kO��֋ �~�܊�6/���%#�ߜ�#o\\AY{VM�mB�Z�*&P3�׭Pz%�ޤlP��B��a��-&�iJ�N�5x��(��i����%�0��pX�e|��t��ĩ �~��Z�M*���Cd˞�`t�p|l��	Iz�(���v#h? ҥ�n7���cJP�.��<��Rn�|��;OI���?���tLE����r ;Ф�h��u��s��eUJ�@�e\@B\2SΪٶot.¯?��u�yy}�Z�J�t]\@<i��/R竛����v���P��_��VS�>��5�b]�粺`�[�<8�y�!
�}�U<1��l��.�pٲx�SE�����K�B��d���3|T���6� L�f��ӎk�9�t	~�;�W4�}*�E�266B�N\a�5f5�}���ʷl��y�/�6��d�~c��#�i�a�-0THbRd����G����p��#V��w_:��7V�"P	!/�����F���.R���<��O�|��L�;��X�����~��t����SD���b*;�|Չ���������΂�	�*OGGVș�F���,KDbH&_?yX���������������6~���ę���m}o˾r�B�����h��{���V����MI<������X����,_6�x���#,�d�����ԁڏ=y��v�m�
�*�\[�HhB�nذ��2Q$�
�n��0���N�[ �9�K�~o�F��+z��/�������ATWk�4��ZU�ln��f(���
��:9jO�'�����*Bn��*���Nn�;�Sǚ0��G�9,��5�l�/�X�W�U�������e������=����O��j{�I���x�&4���T^Ϥ����{"9&�e;�{ �.X�=J��+9�_����[�b��1f곍���L���}ނ�{���l�K�B�R�7WR�,<#<��J{JX�\���)�-�i:��M� ն�WXp�N�?��j�_�L��B���P��F��)��_�M+]?E�2r���H}QU1Z��I`_�n�� %I�w�U��ey�.���<�f���ytU&��wʺ
5H���07%7�^���k�>"�n�o�m'~�g�L�X�Bǜ4�������g�WNZE�V�A�T����E��;�p'�T(�=�^S�>���>�2��9�Tr�����@G��mjrO:�0{B��~�nK������`@P�D>�%h�jV*�� �>6$�>1�b%��0h�ؽB��e�R�A�[Ջ����H,�R'�V���v7����ў������I�B 	y�E�[m�}+�l���U���ͨ �x��Z@����ǔ�����&pF��^��z���� �_���J4A7����s��}ܤg?�B����Z	H?�>l��ê�� �t5�]b{#\�QZ���
� ����]젲_c�ţ�r���*��_���󌱬!v��h(>_l�w�{�c�b+�$�	�f��E�-�5�/hof�u�>��g�z����5�W�x�`�Gѐ�<ZV<�"���i#	����� j�_��(CeI=�:��÷X!�BJ��E%ښD�~Uڿ��
��[gs��ed	����gY��������iJ9u�6�����@ԱE'|j��1Z1��UJ��}+�D�ϭ�XF=Ģ�ٵ�����u��.��WS3�҉���»��f��C�4����꘻>E� ��4�9�Ѵ���Р,!$4?�D"�Zq��2��+�T�g=IX��,�%�O3�W�V���ǊG�~)y�F��_� ����<���Z�^Ɉ��R��Y��s3��:�QT�
�f�9J}�5\�_���^�?���ۮ.��Q�[<�*J��z�ץ�'����9����^�34��G�&�q�~�ҿ�y�$�c�M�(z I}�Jfv�Zy�jH�[?ܴ�ʎ�������\�7��S8���T�;⹅����V)?&�a�����s{1��uywi9�!�����W��Q�T@�r����I3Q�׻�>l5��D�3�m,:b%�]9�̥�R���l5l䣱������/Za	s<���)����u�BYROY`��㵑���Ϭ��e��F,[\�� e��c)B~+�Ⱦ�n${���Z�KB�r���_g�� F�̙T�
�El �����&;���0���e��'��~�^{g��F��^�=1$�Ky�˃r�AБ-����I� W�"��Ș�>>dm����:|颖"�xT=�bY&[�9�*�9�v�f��K�\��Rቈ�_��{V��@���B��宔�j�����|�p5��\0w	�.���F}3��;1$�2GR�Yn�I|�˩!�fͿn��+��$ߋ�!�a@���N���	�D��T��|{5�<�he�֟=)m>�K�	@ح�Z@�T�_�y�<-�k5�Mdhq��{��t���.-�1��ꃤJ��JOjy9n+8�7�:�rej������[�M� K���޽Q�o���r����g��g7���]���0���8�/��T�����.!�4�c� p��HVn�@
���g]q q$��q+ *u���G��NJ�v��b��a�W�!���w�s�|P��R�Q�(�pt0�9�������v��N6��"Z�m��e���@�1���������ӱ�d�K�1���A��#劼��+�ZK?FJ��+]h:
��b����lޑ�8Z�}�IVU���>&L�ٕ쩓0F�  �	ّ�=*+A��k�,(���g,*c�ZDeAV l�;\2��2rG�qcCP�u����a�����0U�R����UW����{פ�Ԃ�/� �(GCz*x����J\n�6D��^ў�������e�0	X�]��97zp��r-��9"�G8l_�;��Ϻl�
<7���Tw!�!� �[�$TH�����o,�#�O�>"/���������K�KF�f~��gsäg}9 �o@i����L��f`�jE�q(�3�ĉ*$� 0��St��4�b��Tt`�*�~�<*��=�+�o��@pٻ�ʝ�!kv���wg��]�Pp���!���!n�l_=r!�@�jw7�n$����ǧ|��}ɴYM�]��.�cny���~�7�F�2%�2���G\�B-ې�w�bZ���L���YOa��������\8��&uo�I
)������!����R����wB��z�M�4�9a)�����NX�z��c�]0����'�9=�2%�vZ7��� ���y�CS��c:Xd���2�b��\\���X��O��jV<��8�Pv�>sV��9"��\)H��S��aeS�m�V�p�TH3��!����v�#V��)|D�*��Z��9Xz����G��O�9���'j��s�͗��&�Ǧ���#�ų��஄R �B��`?wl�N�-ڢ;���_U�b���F�V��u�Gr�1�N?,�d�jM˭Ȋ`9���Gw�9��E�B����ع|Ѓ}�e�������+޾�;{7�3��Dg�{J���_ձ���^�t\PLp�#��=���~H�)�j�,������bo,��66s��ɍ�-��+�����6{E�q���{r/����Q�[{JH�n�s�cy9��W^&G݄�G^�Ӊ'}?/�v���	���F/M�xS(�Z[DT���9�L��i�x#Ӽ���]ݏ<�7����u��$XZs^%�	��i��
ʼй伨��0O�]S9Tq�)t��'$!�c��cA×]��mL@g.چ�	q���|��Q���ߑ"��l��m��e�t��,�� .��)[<����)�xk�]��=Z�=�DC�<M��>��^#��<��h"%&�,�:D b@��爐�٤@�^��9�CU�o�RN�p�kLG(ƞ�`���U.���~Ep��V�*d������-1Fr�":-��s�ޣr�F��ωL���(!�Ir���;�����"`����r��?���$ ��S��������y�N��ig��_@L_� $�bO��pm�F;�k�c��������B�>6�]��:�̈́�>��?P-W�����Ȯ�-)ד4}��^T��n���Y�z6�KT��P��o��S��4��r���s��?@M������Q�ɫ����aoF)��P��O3��u�Q<��wL���>���@��+����\	Cҙ�#�'��gL��t��,kr�;�E�7���D�9R� �%=l�/�0�x!�{��=͕f9��������\� �à�x/q{O��At��捯�ǒMl��?>�@�#���L�&���KĬF[��`fOԽa���r�ӛ�~y�i\�>���!=�=�ʜ��󰢇z澁��1�9p�C}����/z`z��$�ȝy������ʖ�W�;��%9w��������f*3�0i�=Y����.]�џ�
"��o�!���U���x3U"��tD�ǫ�@��Y�mKg)fy���V>�@��4Dtl��3����@0�Z� �\����iV����xl!m��BC�4�R��3K4i�S��V�ͪ�RX��Ħ���_�ݴoJ�^c�6������@J��uO�H~)͸��ԬcTw��e�\'z���.�ܓ�ƻh������A"s�߳������N��^�����#<gu|�@w�,c�)
:�H$�P�ߒ4�Vc����u	 ����t3�!��1�s������w)B�����?�LZg�J�e�"@����
�zG�be�R7�_?w�)�B1Inj��]Zܷ�:�����H�srм�c�CK�"1��C�QM�9G����T�ѫ����F�4�$�Iq#� �n��C�g�������Lh�J~�"й:�F��M"L@V ��5���E�!����eq{�:4 �'�A��!�ߴE����1��.��e��HK�'���"7�%����<,c�xP�&Y�%��-�n}�+Y��{����@��G�4Ker�<�1�f(��+=�b.c�y55Գ��d�8|;%��(���J��e
b�Q4}�@�=g��ov��<��{����T��os��z�{�e��z4�ͧf�ǰ�����JI�n�{�}|л�0�(oXK{
����J�J���qԲ{�����ݓ�� uBj�X�m9h(��ޓ�R0�q<��	u U��-@�t�"ĉ��w�5�<*�(f!k���1M��������%�O���xy2R�U$���m��X��{�5�-j��L�R�s@����Z�-w6I������N��tɻ�39?:J
�q��:�`�#8�S:x��v�.��a��d�����|A�KD�����5��S�HR���I����&FϡN�{o�$|��6��f23�Y���z�vtO
W��(�\s�Æ�]� ��
�.�e�>�$.D	�Ry8n����I�&�e�a���>�0�6l?e[��i@QXX02�##�M�T��i�*�J�IY�j�W�U����.�6�������u����2����4l����� ayZ��<$=˦,Ycf5)�pS>�aZA�f�W�5As~�,̮c �9��9sA��ٽ�R�Z�51��iٻ��@��>�Z/������n'��<�I	�@9��Gzic�p�Ϸg����( ���z��Ԯ��TN m#!X�X��PK�E7�Q�>�3�[X�>W������I�&'���tG-���]m6����Bo�+ᰶ�v�v�FA�=������]~��[��kN�j4uW�$�H���xm�FDOe��%Y�F��J��MG��O��5�X[�����M���t���T+
����i�`�'|�>�5횦v�tf�X���;��ôP�jv�e4l�y-�onr�ܵyW���c3� TC�xM(�����G�s�>�Q���x�i�!a��σ���	w^
J����x�ƙBKx]�(qB�f�@7���)�g���ZJoL��L�o�+�%Y;��jY�rQ��VU�D��BM|l�.^u���(�8�R�
d�8T[.������v��Y~����0�::U礘���YD�n�$$��C�a(��v4��tX([��g_(������','3���c�HCԤ�%Yc�\_Q�F$��θH�4M�x�RM�ӎ�6Sӏ� W>�g�)�8�m{>Y��0���f慝��b!�����[�q6���S����2����^mK�")^Q7���A_A�%����ΐq��:u�#�~;�7�yM�y#��#�����X���"������J�e���O����>�yo7b*g�(<��ş�O��L̐ZF:_^��d�����Ͼ�1�vE�+'��W�1�b�[Rx����ͳ'8�BUʹ�y�'U�cU�X z�_�+�6��_�-�?�3�*M�P��]tF^g.I���%@2F���i�1b��ˆV��؞�e�A_;�69��$ސ���|���+�~�#�@��Lr�|��#fap:v���Le�&�F�+-:&���*j�֚�q�(M�_�� ?vg����!D��m�T>P�.1'���%֑�m�A��T�|Yx��,h�Ŷ蔼u��L���^ `��g��L�j��G]�c���-��rfS�W��7�Z<���k����Z0�j!����|O,e�,�M�GǀR%�o�ٯ�{��E��n�ˆ<�f�W�w!S�Q ���2@�rI;b5��)�1D����S�E%���tIF[��Z�T��bcQ����82�������ąK��a��
jκy�?�`ӡ{���������r����K�[���m����%�jg��@�[}{:�.7��?�L��n�7�n�fG�JRB8��o-'�s��M��&A�$�5�s�"�s~]��ՠȡv�\=�j��b�1�U���Fn���Ga6Kc�E�` �~����Z�l�S!e��cP�?e����	��r�H���!�Y��5�$����6����&L��5����`Ia��L���_R	�9R�7d��W5��g�qC�W��~�%�B����F�o[¨~ _�j�	���sY�͏��4����_�vǟ��"������_��^YBՑDxuTy���M#ݠ(����I��'w�E��M�/L���I�[~d&b��'�]96�!�'���p4��)�p	&n8�7�j�1�S�)ê�O�6�oc�c�XY��F�w+G�����.#�U�۸Zy�уgN~l�L䆁�c �1�J���ča.1���hV���F/�w&�{Ϧ�\���l�$�0��[<]?�{��<���h��#�"�ͨO2e������ln�61����9=f��Y�fH�S���Hъ���o���pI�U�w�$T	?](rK��r��ީE��i*�!T\��񷽧�37 �J��M�����6�k�QO��;c��OȦc��[;Gq	����\����4r{X�wbޑc����*`�=�7��/}ȁ�G�ռ0\[�u��n�v5�v�i�_m���⯸�k���_!]_���פ��=_y�P{ā���.�#�5�?%�i>��*5_I��� �:E½�_/Nؽִ�	���K/�xj!�Kߍ��s��B���a���>#m8T�Խ`�I�_8���1��~..���ξ/y�yw/jE)�hj�	�z%�$���~ڑ��Δ�K���s��E�Z#��M�v?ī���s��Z���ҍ�^!�����c��H�~�'��l�:(�E�wƊ�r���&��'5���>/�
Wb�nK=]�4�:w�Hg8�qx?S-��|Y��g����E�G��i A*7[��8}�ќ١8��{����W�����5�2�y� _�C~L�R��]�(Mk'��um��O��o��yV�=:A��MŕaA���e>�A�'e����'�1��t���|�1C�/�KO��G�Jf:�zq>��D���
cҢ�ҭP �F�����U��VC�������-�x��z!�{�k�j7�0ۂ����������8Y-R$�b���Z������m�$5g4-*N:N�4��	8�*�n�x�~4��2�h��y>7 �hvW3�+��E�m���Q(W�T[�o� MS1u|+��M���M���t�Ng>�]^"�"�"����U^�k6R��V�ӷש�F���0ef�#�p�-�}���� �q�.=*�4���A�-�Ri�
 ����wFV :ZW��9���p)\�e#���ZL�v����xa�l��w�`��8�'�8jvTe^�ͫn���C�)l��)٨��i���e���t�G������9�6��(ys$l��������;�]]�w��+��z��-�V/�ZT�����f�Q��r�T/n ��+P���W#ls�U=FGaF�qY��J.L?��c�M��s�'{�Y4DC����A-�G�[�)�B�d��kk~!F_}K��6��F���~kͤ�u��<��m�Ua�"X�U ~��	�������>����Ǧ3�� �v~y����O$�D���\A�*���p��d���9F�� V��J}gG6���ώ�V)������r�eKoT
�^�S@	"���]��r�J��l��u�ؒ����D��N����Z|�������M#Ui��*܆�b�ߙ�,��´��>�7iO[a�ٿH��֚z�v�?����A��G�*��y�{M�kl�10�J�����
�L���q0�B(�!�TY#�V��c�{s(꼍�����G/H�N�Nk��S�1���Ō&=�=��l�Ұ��  O|$�{�.�`7e���TpC/*2Jd����F�u��Oi��PAN'�E$��,�Uq�����of�\�U�oWI�&Usax�)Ͻ _ۅ�Ƹ�˃K�MMS�
	2%l�m�	C5����d���)Z��u!����!�b﮹P�5�И����ܾ���x�Y�(�����c�!�?�����l�2(7XD��w�'>(���E��q$3�q����[!q��t��1����X�i]?��X"�|�pi:q,������+��QAd���m�]4��]O�JU���܀���]U�������ʭ?'�\ �T�)>��-ni����be�V@�v��p��m7r%��J�9i�ZU���R��)���B�@J@��i��8�����?�T�@*����ZCг���<�`�Be85�m9%*�����{.I���$~O(:�O��)�H���)^�[5�W���kS1m$�e�{���R,ď���VF�FNAE��jN�(�Qb�r:8�����G�� ~�F����쬲̧����ݿpޞ��|h4l{<�ýGF�:S��D��~����ηX����kG/�-�����TI)��>Ύ�Bi��"�6�Ě8�%�#�h�u�ƕ/j�«;`�����E����Yvc�Q�7������jSbao뎅�s�UG5T�f3��P�k&�/��̡�c`E�G���Ț ��e<�IA�e�V�剪 Z�(ĭoٕ��%�^�}n�=�b����z�Հ�(CM�#6����i̍|rݶN�{��o�<�9��?��S_Ut��R��-{b<�ͩR{6�u!+� �CzL�����F/��C�ɠl=�}�s���]0�M������K�dK�z��]d�����E͝!]/�&�J�v�)%.(��"�m��q����ii�&L��y]b��(�f,��4��H�j��0���n�C�;j�:E��#�����vfߊ���5TVD�o�Ӟy��P���q��-R�Q*M5��5��$XR��a�c;�����h!�Y��\)��T�*�ֱKZ?���u�=8���~�~J�zO �X���M��o���w3t�΃���)�>���8Z�� �C�G�h�e�W����i�*)n�,k*W��a�?���Tj��u�j���f��/N�%�`�#q	*�8��iO(秜����W�|��衤��i�-`eV��ă��т�Ŀ����8��g^,Y݂�(�"�1S����)5�#$f7�L	t\Ay��m��f��|�Y��0�I�%r����$\�,�O�E�p}+M�Y�G�4ko�G|��;�>��(s{�4�2`�-����N{��Y+Q�W�h#�K�ݭu�d�J�죺 "h���s0�<kǕ�#��R�TXh�^E�������6F�1��[s�<��)��̓��| ʁ�&��"��D{�{F才�;�M�Z�+&N�]b��]�9��w��3��Ȁ�r.g<���'c���K���	D��TGC��M!N���`�� �L�چ���T9���-���2SuƮ�<9^�e�-������U�ajû���)�Tu(g[�������]��M��G��7"DB�����Mcmm���]ݽ]�4P�F���M�wQ�ߠFl�i�Ż%2pe��ǸX3t��7�x
�T��Ui������J�Eթ�6�\*B��p9Fx �^���}F�1���l���2��@�I��'���K�a���jov�d����� �����.���s��C��V��.��c�ؔ���B��T'-X�ߎ�p�x�3�4	�<zq@��1_M�F��[H>@
�ǵ�8BȎD��n�X5n��?u�"���0(�p�_^�&�mq��*���K�\"{�~��-tH�����뜃�׉����9�ϕ�J�Q���N����\qد-*��il��Ʒ��S�����@'k-�+��:%� � �'�Ž��K�?����K�k�u$�"�}F���Yk:Ej�$hz�!��.'i���9�D��xF������R0�E|�y�K$u�2����8Z���K&yA��>��i�ә�JZ*8�Ye��{��V�X�H�� �B\�\E�����!3Pu�l�h䷀��x��%�m����/�im�F�����{�s7B�H�m�5%%*>\c�hzx�]��Z�~�	4�P��������S�.\1�
��7'��F�E@x_��s����9���NRq&�N!�r�om�F��	��uk��	#T�
�m���w,�l��b�TdRk1��N֜]��=��'*�%�;��u����l[��O�%�<1ɗ�<D;J��sy���@�ET�Ь�&*^B M++����@���mQ�j�"7�9�xp	� ޵�Z�k���!%����^m����ƶ���t΅��?#tT�׿٭nL�����G�-t4�-r(������W���䞜[T����QHI�Z�E����d�w���L�O�D����/�Y����=]�Y�d*R�q� \�fv&N˓����r{�����rt�Z[��_����8oU����K�������x�))}��C�DVXX|��\�Q��ւ]�ż퟾�}O<S�t�H�Ck2ŕv6��y�h�B�����TV�t�!Q�������έ:�������ZH:]F�Nj/�Z�f� ���\���K���]EKCb�`[������L%�44$D,�DbUa���y�h������c���*۶���r,=	/2�e>=룟�M:5T�I���o_�A�5��}��5p� ���s�:��4��Lyr�k�Njh?;WU|���>�E�u]x�c��Uu�X��ւ�N��^Q��[,:g��>��K��������I.[M�T��Y}]�#��Cю����q�NΩ������T^QKZ�I�7xz���Kݏ��
���=��b���������9�I��>&�~̙dֺl����n�Vٗ_��������Z���7�_Bܧ��+�����)a��]#KH>�&���]-"7c#�����w��X�
�:��	bֽf�HL]cb���^��c7$; 4��<%�u�r��+���ݢ7��0;�+��Z�p������|�,T����)wA��Q����]F(䍱����5����ءzr(����=���K�Y,"��E͜z
�T�ǭBPa�����Z����eY\�_�?����PE��v���Lɫ��аTC�⳶ԁ���)섰�ZĞ���K��.,?�D�0����`T �ǎx6$-z{�:�Qa�''�J�`7PCa��W%�e��T��}	غ��[�4���4ym˯*.�s p��H��TE��ARM�j���ʸMgUrڥ��s|%Ǉ� sT>��a]
����\d1؆Hm��r�����M |ip�Hvch�B�k����ܻ���紭�C�_y����:����������+���ɧ��J�x�����: ��׼���2A�'a�?=�	��|�N�΍��aD�����{�Vyu��Pu�À����Ka�2�Ǒc�j�k�1]AP[U�A{Ԙ��#���#��1-t T`z�!��}���<�o�p&K����%F�c����C��S��#��'Հ7w�d�K3�lxCR��B�*��ݥ��%*�{�ש=�'�'1xf���3�Ak*A"#��ue���%�c=K<#1�loO��ąq;�KG<|��K�h�/�"��9����uB��G��Ly�s��K�5�A�p��00�@�=Q�}M@`r^SCM�i�<���4aZ��ȵ#5#�m[ޤ�ˍA}+C��{C�=��FPp��E�H�(]�%��>|mDkʝ��3��tk��XhP�B���|)����e�<��&����h����-��]������E^=I0t�aaP�����$�X����G�|��8���!�V�oT��J�K��ߌwff[���WS�b˾���l�Ko�3�7��°Z�]��@׫�]gm�DG?�K������o73��$��:��=�#l���齈I���S�,����n�7!�J}s||���j��#�)v�[�EV�om�c @��d#��~�/�SiM�������/�Y\ҩ8:` -!]xYQ�'���J�ĕ��f;�Nγ��]��2{�f�"9U-�����BȜD%�����C��~@��O;����"��6 ED))�ᯏ����@{�˃<B5v���'�IcF�+��H��U$�k�(�N�L��T��{)�D��76Ī~��?�M�A<O�"'a6{l<�b��r(���%��	��ΧKF�y	~	~�h-������V��;w�:�R�/(��.�T/̭|��`\b�l^Ћ6��*�GK3�p�^ɪa�UtS&
��ȸ�͛���+v�|CJZ�*�:+�n�i��z�m�Dp���]����bt�L� U������"����u�/Tx�U�;����$�d5��D�Y!�^Qx\����Y.7��s�n*��_!sbhjwɤ�ʄZ3�� �_U�b�\v�(C�יx*cH���U������Q.i!Ǩ�k��;�j(X�BuȍY+M�80sG�ӳ��I��y��'�;L�K�q�d�M�q�Kd~h0��?��`}'W0����8)P��e��� ��a�_�,*��ZIqLB�G�jK�{dG.��ʱ:�8�84�u���ֹ��Q��%;\�%��t69���C$��g:�5�$5ū,j�Q���>�^������0�	�><�}��@#kaM"H�vG2��k�����쒠�K�y,��t��cg�:�KW�4�.bJY�p��P<�S�b�BL>���O�`[`L�2-�.FT���M�s"s�Gb�XNwDs�+6yP]������+���|�G@���G�5��C@@3Cdoe�<��`�� E��.L ��3� `P�&��> ���fŪ�O�A���=�Ʈ` u���l_��v�λN���u��:� �@g�&b�tj+�YWj���R5ݼ^���3|[z$rM�/2���f�0fs�N��P6jV���Z���v�n�����Q�,39D��?ђ�����q"�.�^;�0Z
��//6Yk|�E ��p��l���FN���E�N�\�����L�:]eՋ�9Z�����3���lβ	N�Y�z*��`�G��c4
���R7��`��"����}n>�����4������<K�.��� �KF�]�K��g�7:HKUKCn��0w�ƚ��x&'�=��б4}��#�\J�M�6NƦ��"�Z��fL�^�J	Z{w�Xo&�� �E9��&k��er�*��dF��~+�9�����]�g���{}�2t�V65���z�����?[��1[H�*���T県�����k�3׸��IO���%������J�����t��Z�h�έ��c����z܁bU��#�������T�����EU5K����D����5(eE˭�^���g"�s�o�=�}q���DaF����e�+�8f�û��9'���k��.{��q������1x�̇`���`"FPg�f��;_96��	n�?��f�J7�N�hlj�{����v��LѪ�%)����
���3��XEL,a� ������\Nx�	ɑ]�(���P���I0�j��/�U�ɏ�{XnL�����r>�c���*ƨ�<d��= r3�p;��1-L���2K�Ǵ�A�I&}P9�ںUbcw��{Րp5,�T"vJ�Zh�`j3�{ 3bsE������T@B���0d�Dv��'���_�����yj�
[:7�)
�4|c`�<��X��S����EH�p/���Z-�[p�c(]ոe,��C�e��	}�Q��@�wI�Ŷ�5����
�c^Rb>Hn"�S�D�[�O�����@��	2�hk����%l t�@yn:�uT r[����Xɒ��� @���<��Z��c�n�8�-[px�7�3�7�ve
d���TN~/��T�V�zf(���������&�y@�GOu?xA�5�����_�p�'Y��58��;����u��IWZ�˵'��|M$��� ���yb*���7���LA{B��7Hk$����#Y�����y"rFo�#)���-�0��Lkv����6������G��R�.����(EA�}�*Z���QP}J�/3pE"P�?�����䝾vV�,p|�!Pڪ|�̱�٫4��rm+��m�p�.j�.O7Ư%��naR��ľQ�8�,Y��U��Kscٶ�#5�L�c���
z����\��~ﳷ�P���BFf��I�-tB�����������;�
�WNp�.QXT� ,�'_�-F�Gb"����ٿg�t�$��J������d�m�{������Z�#�]C�wFV�U|��/�{t���2�3���N~?�:j��"6�0{4�5��O	V:YR������)�ϭ�"��elrT �8c��Cڰ�)X���:�����e:�Y˒5c1���NY����0�:�.&�l�`�����mW����.h�]`�t0��/���ʐ����N^�W0�iK۳s_r�ޭ��0ߘ��P��3��G�4�f�h�߆�_��.��:V��N��<O����� ��^g?�~�s��nS��n����pWĮ<!s.2ϐ��K`�۽5O�`��r���:�����Y�i0q}y��J�]hW[f����u�a����d,��R�r���^5qF!�C�Z��ٮ���>њ�.Cp& �| ��~rO���2V��_�oI��G{�v/kB ���R�Q`�܀�59-!�w�|"ڢB/����6�����~�Vg�����-���<�ɰ���eU��a�N����1�����