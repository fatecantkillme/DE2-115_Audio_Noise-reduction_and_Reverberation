��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<��魁�7�f�I��-8�����ȩ�[�����>R���X]� �N0gޑ�.�-X%��=S��k���R�s�f,�uYn�b�Q'";X>sk����H'��hSE�z�I�r�����Fc��Bx}�O��~�>w�5���q�Q�	�����x�ݮ�*c*[�U�&{���jS�{}�DZ�9f����n�FH~��~Qr��~�b�^��ǆlվ�zT#�va� �u�Q�֛{�vp�\�V��������u��l�9i��9֚��(�A�Ե���H4��i��6�W��/�9����yEW^}���Wn�|��wW��~O��/���L������.��3��d���u�#�=��%�d�-n;\�P�
��u��\�@�5���w�Pw�#����j>
W!�%$�GSP�q���"�Y�{���u�ߺ�I���_���H�]�8~����8�C^�Jdt�fa��p�o�hf�Tlq8�$�����C/��w�����$y�WD����G�g�K*�u��rŇ�Q�3��6����Ɛ1�S��m���^|ǜK���(q��b/�}�wי�u��n�������YbDRx5a��m�jBpm�D�י��j�:*�~�\)Д5zj�NE������>+-ǅ�?6j�*l.I|@��{Q��ɍ�=	��>&r��lo� �p�>41*�
��=̾F�Dղ��Jh���4�|�^�ba��*�?CtKG����_%�%"*�&�p}��[4v~���/�l1����?��lP�p���Ģw�-{�mȑ�ú��-=�"��Ґ�C��Ҙy�׎��Ɍ��С�!O�N�CE��1��؅���(�[�ڙ��$�R��J*U�AsУ����:�s������R�2�TdD�S�Z�	�c`��'X	�[�kc@<���]p�"��=�r
T�L�͕Z@"����	P�)h|˲{�
�V�yQ�D��QB4��ݤ���/C0�FLךGp�:�-�c7�:ʚL�	��m/�`�F�s-6)�zk��B� ��l�X|�7���-��Z�\eB�Ta.y��F��{�_��͇��3%Gɣ��ґ��"�&�O<��dS����c���CP�g�8�EV?k�x�qh�խEe���̩�_ց:%�2 �4/0���KL����c��7:�n~��b+E����?�*j/g��Ui ��#���DF����ƀ\�U�Q[�l�q�:����Y7��ޥ�P!�6ף���g*t�'�0+�?Z� �@?�ax��pգ�/����LL�����{r�z�#�8~��(
Q��6ۉ��,�{K�
�^!����^�=X� :�Yęjơ��*"\���J�����	"�ּ_6k�p�A=M1�ǭZX�P�׋�pH���-�3�
�g@F���뱢����X��1������`�cQ�K0��Ū�k�*2��/�Y�g��(Na}��+J2�BˆL�0����ħa�s�"��G퍷s�*���Q��jՅLu�d>{�y��ԦK!�.�+C�@�4T��#~�dhl���`cb��ϦB�!�g����	�ki3sf���W%��	��I�yɢȏ;\p6�lۨb���1L��+����Arvbv�Ş�A�pz��+�f�z��7wr�,*��Cg�8�J�OBK�/x�޲���5������E� �֢�=��σ���
9��.2ƭ�f�b�c����M��Ы�2�l�w!�I�&z2�+�8xH�o��$#R�8T�5�ƅ(8��K\��q������h��|�lJ�tK��t�%�E_y���ȇ��a�0��+ ���ڪ�SfJCT���"��dׂ��[���>R���������n<����P�n�4���Wi	����o�]Ad�.�����T%Q9/Ӊf�÷v���*�E��'�|��>O