��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�8k�)9�k���J�f ۘEN�R��>�Ug:�&�1$�[Zw��>�E�C�f�fԓ���c��my9������;�o����'��{�ȷ氎82�9��7f�� �B#Y��?l�m��*�O�~�&�,�+T��+qq/�lTj�0���	�}�krh;�hʮ�ʙ��*�۩e��ě�
|$3{b:�Ss�#�AU�`�o�[�<�2o 6���7�0d�Q�B��_��qܣ�j{�;��Q��m�
k���U N�$��<i�vF�-����'��Ss$��Q}�1�p�9�i&�4�[V~��)l���s�^�ݵ�Z�ir4W�w7W5	�6�`C�1��k}�S���
��L�;���	^�7�'�!���#��މg���aW+�ľ�f�`���I�Ջ����$V8B���!�fCV�����,E['舱Z��vCF��QG��a�#@�?x7*�Kzc!�ܳ������M�ˤ/\J0�>+݌�jrS��V�Ql�� �4�W�3�f�ʎJ߉�����h����5��JX΄\Q��,�-`+�;�q4��X`2�s��$�s��R@��>&�t���+!<S�W�����#�w��j㫞�=��wS&
��~�'�9]sS�WF��ˀ���� d��a@���\d������o��՟��J[�ɴ�S�v�~
n��;�ZV��ǿf��F>\����]����Ԋ��5�����ߴ�$��ٛ0�`�Cxv�=�a��vk`O/#ڦ����d���x��y�[��Bzl|�sM�R�,n��;.��F�N&ɉ�;��i
��H���3�N��G샠+��,�l~�r�+��x�����2K��>�G��4���5L �ޞ�D$�t�TyDiWC�8�"UA=�
��?������Q?��gBZgw�8���8#���>{#������c�"	���K�엂K�����%@@ĭ&>�v�S1kL�P�D[B8v�%9�f���W�&�0ߐD
�&*����?e��`C���-o�hCUD�u.�=~2/�	/�t,	j��-!?g��!שϓ�3_�O�p��pT�5I��th:�K�b̚��bz���pb! �|D�T�+N�v�������]c3���-�#��aУ}hd4ú7|�����S�:��zJb�O�(��$lU�>ۈ��ԁ�!��*���C%�&a�����T;���ܰ������if��mgp<U��
L9��q����be���ќ���Q�?�sC:'���_H�/��(��K]^��b�x�'5���~H���|���@�Y�A�aq�����i�������vH?����5F����jP�)��R�3����$%��tԻ�t�m%�5�ktR�d���0`Ej �O�Ӧ4S�	��M��D&#��bZVͼ�˶x"�4,2�䨖ۿm�|۫� ����6��O�e�ߌ���)LQ`��q���ۡ�%'"m�G��a 0)�J�����
�����)��װy�� ��i�T-W*�.�`�w��ֻ�en�2��W�$	NL�x�� a1C/�-NHy�U��E\O�����C�	 �t��!�(Co�'�!�ѽ�^G �D��&�E
��~4�Pb�-'�>s'.�{JRG>��%Q��Aȳ�=�-�3E%�o�v�����b���cm>m�T隬Cǳs{p�V���7��d�A׵5l��xlU?!�43�	X n��.���z�s<B��S��v�:�-$|�?P����^Ƣ4ҭ�[���"��-=��x����1sĐ��P�p��{�
:%s�~%p=j�\�+��;%�/���P"\��������e����y�M<'��>XV��5j��,S�N5��6��ϛ1���]�F0�1]3>]*��?�<�if��b~J�`���i)��gYb@<ź�ȡ^k9�㾲�SD����RB���o?��;��:�=�S�.�&��$I�?2ek�����1J���Q�����m7���?ʴ�0uk�EG�\� "<��zb��w*�>�mg�(�Ad*��5"��Iv���O�f�9���r�UC�(�B0F�D��r�����Y�ƅsg0Ywh���|�g���k�u���+$���-\;<��r�p�!�H���(Ǹ�����V��cFZ����C�L�����o����/����C�a����_��C���}+R��/��n�Y��H����WH�2ud!H��'�� aB�"`za�^c��zGt� =ufR:�u�����@X9�	<�ovBO-:�Wű�g��J���K�_F��o���@[��N�����v�sW݉'�*������ �oCJL���F'�G&�_/!%ц��jeH9�8�Ҡ����7Ǟ~���Y���V�9`B\���a$OD�M��955�ع�Qw�`V�g��Z��~��L�X��h�0�[�*
�f~c�A5C�#=�
Y��d�*&�4�y�n/O��ByOy�fjŸ<ٛ����D�}��4JP��8�pq'۝O#��5p �'��B�>���0�V��g��m4�q<���26J��$p��j�q"�V4u���+U������Ks�o��B�?�4z�h�5/O\-
T��*��6�>�/�K!�*�P�ݾcmjqCB!|�-Rk�������|c���ÿ���)5���I$d؁!��X:�<X�Fd�N]s/�E#��� �@��{�,�z�ͷ�nvv�4zXTe��mm4� cз�jT��
�n'�v�;IX��_��Îg�S���5����@?�h;�Z�sWН����8��U dS�tX�6K7�x
h��"���'�(VI&��?��KU�px��&c9ιW�v�9Qr�{�����de.�*Ĉ��4:�I��0Z�k�������
\�Uy	�1�Gs[���{�H��5%A)-�o��)�����_��U����/q�)C8�=h*2�m��Q�������\o�!�v��RK�4qc�?j�Ij��Ly���.)�^7.R��
��z� �i]�3WCȓ{h�f��2F� `��!���`��ۧL�\όI7�{Y�E��O�-_�?�R�q�`,��HK{���(щӧ�c[��+����;֙�������8�1Aةq+��"��؏!}�/��i���"�v$�k�%���45oW��6[֖���RtX�KY�G�����jQ��c=Ja���\vtЍ��C'�����p�>BZG��O!n�aO�1Z��L�}�Uɩ�!�Yd�C/I
��0Q5p? �OA�u,���<��f%�M���
:6\��Bj<�ǅ�>����vb��M{.���9m�TAdDa�ﰘ����8e�6g�r)wc"��^p?|��<���NU��g�݂|�FvNQU9�H���7�~�9 �_� v ,����ـ��Uyc�+Ց����e�s܇o������8�081",���2�6�㢇<3 ����4�ͤ*N
�5-d��i�"����k��[/�zٔy����H1�����a, �RA��
V�e�����\ު�։�ڤK�#����i��� ���o���Y#*�p�2��K���f�wD��j���Υ�*�!n�*���v�ۿ��Z-Ic*��e����梸�kY�|���R�����D�	g�h�����7ƃ�`�O��0,�Eb��8�Eqp��W&�r!��J<�U檡��s��8�ם���x��n��[�p%_�o�L��J�l���{�n��{H�� U���:i� ��tC"��?ݾQ��KR�Ӻ��3�K!]�i�%�����5KՆ`��
|���K=�3�`��Xa�9�+'
;� o͓�(���u6��$�a,�1��;�=�E�5Q�8s�E��?�U��<�Ͷ��ޜ��l���w/)t��Aё��T�'�W�����L�#�G�.�Kp��T����d�sǈT��[B��@��<ߏ��7@�|׏��OG7�
$��'��=Ś�,����LP��m�6Ȭ@/P#�t�A
���PǦ��E4��w���0x]�M�(���so	��z?ԝ/�У5r�S|��?���g_q��݉���g7��B�!�x�t�W��d�G/$�.�wŴr��?Ŋ�r)��ALv�U _�K��C.DJmA���%DŽK.�;f���]��P��`ZU��^g}� �2[ݩV��iK�늕3�����BOܬ�rz�`Ȱ3I+<��L�le����_0pw�(w^�+�������S���	])P1�]v�׍Ar��F��0� (9�Ǣ��<��� �MΔ��
�Gʣ�&�w-�!~v�!wYX֝�����3��	ڴ�ټ[�0|�8�k7��[%4�A�p���fA�AV����\�lb�z��Ԥڐh��q��xƄ���j6�קl)M�V�/.�� s��_K�u�'}�?b��i�H}1F�h{��İ\=)'\�:��bH�&T�a{	���كf��E���� }�P�kgI� �&�縅N��"�;����n	tR��BG%F�Omo{�$J�҉��s�G~�vj�"���.Ul몀�	m�ajG.,��j�d,�'r��s0�̌����Ym-���1.���RKp� ��N�)���KQ����/��w�w���Σ����6VD:;��l�YW�cP�"�:�4&���i�g�,H�o���t˴x���'�v�u��:ܶ�*S)����+&�C���t��e���*ijh�.�MةF�ֿW?2i�_�Ö����=�����_L�e����)��vH�U�B�.)�\�l ��)�[��~�|�*�(�(CZr[.44�~��-V$	m�:0�xA��?���ħ���GM?܊uo^�4�GBV�^Fޫ�3����Ǧz F�I�@����LXu��l]E��ώ}SC̎��E*3>I;�P)�i�ƖA���#н��A�@(���� xI?x���P��~A-�J~'���=��Mb�2��m00G��ע�I���8h�	$�G�H��Zz�Ѯ�7��Ԋٶ�7��������Ͷ��ȃN�T1��L�^��وf�}�:�Ȩ�4Z�Z�=݋�������P��#���Ҡ�h`��r��������P|�pw��X@`��+D����Q9�]�ߚw��e�$���6ŦY�?o��dJqh ���*��%
��T���nvB�F�E��ك��A��Ln|.o3�7��c�&Z	�~�ht�l6˲�|"��zI"8�9�<v�}x��wP1o�Os�4��D0�l����pd��ཬ�Ъ����;�i���O"D��*�V=xK��_YA��Q�1�0>�X^$�U�An+G'p3�&��UI�P���l9���U-s'`M�������G\	v2�I{�7O�>�Лd�"_�zD�[�ۀ�T+��%3�V���;���=�3��C)v[���}��P6��gT*�{΋}��d�=��W�g%F��m�.�.�"<={Ic+�aaB����Q-������~t������Z���Ŝ�nC_�u&�����1~����5�$2������YՓXjI#f%���tFы��jZXKR��WrrT�� ?�o@H��Ə)�����_~�1�$u`07�߈��y�@���ʣ�߱��am5��kuԊ�<�N�2,�4�����.��@o-���2)�9��9.`h�u�}��[�xk�$� _�f���Ju�?�h4-�BBv������0��5�n�7,0���/>���%F�⃳f��Vy�6���3tb.�s!����i�
���k�YԑS�a}s�P��É$^����#fQ����y6X�S�ⅼVE�7B����q�2��l~B1�-/_0�����([$/��;�G���6E�Hrzj�Cw�<&�	'|
���������;6� ?ԭ�f��i���Բ����0�)���	�_Б?<�w��u�fb੭h��ͷ[}�g���y��4�Yj'-h>��VV�TI�Є��Uc�T��	����Q���d�\a~Ա5��}K�����"$7�gRlLdg���>��e��L�A�f9�ؓ(�?��sm���ȴ}/K��&+F�!C��lA���R͍3�>�N]�c*��W��3�_�y�u�=b�H�>�l!���~��IP���hG����;�g7$s�s����I;�\�����H�/�q3��Qa�"��}<��&�{Y}q��N����S�"�k|�>XmS�W�G���>:�`���c�vj�Pq�K�ĤHV��xV�FSQ��Rv��P��|�D�E?3�H���H�ۢ���܊�n9��;���r�U�������.�0~�P��� ��?�vg�8��Kd|?��K�=�$��qT�?�
�9ă���
W��F΅��Uu��Jv~ �y;�k3t�ie���T4m/�"�I3@�-8���o�ܘ�/�g�D���sn2���5���d����vev��H��u'��'�V�Z�A�I��ޠ�4VAӴo{�UR�PG��`�
z���t�6"�P���6�VU�R?y� ��y>2�UV�)�՞p�0�I}_�!�)?��eT��}�;1��Æ�e \^����������^�  �h��m�I��׳���b�f�̊�A�`�h�tlv��ɑۡD,�q�fE������{�����>
_���b(��>��2�����#r3n1T�H�U�_���}n�@����Cˣ��^��������/M��őWs��/4�lCVI*<��mٸl%�*���bP���W�WMvM'�ܶ-i� =�z:Y�I8qN���\-~$�/5L�˹�iHWndP��c*P�CU��v��o�K��pLc~�.��a��N�{;0�5,a|/���������Z���ĕj�I3�W�d��`ui�Rr�ƌ����ApoE�s���iO�_Y���0|V��h޼����9��$*�k�QjDu��J�j����}Y �e��>�/�U��y��c��׸l�����й�e�t�U�����������Bi����c̖{�;�\>8kd�����p��֒T��j�%����u�~��Gv��؞DSJ���z�N�YK$n�ȩ@R?�>�h��wߓ4�} ��1���.^	�`������3�f�}��C���:����+�Q�5&�G g�=i��� (-��l�ǩ��ݼ<�t�:\-	�!�\�ݰz��ƃ*7,�`����tQ�/<˵K�~_C�wZ���o�#���aF�x&;xO��c��J8��v�zsR����ka:�Y0y?���a��l�I7D�RC��s)�D`"���vպ� 2��(�Z���i�(HV�"��vk�{��V:MA~�z�,D;մa�/yz]��ɝO�^�I�Hrʢ��q9��]��/�	��h�']�Ӄ��I�# r-���4+�Kvfq��ƵpL�\l� R�0]W0��v�&�|���n8U����d��?��݂�h��P���S���:�6�3�;����HI�U���M¦ـ���`���#�&a��hǅp�I�["_�s�c J�ڧ���x9��˛8�I*�f�~�	�J�]����Mt�ԨپL�F/9���H���������-�=R3o��R�]N|�^+��ȋ��l>+h��J/���刊MJC��c�t�2IU)�}(1|�:�<]�>$m�OEbRf]Y�VoC�8����tqb���{�k��2�݂Oz]M���kW���	�r����P�Y�}H��*�z����c}[��o����������'	wC �ٱV��ɗ�����ggκpf*�~�K'*�XU��c�P�!.��C]<E)�<ĩl�/u�9O'55���VY�]��-�j�4�p�\���D��6B�#n����Q��hm�n:�/�������;��͑�b���������������x3�v`��1s��2�5��H�a)��@�w��o	�T���0?k����J/�Y�D��&G`m�=�BD<-��}�'&���9eg_���VAa?!Ĵ���}[�.3R~���XCY/���՞9�Q`;����p#W	�q#b7�	aU���1R��V��E����"ËR��yx��5�(�x��'n�l��%��\��@f9�9��L��Xޡ� ��h)�����LX�j���a��8��ݲ(7�'-TT&�������w�O�.�P��57�Y�,@d��������/V��,q������s6Z/26{@G_]8"�K���kp��+�$^��'�
7�����k^n��ܝ@u����+^�3���7����ntMϵ?�������Y���Z���� E�T���tL^���ɍS��/]����B�Ҷ��k�(驁�٤�2ϴƌ�Qp^G�
+��p����<�?9�%$䛴ƥ M�뫭Uc��oQ��!��Me��� &�@r��'���r�r�L��_p8�X�mD1"�.����ʠZ��Sv�Q��Xg?��+Вb�`ް���!S�)����J�).��6{�Ё���us�ԉ;�
�Ȍ%Lne�Oy�ڣ��'���<K�S���@�[�&���*�YJM�{�r�S{�n2���r������`��D�;E�����
���F���^�0����J7�(�v[[�@8���v��򎔮�7�F�l�֙�r�7~��i�K�p@2k��!O�F��~����+�Q2V�k�<_����@��tI���4R�� �j��6`|p������{�M���S�6��K�HBq1fd���	;���D|p�߃�֌A朢����j��`<HU�g��QO��>���L��;Y�@�oxQ�I�|ya>C3-���� �ƍ&wz}w@*4H�h�8����9�<{��l���FWJ�N:�K�ྈb��h�c������r��*�`g3o�����}L��"�Չܔ�x�Do���"�A������n��B�{H�r������?��]Ep�\c?��%�h*R"�U�r���B��8L���W~��.������T������B:�9FN{�T�����75���5)ϰ; "�h�g��|���0�&�Hؙ�a�7���yF�9��4����O��B��A����vy��Ðh�����w51,�8�k#�򐜺.�q[�O��"��ý;��pb�����bz;d�H��@˸��'P�	�3]�����<��¿��glkI�a����P5�`ĸ�c�PڙW��� ������uM�֠�1+����C�7R�(���بl
�4\�1�e��~��1����)���q:�9�F{' �NG�kԹ�N_8�cFۡ����s�Ӫ��Dl��c�����1���[��?�y[b(pAp��F�fE��h��iL�^�E滷fZ�;���V��2Z���)������Mz-6�M�ɔ~�.�����߷+��LiN�N�.%��:����)�-�"��d���ЕZe%)LS�(�S�5�ѺAt��
��	�z�uK;�۾��+���3���1h�7�xnEk	=ul�ōk�C2T�ׄ_�T�@�]�UZ�z�_�KM��֜E5>���	Uƪ8T����`X��o�ܜ8���$�A0{��i����� ,x��3Et\�@�Dg�������y�e��w�v��`��'��43&�Bq����?u%t�44-Z��%��	��c�斯O��	�s�p�ŅL����")���r3��F�V�Z'i�Zl���b���2c�L�����T�:�o'-7"��U �o	1n��|���x#6im���f[(���R"��,���V���T�����X ����N��l��J�<͝���޲��LI�V���ye~��c��`ě>]7��2�i�!���V�$��e_�����(�0��e��9�KS��%"s�ЀP�p0�6���+���O�Q��k4k΃�d��A��_.�q�B�.9��-�m��8ƀq�(d��s���ݟ�X���ާ��mh��:���Xy`��^Y��hɚ�y;��\]��
�~BA�R�vx�J,����.90�Ք�cD�����a.��*����d�4tJSv�t������J��`jޥ}V�ZV���i�A�+��k  ?�Q��F��G���tՕ��@FÁ��2
Ui�h��[EҦL)l���v=P���f/9m�ҽ�	���W'`O�3ж\(�s3_����1˗�Ϛ�Q�G����Y����&K���7���B�lz�I�hi`ଋS����I���F�/��Za9!y�l�=�:�7^�e�1Ĥ�4<ŴI!��"כֿ<o��
t���Î^�y�n�i��1�-���t�8p��V1O&�x�B��UN��W~�P$�(H6��ï�@�/*�	�#�b#V����)�oVT�r��+YKz镛�)���9|��zĦUa�fC�y����"��\^�eZ��A�4N��.�^:�Du��n+3f@:�e2�^���p�Ԧ�8v���*w����^�ZnL��BY�*�m��!UK����6���"�7��W�r����S+�D��&]��f����x�&��	}U���R�&)�\��y�j�
��7��Y�99�å�Y�E�s$a1v�%�+�-�t�X1�s��)^�Dp�ǃ�%���M���}a��4�+!��R��)e�����T3H�P�bGE,��Q��*�3�MSR�ZW.B�؞�b7��P�<� .k�ǭyP��t�A��i�z�%��F��T���(]T��LL������A��h~��~,'W��?!��|���/H��	/�nS��`�7@@?��J��m]�H����v���S�|� �
8lpS��ᜇ#Ĺ��k/�6�#��߯�Ǘ\ؖ]$�1�J(+v,��[�o-9����y��0�����جb]r�+oX�uwU��
��r�v5�uW`��7}U� /xs�������[���|W���3�rU6���<��+q^�)a��M�θ����k���^S��L,��k���:�?�lY3C&[�������yUe�i���ش��8w���,|�����!���ҽ����^C�����6�yGCW�[1����4{_${�Ӻ�Ը�y:F��69����o)��j�_!��u0L��:�������G:u��}H1vV1.7����
�wߝ�;�Go���$w��d��7K=K'���T�1��9�_S��vQ}`Id�NOTƚ2��I`�횪����nP?>��$	x�/��M1`�im�E����4�i������0����!��6I���q���>tu�b�f�ԕ�\P!��U�y�/a�q]�!��\Фw�K��J��9���7��iD�W�v����$v ��+u��1��t����h��%�ɋ�,�]T(�cD��-����j���2�َ�5崠���zA2)�qGG���R�Sk:}� a�҉�Hsh9R��[h��j'r��\�
��iG����:���(��+�.�p�?�m�Z=��zb��O!ăT���N�J�ae�I�p-w��'c�Դ�����=�16���;8��&�����aT��aC�y͵�B=���?*M�����h��8|��Nb׍d}/M�|�����F��f�%�<����@l7�=�a��h�Cn�=�*D���ZPw�gG��g�j	Ҏ�N�}e�����B�F&�����Y�0�\�"~��eQm�Ν)?�S@�aq(��tȢ�Ii�@wǞon�БS����V�_�zit)��N�c������3��X�EȪy�Z��������WDѷ�(�5i`O-�r��X[�GY����#��b. ,�T�ݿL�$';�p���pb�L*V��tfgw2"6��7&v����wX �6�5@�<�t�(�k�����>r�Aƺ�.x�&\#Fєa�)}'LW�.li�sӝ���T� �_1o���|_�> 2RvfOy��H%L����S,�0,d��m戅����1/��u_�ġw4��K��ʻᰤJ^?|��q
~?hB�.��k��h���07 \Q�>�v�6x!!3+ף�f/�xi����8DXO��H�� �<�Z��дӈ(��G�\�,i�y-��Z܏�;{�Ws����$�(��_��ō%R���c�xN�9ȩ�XξT"t���(\
;aS��������ɇ�}��]���Cg��{����8`����,�N����o.�?c��͖�t�rj�U��%U��/�I�[�[W���� &�и�!��TO�/�]<�����/UӀ-��p��3��*�B�`EM���J�3/0Y��l'S�3�W�kO��g��7�wm���!$/h[BY�L���5�H���u	ʵ�Ƃ��� )�R�&��c�lPѯ@ 7����k�hl-C�s!c���e'tV��!���,_:n���s�r�`���q7���Ւ���������U�Bs��/?@���t�+�/����NKc��h.�QZo�$�xQ�Y��5B����딗����f�'��@��J�w#A�y���U�{KeH���8�ߋ�A����u�	1}�x���^���b�r��4 g�䲢�RLaô�_<�z���5^��i� w�c��O3z�V��?���b@j�C����Q�H�9�(��o�s ��Ͳ��\�2HL#��������,Gz�����ud|�1v�S^���M�J�����[X&��t޿�PzF�~�͂�� E\9��_��Eos��ا+焩�Kz�!W�9K��z��j`?���MêM>R�a�^�CN�2���m�SG�O�Yn��m"c�b�b�[
ܹd��|Nr@hI��~e����)�&����2�2jh��)��s��q����7�Ӻ|�6%q:�s����kն�2�6J�?�#��|���A�ϩhKt�k1�]x��f灖+�^��/=����e��p|�fx��N�F(<]�1�1t�[p����x���j�"�dO��	��I�1���[��'�Q�Tj��a�k��s)N��J�W�Ȫt��,6'�-�@�6-a����䉚j�[xJCw|(�do�u|�@cl*<��?ɳ8�`ުC+m.)�r����v��T�{�D��Y�ѩ����H��{j=݂�Y���o��)�w��Y�Ik?c�k���a��F�I�u��
�no?�I�k}��p4x��ż�	D`��	��N(�q@h7~	��R�G���1�qQ�§t*i�qD���V��)�Q���p��>7�[���KG�������M��ަ���镘�:>};gz��.��F��v�y��8𾧄�OG���������L��n=A�o�M��
�5[W�j���8[���F1��ˎ�FI��=*)>�C�ɺ���"�uA?R��h�q6B�����!���ǥ}��F�YQ�s�o�N&�ߝ�Y��?�:M���xJ0��~7[)ݦ#��::θ��8|����P�+���rXW��f�J�f'��8I�>�c$A�tr��"�K���,?t)tSRk*���MY>_u�̈�P��k�`R���{���;/=� }��D�����Sʎ�QC���I]f�C��Y���򼻜�r�Ћ�s�\Z;���)�A��CD�������|����ug9&��9S�9`�Q����s�_���p}z�����ҵ?о���G��?Z��?�G���D��ɻ(���al�9S�nژ�1�i%�d��XZ�`���Q)5���M�i���4]����,g^��`�$K�d��������o6��5�r������g�z���*�$�B�<�\�5�h�0�������(��.uF^c�!9?أ�yC�K��&(<�	G�9]�?��0���C�X{a�L�o��A)�׸��ʤ�8�v!@��SW�~�=�`�f�9ܢ���&�~�2�Z�Z����Ɨ�;�c/�9��:�v�<�7;7Yt��{ϯ�Oz����6g;$���?��~��#O��#X����jE�b~��˟�R� 4N;��FrX�W�����ݩZ
�p($�����	jw��t�!��;p�r'+��Xp�a򰄯��T�)7�.8h��IƌKe� ��XF���)��K�x�j��>�W�)/[��5�nͮ��1�_�s��k�JnL��9F"L��;a{�h��OBgI
�n-�Ϝ�d�$����lgH��sK���{�����P�01�i	d�7n�f}G��T�]8�*C2h�j6kζ�a����k+l�zBA#�����M�2O��M�^(h R}�i����CO��HPL}��p^��_��~��vxP@d�fs��ev�غ+�k2�����Fx=�#:瀇QR4�_�l���,�:��*�o���~�]e`498^W�	��ÊhJs�c�]BMNf�D�*�Ͻ�K'Q+N��%9�I���D��Z����˅��.�cay�;0r,���c�լ�	:Z�z7�b��!>t��H�?ђ�룢n�����B��̇UM0�� ��Yr���.����W�X3��}YQ��ĪA�"���.��%�>�/�Odex����e��@w{����Lӆ8n<j�y��G��
%��&H��Ǹ�9v�>
���G0/N���j��ʄ5ĽjG�L
�'�ͷw�'j�)jY;����x�!�9Md�*���,����PY��<yɮN([���x �AacىV���w2�� �`���i�B.߂~�+	ϝ���tT���o�kF$&^���58�cZP�&�k}v>������j�3��x�����@(�3V
F8�(�L�\�K�*�2o`0�����M�	/X�SP{W���ȿ��#�Y����(�A��g(���R�0-�e:*ߋe�T��H{7���	�X��o�k��k4+dC6D����_f<>�wIՅG�h����s�=N{EN�����X�����L�u�Ę��R�'�ѼE�Gb6�?���h_@�"�o��VnMHM��G���Bg��)Z��dsW��Y��h�xK�e��x��K��v_?�� .Н�����:F�L�a��Z���������9�>H��|�[���*�Y�"g���3�H�:$��������5�A�;��1�-�����_7lm� �Wsi�vXT�|�6��>V5!��o��8��j�8*���aM\����@�c��û�Gή[7ٜ����a*9䱞	�lFZ���eC�����Dr�٪��,8�՚��jU����a��
�(��s`t@u�����U��D�#樊�*˖������*#�R�Z���d�_av�|.!�4�PK��cGp^�#����Nӳ�Se���a���g������"X�SIq�އf�\�a)t |j�2��+(C�Z�JO�'H-�.��ٸ�Wjk�vND_ҏ�m�^MLAt�i��3��c�X���yE<3�Y(�B���@��wq�M	���k=c��vl~d`��~����& �!�X��F6>`��_�ٶS��I�6�'�W9�-Z�I��ʧ�ܙ������y�W�3>�l
�\�+ۉ���2u�$��Y9:��>�t&�7܅��E$��W!,���w{��	Q���6���p�HFN3��FM�p�}w������:̉.*��0W����CGlL=Oϵh`�եr�Q_'��r*�|a��#i7�tμ�e�ݗ�Pb�(���B:UŖK���c��a����*���6�����z�r�C�u��N�G�(�U��cdB���K������l�U�CgpԀ�g�����*_X�T�s,�G�]�:zbm�����V�s}@;�c������i/Tc$V��� s�n�t��W�&R�ۄt��Mo�sx�� �� ����	�ީBޏT���g��q��u{r�V����-+���\��aǸ�o����ϯ�����[5�;�4���09�c��DȂ����Df׭h�>O ��B1��A�d�\`a#ۇMbx{���*���[e�l�	��jBԼW�~8/ �ǩڂ�ǐ���ç$��oγ�.z��ML�:��g��{�(+�
�"2���Bj�����j_p�,�S��,:ͷ�XR@Jd�^�bمb����0w����y���!���O�{�Ba�fb��7�;����uy�_*ϧ�z�_x�}��&qw '	�&N�����:��J�W��_�����a�H&������K&D��+n��m���Ŧ#6  �R��A�؃/�#$�K� ��B�~Ĥ�7S62ǫ�;��D��5T]�gE|�� ��֫�\�R~aO!�)�V{ϐ����A�v���}�;�ܨ��)�5G��h�6X!N?r��[[����_",�a�1X4���'Um׹M�)��1v�u���uގO�5�]�!�����MA^ĕ�i��@^ϖ�{���U��Z��3���[�n��b��6+��狦h�a>f<��ȗ�<��z���*��f����At��IA�G�Ft�m��|��G""r�f�A��)����H�k|J��M"W v�@];�fDhQ�r 	���lI��� '�>?���bv9��хILk��:w�?$"�Z�h�����3l~Q��02���%��$������=rɰ~O�gy���IM@�^{Ǫ�9���	��<I�%�~�)�"Õ��N�-�(�;�gO�vd�����/Ѐ����̧�	�J�2�,]��\�rJ���ԟ���P�v��g�~ܑ��ܺU,${o�Q���/b�[�]k��zB�J������(��>��I��+�r%=:��;kKg�w>��+4����?�q�ӆ�'1_r�tE�����5���y�c5��`zM��pL�ECL�o��.Ҙ����e<U�uk�Eb���%�%�$�|������ҍ �-�e���ix�;�=G���H#D����A�OF�u�:b�iR<�:]�oX��@�F�#�Y��ˑ:ъ�"�d�^ls�y��Gfr�r�>���a�tt����	�)_��`��%Ԓ��@��>���1��$�bh��tx<wD;��:����%��&�#�U&&:Hc���Xt-Y�j�:�I9�#Ng�$6��5WK��v)C����	��,����&�Nx7((2�΃�l�7���X�����+��y*���%���
�f:�?�텒���ok�\�K�[t��Ӏ����)����8�!�&bQ�λ';\-�再O5�7���x�D��_�Vo�۪Ԃʒ}��m|��AuBU��\�(��'P��>���P
�u>�瑬`g&#���3Ց�����-iG8��@�M���6=�k�Z�>��PE��rmLU&�غ�;��½)�� {A���c2u��M�g���I�E��V��\*;��I�U|	w������!]u�R���V!��Eʢ��ev.DA�V�]a������Z~��~���	�ezp�E�΄��p�D��'��](���e�^0�L�[�w��5G��]�_	K�r��{������+�gJ���(>x�J������i^~԰��!FI����ue]�@}�N�X�y������K-$����.1l���I'�c��H��Hl����q�e"�n����ֹ�s��<�V:���#��2�4���4G�$�Y)��=�=�\�F�0�hM�R�9�;�+�����Q�c�r��LF�u�F<o�)f��x\��f0:�7��{���Z+�Z,&E�GR�έFGL�F��,�3ѢUO9f5�#�J"}'���^�Y�2���Y�V������5�"���Y6H�'��t���=C�f��N��榳>;K[�O���G'u>"%5J�o2�0���:O��ٳ_��C�"�y��
:����iUF$���pALن�۝�*O�ޒ��P�=�/�a��`���A>�ۭ��d4A'�%[�Ik�#! �i�ǓC��O<7+̇�@��?��
��y����p= �����P��
$�����*x��_�-��P=�H�S»ț �6:7#VD�=S��3��:�������e0�j�[oR�Pm
v�(ă�A.'��@0���߻���\�������G"��E�n�Ӡ�l��5 F�w�K4�TI�{�٧eE��w�/13.]�%��@B�Rߤn��j,+T �`2;FŐ�q$��ޣ��x7!��E��6l7�����szE���h����G�,L�W/d�Ӯ�g���P�1�P�z��� A���Z��s��/ɴ���q�Y�q޷ rfG(�`�?O��Aނ8 �{�r�Pu`���F-,�)��{��Q~��ǂ�ė�'��NZ�k¡Pyį���i>�9�}F/��?"
�N�AeǞ]�7]c/5?r��� ���8d����No�v��
��:t�s]O�P�m��/8��5nl��@����LR�
*��"l�����M+Ж�IP�>㿤���[^�c�4l#4r�;����K�@�xzc�O1#��+�s�C�x3sO.:F��޼N��R�w�n'u�'�v�'�	�v�vU�����4�>Л<�
&fEC�K��h��t�}Ev�?,3�m���RL�̑s��,yw�J�cs�6A��7�t^���\L�Mn�l_�N�J�5���ͽ)�T1M|���k���~�8��qv���#��ƈ:�N�2��ϝ}]\f���z���#ZaͽK��Z�~.mKϯ�����6ޑr9 �!��%�}G��^�ؠd���p~�m�^���,