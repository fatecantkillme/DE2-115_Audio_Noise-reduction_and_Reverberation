��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<Ph���כ�� oҺ�����5�B6���JiF��?�;}�xx�>̜P�7��&z�1~����w��k����?���m��yn�f�m},���D��#l{ b�?b`A�V���ՕD�(�W}	���kw�?��t~�삣ՀB��y`>,��+�PW�Dv�@�7b{K�uF����$$E��;�zQ9hV�s�$#35�e���s
*�'ǝ݋L>y�勱0�3�a=E"
 ���Y�j��]{���j�2?�?F/He�(�=���(2H�T��O��C�s`}�M`5��_TU���C\��s�	T��FpgǱT�tN�!�lz�r��x��P�])���5�Lz��m�V���jm۰K덆�B�S�^��2/�;� r�"h�N:���!�0��l��W�z0�8:|ɟ�߄q��q����:Z6���ƃv�����4��˞�Q�F����o�ȗ5����~L��\q?��$�{i1��k%��b��HO�Z�dɗr/@ѯ(�[�A֓����~36JIg଺_�S`�X�.���#83[��$���+z�LFp]/�zKw�ߡzS�t�v�����.�ݲ�3a;��Ac�\al�yw�K?�P��Dh@���%��P~X^�)��)�a=�,z?�4�VD|��Ym�D�y����[�,��X�]j�h(�s�V;<k��zE�-s@U�+��?�I;�kƐ�;�f{���|> �&��
��F>�P�pm�m���x�(@uL�۸�E���	���0_���ۈ��H�Y*kKB�b�ϋM<θSGw�ɶHw;9�}yZ��X6�[p?o�\��㽝U5��=9��oʅ�G��� ײJ}��Lq�,YIЉ5�.��x������s	z����rSX/�:m�9�KA��y�-O�Ԗ�G�#�W��,�Y ���4�(b8G׈�":_z�"K�������j1��"c�N}܂^e37&����!�f���J���	m �n�� G��Z�ג}�\�+��XvW�<��3,L�������dǅl�=�9�g���0�������R��Z>���/Q)�v{􀾊w�S�i�Υ0�B��l	f�i��/�ކ��,����@`?G�Cu��}�8�k�/�o�L�\u��J7��������٬�����M��9�7C�<�1����
#�T��~58b¦�@�f�^���Bb��T]&%�=n�s�s��A�O1�`��8��U)���W+O*J �d!ۍ�x�$�cL����ܪ��zEtˋ~fv�q�>&>�t��_Ţ$��t�4��O���-���:0�zբ�;������R�NG�,��ІE��F	���G��zSɎ���7)�{}�η��i�(&��&����(��1�0���B������9�iQ��W��	�B0��u�g($�!ZL�����+�/I˰O�V����ʉ8hWҕ.�t�uߜ\e�}��(���|���Aj<�2�%����Ok[�(�_(`��S}�O|���ǃ���85'g�0P��ލg�N�����A8���U��Z0$��\�췪B�P�iVh���ur���������FK��91?���Tr'w��|�K�O�Dd��Y ^�qM,���t���z,w��>����<� Ҙ�_Q�:p�w���̆1��=~%& C��U�ܤ_V)�9~?B���I�h.�B��gAEXFNӑ������L�a��;��L��!7F���w���k�<^���)����\jv��'���pqf��	mc��57��?����t�� >����v�O�����]�Y�~hU��M���p�<X�����%�`�|�8%���.��^NT/7�;$ʤ�d�{�aK�Y"Hhy�P�}X|��7g�NV�-RIm�>(�����j�S�X��7��#�o�'(ƴ�S�@ ���Xfܟ]s��'��׸27n��J�HJ3�L�4I9�|��_\��b!�Wkz�"�d��n1�A�6^��g��(*y�p���m��%�	�efL*\�tN�*X~����+��BfS��9�	��v�؅��� �G�1�䔻y�ȠU���.�ϭ��k�x��Iks���p@�h􋡀��:��T����*:W/����ސ
�L��ͻT���Ql��I��[��z����x,:Q�3���m��Ʌ��Tߖ}f��l���hK�u�`��	ͤ'	F�(�e�#�]\�i�e�'kr7�#�� W��!A�R���9������g�D
V,Ĳ�S,9i�$:�n�d��R2Qٸ��zj�߾�b#!DPǗ�w��iv�C&w/x�|#�1k⨏�����YM<��7���<	M*�l��W������t��ޣҐ&������ �9R�]�y����7U�	�k��2"Lt��擔�k�&1=T��-��,���4��ɖ�,�r�,�ZF*'J$g��U�b8��z܅V�1u���qq�'�X�)���ُ؈�|��~-���!��ͥ�c/�(I��CX˾���qM��0S��	Y�z�ы���6������r���2�v��O�?�5�jr !V��A�4�G�����
�)�_Ϯhv�ծ4;��PٰI�H¶k��Y����"͎��fQ��.&�jW��1�+$���������GV����:7a{b����6"��^{E��[坱�+�����^��%"ņ�Q�2����Ӣh(��ՒWC)͊��b�+�M�38x;�d��å������2.��V�Bh�W��ԏB��I�k�ͳ���e>�nd4�q����VMI����V��Bco ��?-��J:���΢���e�*�J01<A��Z���.(�԰��O�}ma�Z�+�jr�0t
_�7�O���� ����uJ7$tܶ�c�'}TJ&j�]SG��b8ҥ�a*τ��uu�.��ݪ����Xc�5�?'�T � ZKÚ��%rb8)-k�L�5b}���ῒ�_���~
�rڿ[�n � e�9�tV&�c�����<W/��P�z���7�
|�j�u����K�!�,�Vԙ��Z������C��=�� �A>B�}��5��D����ϑ¬4���=a���Y�v�~�Kl��m��.ǲ�ܸ"T����}�,��ưC��h��
5�K~>��X���� �a�j�
�DS���@p����1�YL5m�Ĭ�h�R�`{ߠF��-�%���ւ�? 
�ռ��,!)|��\�:�1��y`��v߬�, ����4�m�C�%d���E|��x�&B[)��	��F�^���CH�󬋋7�^�"��rM��"%#�2ĎZ��1g�ϤLQ����@�y��|�9�Pv�655>jT�c�q7��l&��J�R����Ռ\�&�Lz{dڜ�GW��+S�I'����}Gg��{�UK�������b���I�Zj��b����>�h@����<���^��Q1�G�		r��&1�g���rpm|E	ݏ�X��Of'�N�o���k�6�(ƪ���\.B ���<��~��D[��o2��n�k��S��L}�a�'��Lh�i�`��N�S�e��WMW�"t���vB�_�"E
�IGd��̅8��~׸<��p��dF%g/C~o���=p5��Wz���&�؄�r��Q�'���+ �����pbc�|�[ɏ>8��آT���䍰�k�'�ӘG���"����>Ing��3��3�0 	fT�>�Ys����[����KP��_�[��o=���]�����u�A5��d�=���]ZH�T�hx�d0����[����e_���:Y����w2w����&=y6w�kB�L⪤o%�5gZ������e�|�*Ȝ�a��?�7�}&w٭���Ђ�-`��s �,pz_��0>�i���6��a�M���p֋��f��Õ��T�u�I���l��Oh�D�+ھ�"p�T�5|�͖�9n+��9VVޤ%~�u��W�����?%�l�%*��v��U;+���7��>�0U<�zx({��/����"�Y���,J����ާL ��d�E��>��̡�(����q���璊��g�hrf�ji�!��:4���Z���b�x���M�(.!C a������5Q�8a籖5��xiy��ڄ)�
�R��B��^<$H�d*��Ո|��c;�ں;sg5���Do�7(-ڲ5��_@X��,6��K�Za�(�eJ���(A���݃!b�|�G�VŘk��G�'������ qFW�!I��m�
���$l� SІ+������Φ�zI��l�Q�9`j"[i δ2�b��[��(��o�
�\���k�,k�\w�T����M����|�Y��ўY���$N�W<3^2N5���ӵ���A�_��9���Zgx�!���E�	���[ͣ��S��y,<� <eA��(�!&��g���k������7��
`�t���@
J)�ڗ�\��љTwߞ�^��~� -�J����+�h��0qH+�a+�܏@�G���z�~�ˮxg��?��D:�OU
��"�tϑ�(�p�)�8�%��'��!dg���B�g���\�[o�H�@���14΁h����`P��Ih�=�:� ��x���nBL��zϷ$�!�H����	��@��"�B�7$M����O�[�P3pҕvA�}�e�m�������p8�.�b�Q�VJT�	5*KO�,
���-`�oɈ���_��3����X���}��Y�}i:�� �6$���ؤ�J�������b����'�1�]��8�� �TZ�-(��iz0f��1zb�Q�0�FJ'��h��|֊��4�TrP2%<���Ln�Hm_=��;���R@dG�aê�|f9H��k��A�=,1#�[�$��~�P��
̜#x�W�3G\G�f�6C%�7eI��6QS���2t����+0�9��}�^�?#���"7����O)Hs���ץ�V��l?�{孒&]jLu��������W;�،����N��/wl'���g���ӈj-ٜ(�?�m��Q6��^�=�@��*^�ʰ��Hzd���`�u ���3�:XU0��p|[���%����*L]�������h" �TP�lm1`>7|x	��WcY�|~�V�3q(��'^��Q��=ʐ%�5s���o[ќp�a�ڌR�96q�U	8�{�1��c�*P���U�?ݘ)��7��ǿ �TC�d܄e�$E�8)!��6q�݆�9�I����b�I�9�t��ˢ�&=E^�'��b��F?Ї��&pO|>ʘb�Hk;.�;�S�qQϞ�3�
��������6
����L�e̱�̮Ŕ"X��b?;o΍:ɚ�k��6c�%Ē�WM�I��M$��u�n=�en��敼+�7P��"���܋$>;S��F�\γ�+W�9�\{�����k;��)wU�aE����%t)�
�&�����-2\���k�����KZg�;tR�K	��Us��ڊh?�Š���t&���Ʊ���c����61:>��T���L��M���>��[D���}fN���J�hA�+�J�WvN�B�o���Cj)�^(�(�O�mo}�O^-rh����_�-p���tK�j��2�3�<Hkv�-ܒN�6C��/���ZG��vR2�&��b�:E�s��=WiD4[�ɸ�/�< �?�!$b�D.|+�rmN���*خ^<�}�?�Y}�#��#�M��Go��k<y��
E��m��Y����<em=����( ��iY�Z���%Q����/H�E�\�~������!���v��r�|&�L���s�F����Bq�]#���d_�ͻu���?[6��䟐�ֶr�B�fkW~��<���NJfmnVr/ӡ�Ύw!�7�@W��e���c�%H�Lӈ��A�ޫ��&y1��)�!��+�PT���a�-�s�㚵7���M���c�Do�^{|���\"u�2�P��@3b�}�!�8}�#v�����fm˄�"X�VLڶ�UN�@�$�H�o����s�7T 9����"�"�|�iq�	�]L�5ut�ʌ��@�I�܅�yT��~u\�M@r�)U�@%-�^h���f&��W�(B�1�f��·���-R���5�t 2����+�z�E�s�PԮ�Т�"��ؤtXOe�%���+�e�����u���mz��SWS�%�[���	א��|,� +�����9������~�P��sOk�*ސ{�F�6BѤB���=5��9�����Z��9��
���zPJ ������ѐ//!u ջp�Q��=�͹��%�w��_-Y�H�w+9+E�w���)x'�9�� ȩH.j�z%�!g�6���q��u�$L��4�t<� ���G��d�����eV��1�XX�܂11����ǒ�Y�DA����ɀ&�A���ӿ41*Τ���X�$�|�p@����P � nI�� @7>ޕ������3���񮐘�xvֻ��i�fBn�'�8��ub1���DF�������^n�F���N��!��Թ�O��V �!���J��[�_�?�!��G��r8�R�O�����˓~��S�h�q���JkI��+�O�}7z�p2�-J�Ub����5��1`���-�R$i��蟝��U�[	���	1��+��>T�W�*�(�*�Ƈ/
�lZyg�P��Bh}�[E��c����lCPm�|ޖ���~�w�
rw��N�?�LXmQ��{{�i�����Q
g�H_U��[�I0n���;�ùd>5i�4�3�S�?Z�O�ۺ1@�S(0r)Z��)������6b�Qf����5�̭�n��cOrO�Rg=�$���@J�Ί���n���[V����]�GM�RBKh�3�EȰ/����iDA�)#�-���&츽�����;�۵r�e�Pޜ���'����0"X5����b�@�k�E8L�;���&:����^��Yi�L�tt���W����A҂5uF�<@T|��%j���vM��G��{��HO��I�����{#�J�u���6iu4;�&'p�b��F�c�tC*et�������@�j� ����3�z����Z�oe;��A�Bk���oe4��j�?MP�#^� �?h�0*���"�oA�2�鐣l�y���H��G�X�h7
v�5�A6�u���D��
�*΍3��o�/M�\X��Fl57m�]iZ��n� �<�CD�E
5�5Z*HE�"��jpD>,� t�͵E��Ct-��%�Y�p~r%Aw}(����A^*�T����g��y��;��@O����ܴ�W�@����c�>���[@�np'qB�>zg���0G,CG㴋�=�B9PF4wF���.Y�b���5�l�'&����$d�]������-#�$3r���n
D���Mh� �D'3�Onv����]���ϔ{����p����4=.=��y�Fa�R�i�A�E�z`�T��&>̔<{��;\j�#�3�_�{�%w%��A��7׆�Z� �,���Pm���%�J=��2c�f؍ �4tБ�8��K׊�=�#�����:V��s���/��B��o�>Xأ��i�%b`A��[l��o���5�_n��N��!�!$̒.4��e�p年n����{�g	%�	�|�-���f�o���\��[/�n�8��KIEYD�ݯ� S����!�M�A�y���#��_h3Ҋϙ��>Ǘ�#h�a���1u�;}��kgK� �&�+��K�3�(��T��v��4���k�L�%+��"���3���-���'��I�
�՚���AY�y*O']��B%�I2B���'Re;���ԛ�@��c�D�ak*ʯ`��0#�<k��xb����>aH( �9�}8]<��P�dWK��R��M,����s@ijs���nΗp�}�~���&D�KF�D�6��l2��~R(Yb���C�cꊀ+�W�>�s�ٛu`wr|�ћaa|��о*��#��I��n(ˈ�:X���a�~:Bn�=�K�"N;����G�蘼��]J��a�!��|����0(ӡ����#�,xW���΍m[��À��g�g�%�ݧs������\uǔoV)���������	P8���IJ��-�W�wr��D�݈Ki�}��s�B/����FJ����Vl���o��A6IRH�䠎*?�Qp!�yc�=~Ľ�C��a.�IY�M�4��f;�f�Q+,R@a����d�Q�uy���ʸ`�0Ό��lD�C�oK3Y�,�� ��(�ِiX-���2�%�,xA�4��(�)z���,S��L���-�R�G�.��s�W�3�v���m8F�KA�^�߄4�ѽ�GC��;�HP΅*���mR;Nl�RODt8�����x�3!A��W�失�3{��AVy�������G�W^z���~��t��HhT��m��3���u[D?��u=:�F���	c �	1�	6"�u�S��djq����$���-?3�\�Dk�?Ý)�1+�//�8�(��73��R	$Z`L��96�2��1[u�\�ƗP���Of=�q��Ce�ɐU��P&'�2����QP�/�$�bl`�7�y��ڐ6���s��.����_�u�����A�C�,���t1I��ym��M�J�<!��'	�O�e֞v������ͳ��i�&�kjf�OT���[��à�2)xK�*Of�ԑ�=�s��Z~h�����[`fZD�$��Ţ�S�v�K>AoH_���:�9������< �``���"p���vi "��h����"_���[gh��U�v}:%�Y!��"Z6n����\'�9M���>[��vU�Pp�HSXm^�)gޛ��tmd���d��t'5΄���u���\�����}��w �����7��VF F����0���/�u��w�uS���)W*�T��(�sq����"?/g×�/X S�>��[5�7lO��o�; T15���}.���lu,	�+v�S��
E5��dɨ���摁��!�����j5ώ�G���=�)�-��3�<s��dB�z��km>�As��9��d �ږ�b.��N�n;����|����/͟\�H���S=�R��Xט�Ve��7�L:��<���j�p|#�"�ň�C��f�� @�?�b��q9��}�0�K#�~��^(.V��^̟��p=����?G؎�m|qDɝx�k���w{]�:�0?t��-�5�` ����5�x 6�HjC��$Vh�0�[�=e�vj��ZF�P�],<:kT>1,�0�"Q��Ba(�����������5�ͩ&=0�H�4�#���(pxr�\#ଠ�;�۸�ɔ1���8~"�2�`�L�"Il�H�i��)
˛����٢�y��e,a�O�#JdL_�G眘���ܷA1��^�����ͭ���ڌƌ�1SL�$�i��i|J���C���:�̹m���Fd]�+gJ�v��_{�}O����0˨v�6H�^#k�i�Z��h���~����{��
xU��F�.TuIU	&�7k��r��X{>�xͅbǣi��Rso��'{dQ����Yw�o���7U8"�����Z�8�O����
�ԈKڬ,�ԣ+�6���828+H������ �#���?�r�(s�o�=��Ծ��]�(�5��R*ed�%%	�N�zS�0�4!�rwR�T�Ͷ���c�N9$���?�zO�N*cY1����عv�3~a!9�*��<}w�,���f���0��b���� ��x骅-K�7(wc�L�%�C��O��Z��kJ�]Z�	��B6��D0� jL'��������a>Ъ���"�;�.�9��e�
��?=9�������Y��&�)��G�7������)O��;E�u�^�����4���sH_�8}�-?�:��e�ڐ���	��բhWrx`Kb�ʌ$٩i�:'���iN�%�*{Xs<d�(o�j�����"�D�Q�Wr(�%$�ea��ٰ����H�Wq�蟗K�n�p6�#3%\��w*��.ۉv?.�T@޳O_q��=����(S�=z5(��%�=����b&�����e5)����c�.e8��;q�At����j�)ťr��Q�ɨ(�FM�G|1۝N1$�	���������G�Oø�R:���fepC�x
a���޹@�i�{��?������q&��N&�-��-C!�YU�YL�*|�^bǬ�غ'u}�b��P��
��0����&0f�v�O��wfP�b t͔�Q�3l;}��_�2�[Hw��s��=�K���Q��ˀ�T���BuǶ������x���p����l\Tu]Ƅ�ẙM�D
�"l(�R���_n>,Z��4|����Z�5�?\<��r�̸�d�J��@h�� f��o�C���n��*���Υ9�!g@��J��t�_�XYD\�JG�s�Aڔ �:��A�� 3�y�"$���h�$/��Au�s�_R��1���!kz�����mkpƓ3�����n�&-���TU�D�Y�{��o�b�4�*�O�2|����0��"(�>�����"t��Ķ��\;�7�[�ž�B��8o��8$�߃���d�_��I7�elɾj=6�x����/h�����2tc�6���G�����eI0.NׅP�M��-�5��kRz���}� ����V��L,8�
~�P;����Fސ3���^t)�N�oL��R�=8�%NG�&x'���jF�Q2縜�����+��@�!��33�f{�=����xOLp^��?s��@Q�k<����Xf��?%��.��	��k�g�D��3��K��+�R]�~�s�{����tS�V�� ��5�t��fbY.���3��!�2z17s��:��g����>�V��ψt������ ���4��ϦM�9=J����re���(Y�~,V�'��aXز%�bz �^wMꈵ>A�V��t��
2@ȿ�+ٴ�|K'�m������5��lߠۭ%aµ���N���r�6��A
6(�!
AX���:�^���
9����F�w0&���ⲉ���]#vf���5YN���|Qi�?�q���/�'7�:�R� ��ҁX���14X~A%(h@6\�>2P����b�gc�J����I�-(��΄=t��Y,����C�5�j�bޣ��_!ώHZ�E����__SD���0�n=���g�ՁD>�V3��<��
��17������
��m0�z��e�ǰi����N�������"U�S�̢E;��g��2�����G2ikv�ɍ�U�'u��;׶�~���/��w�����y4�J��>�0$p�K��EP��6�q|{,��Uf��B�7�>qQVb���(Ia�z�g��������_L+s1�Y� ��	���2�e1�Y��g�k���=�c�r�1ֆ�8�D>��G�+.�@���2|��eD݆�,r-	���_c���v�&W�@��=�n��R��	� h�NFVRX��K����}�3g�kE���':՘������F{7�q�6E��<�����L�[^\�1
��i������%2��m���<��j��v�lZ�#׵�sh~������)��qW	j�7P����:�D{ĂLxQ&��䵠�r��#�U#���U9�;�w=>�dF(B�rс�H���M>��<n�A�"w����mL��h�4c��������u��4_KE-|�X)�[��J�%�Ä��n[��ˬℝmY�y�vX�u��O�<�[��,�)�5){6ӿB)G���0^�η%T_�I�0�|�F�0�(ښ��:�y?7y��|��&P�N�y��m��*� �m"ěX����r�=����>ꋍ�~���o�8�W{[
Sߡ>��꤬}p�>'�W%Ț��2\0�ēKS�E��,�{�����t�~��H��-���}D�\�oqƆ�ST<��E�A�,�2Y��E#"-wZ#@-eǲ:�|z/a� �7K[��
E��E���7f���ͯͩ��D�D:�E����b�ɉ��g�-�$�⪆y%�;�`��:�K����pU�9�n��4�6�y�;E6�%��BN��Q�>j?fqg���u�/;uw��P�4��$��]BӨ	����*�%�˔���m�Vn��6/E̶X]�p���Ƅ��=���I�3&R���?;G�K�/-��"�[l�(�o��3[�03����[]��2�z���lϋ^6"}��N�����8�ܤ܂b��F�r�+eO&_�)Y��~�O��E���ifm8[E*^�ů�g��8��l��!>I�ؒ�v�S� s�!��������	kv>��P�e���2���z*�\y���I�+�s8M-��"I�B��� z��A#A+Al=�h�i��~S���kJ�td�~1�H��+�i��&�͏�#�L�'�訹�a���;䐰��V�w0��Riw@���r��)�b/��7��2 �O�%���j��mC.���_�Bx�g.����zܲ��M���$κb���f�=�q��z�R���C87��~�c��.m�ݗHW��p%p���>y��L�
b��|&sp�U���`~L��]a�P���_�|gH�J2�i�-��Q��_<���*��o������:~�1�5ߺ�K"��7�	@���3��V����jK-��^x)��雯tᠪ�v2d��A���6d34o�.|����y�2kv,*p�R�:9V���V�T�݂/S�u��Q���RN3�|(�ev�zu�����
�؜��s�t�r��9������B?����A�^K��C�eAx�报��Q=.�L �){짞D�p�CΊ���9&{��:w#�����1{:EGE�ޅvZ�\G�Y�f�-}��37�=kl����3�qR<l���.�m����sv����Ӭ*�6�f���pX�|�8�8G���H@�k�{( ��/fs�M�{������>5�ɺ�脪W�8�`���A��F��|)u$�~�qm��#=���+� e�za"�����?�k#ݢp�, %/
�0"�]��E������B��Kˊ�n}~�k������yOc�v65�0/�Y��~`1f�h��T�ݭ������)�/:{����E���������<����-5etfLoh X��V����6 	0�h5ݞ��)�ﬅ���1!�F��&��'��c�#��5��>Â��N���.�� YY���U�!�tZ�8�K)���R��r��`��O�}���ɪ�΃FAh*�$#$J1����A#�R��LF���h��/Lyx��ь�+�H�=�P��W�gH��螸ULbU��1������j��^��.ɆXП��f�e��~��AC���J{!F�l��+��+�����KA�ުb/�^B�DS@�soB	�I�:�@�T2�c;�|�7|31�۲�n �l���1�]�J2qXϩ�h���Vo�~���1�Nsm�w�,��/,!��$-՝��i6h{�ihn�#JI�d�v��hʐ�\� V,�c9A˜`�a����xf��G���<O�6$��F�����'�V�o�]�q���ŏ����m��C�y
����)}+t<�R���2��7�rf	�Ǔ4i>����2n6]J�S-мZ����m���K	dݙ�j+Q��`ςO�͊{��H���0��a�,� �;����.g�yۙ�\��O9�6U�O�Hy�`��
�2��B��#4�ɠ�� �wYl����瘚�-F�g���M8�M3rH������eu����ǃ�(��������њnq���5�'>�~�IB�AH]��o@fUd ��J�7���4`-�3N�^���h�F5�s���a����2�i��cg���mN#�-�����q���R������e���e��$��v��-ٟL3�9��î�8M��N �He��m���0*��3-O�é(�N��i�	�˹�z��b:R!͞'����a>4~|�0 ��^���o
����w�m�Șa�zM����(�����v�f��U�b���~x�ɕ��M���M�ch��:ͤ�(���?!�1�B�����aI��X!VYQJ�w����z�=Re��zemi�~��Dܿ�(A�c ��&�*��bg'Yhr{�E�o}��M�:��Aꩧ?����ܢ|�Z�R���|V�C3g�!q�b�)<H�����������rat.�#(H<y���(�����*1�hg���Z�tĝ���U� ��8�i[����%xQ�*�R~�c~�)��y`V�F{����9N*�K|�4[;L��m�$��kЏҎ>Du����T2v��-.�B�|���|�����{�I��+'�HF�h?�ʫ��~������vƟZ1���{��;0Ȝ��y`���g$4���I}xfn�I�*[����q#p�W�>fa\	��z�K��{�pI��'h�����{�} ;��]3�n5&ޖ�M�f](y�+T
�vjA� Wރ��,-��Ҿ��U��O�-�]ƢO&��g�F��^��X�h�OxY[�����i��'�m��w�黒a��S1�<��p|*Х�Z}h �޴�uQ&�o����j`�������1�s|��i�Tk��]��t-���C�1�zu�T�(/��Ƚ�q����:k@�o�Bi���FfUW����}��[�؍>pj����A�2�F�f���m��%�L��f=�J<�iy�u�rm�0�05_p�L2m�ӑ���Br( v�(IQ|ǰ0:�� M6��!�/�nfD^WBk�s�B{�YD ������]6��ֆ�Wۧ��I��øU��Zи1�
"����&�Њ�"�� dw�i����\Oږ-�T|]Vg�4�롛7��~aP8�D�9���t�H8pt���d5"{�;5=ǓR-��^L�����]{��-��H5�Q/>S�>l&��Z��1��u;�]��{�氕�	A�D)�Lm�zG����~����w�om��@��lU[��܊e%@��N�V@� ��?�L��*�ʉE�]i�l����3��n�P[��Ӝ�d��9���:�)��켍y�,���8���*���:q)8y���}�M�ؑ-�F�zl�?*^7.����G�{+�-?�b���e-�J�� `�q3]�j��ܟ:�$�.V�兽�0dO�<���Yh,�a@	��H����N#^�����w}9���Q�6Wm��q�_��/ W��M����w���x�G�̸m��J��X���#|�[���6e��Xc��#�^3�뷃-� ��K�2�p7[K�V�C�S �X43x������r]�v"�=RM��$E�H��Χ��b��HP7��6���d��ڸ��(�%/g�.�l
΁?���8�E.�/�,'���0��)�D)��%3��j���VG�_�Q@������Ljv6n�h��+����r<�(^�p�����������O���h��o���]�|����,v��Q+�����\ϐ�}�!y�qO���� YH����:<'=��;5n�C�tNG�ZU�DܳF��GK�����}|mO%� �g�%�k�w0Reav߅T"����sQѮ�0w�9�p�㐣o5�rX��v{ק��i]F��2�%��O8��������B��f�o~�����Fn'G[�u�B�]m��w]�BN�zcM�VT�/|(7��Ivn���KB�^%��SmԶ���M�z/#��+feI$�����f!J믂����D��_�\���rV�ې% ��5h�]�W@bx�z���3�"�8��}��WU��X��L�B�w�e�.����r���f^�J�Tz��CGɑ���\�ڏ@��I�"�IR�C"�b:"[�ZtDP2bO_��d�?�q�GaW�U���F�ϵ�Rijm�r?%�z��lg�j���<��d�3A5�z	Z�'X'�w��P���8e�7��x!�Cd5���?׍��?2%��,�.S�K0��'�cF��Z������Y�%�wO��T��x�{,�&2� DzC���}������,�c����	r�l$N^�$�O_�J1�",�E��{ܝA3C�;�_��}�a�������A�Ve�o����Fǌg�l�j��cIS��zRM�h����Gd@�|������Ȭ����^��.h���L�~�D���ǩJP+��G���0���s��:�^���7�^��K���ܺ�-+|��W��}��*ޝP�"�
&g�.�|����8*�����-0	��=�����K�ɘ�,y�,׬�Y���r����#j�C�U1k���}m����b�3���tk�P8v�\����T3��_��ŪA'M��o<�]�*�`��.Y3�A���s������̘��qUWɕ׊�C��"�M3��\�D:T 1���]�/�1�c�Zg�]�&�̚�����+����)��G �Y�+����;����^�m�s[<O|]�j�6�h���r)�@���ӛ��>ڷ&���4�K�t���T+�]7�6�@�t<��h�ZG~A�d��,ڪ@�pTp�r5�o 
LF����%���J*<�+�>\�H��MuϷ��[��?��+;̓p�b�mh�;�AtU�m����!��q�mp�}]��η�j��갮�z^��{���[e����jI'��Z���	�T��_�t�~\��b���;�s'Ȫq�ъ��X�)�"ྉ�ו�4W| %cO.�E�o#a��E4����Ӭ�=�X�����4F��1R�s��CC\����U���������S?68���FN⊹����Nz��������Lt�'�b�~��<��[��jpg����3���O�诸�K�1X�0�o��y�g��Б�9�	d�Gyϒdp��;�o��f�s���M���0TGX��q��]މ�P֢��M�^i�����>��t̸E��v�
��#XU��"2�����Q��-���9�N���L���ܼ.�B�M���o�b5܆�~5i^y�����˕u/ҹ��U��/� 	�4��]��[�[Hk�ܛ�rm���^n0�n�/c�(^��U`�^~�&��c�T�����}����F4*xV�L����O���*�`���A�EI�&��F��0�O�v�.ri͸�{G��Y5����p���)]	&�GNE��a���6d�6�É�e�C��<����(���#��@3��_��,�IŠ�"��_h��!]�^6����G|�V��9��&y#��g���Jp�ɤ]&.�rOF�^R!n!qZٜ͟^�խ�5����c���h�3��ή[ ?Q��b������=��N�7ݜQ�����~����]�CX��ԁҵFc���VK��ZթJ�t[k��ˠ��w'�p��~g)�ZT���P��Ӝ�Vk_=���پ�3��5l�vR�Q�F�-P']����2�ɂK:�� ��B3�A�G��`Ǒ:[л3����-��D(�U�����qPn��� ٳ��d������Z?�l��B^�b:o,CT0邻sjL�Wz)��藪��<���j�%Q:��#���r��4�}؆L=��I��|h8U}B�61�0����s�cz�f�-T�h�k��h t)��iy�����E�����b/'����،���� �~�� - �lEA�����'��7��jX���c�v*��տ�w�C��u�����O���!���.}��Q�۩��_��H����v��Z{�_W7ɖ7�ef��9�N�bp��:�)SG�k����Z;npG)�����/����d�n�����;�	 I1W�)��5�
�� ��	���#�bXK��a�c��~���Խ1�8�~	�!�n�Ń,t0 �^�J��-F�E�����
z"�~� �[���1|b��]'>�D��!�$b��(1b`xGD{1>�w�u���o4s��W�L�ˌe���U� '���pM�$�z��у��V�[O(7�/E��@��
����0&�[D�&y�_JF�Gۿl"}�et�oX���Ho��E��p	iIt$"(�����'�˧3�Y�u'3��[��1�+��D�)>��4�;(q�D��˄�X���ËU�;�B�
å���Nu)�HT�E��4����Pu �L�G�b�GN��y3�(QSH�U~��e��J}ȱ��t�<8�dzp�K���!����2ˀ���s�0A~����ͻ~�v�PE�����t��Uݖ�dբ"�ՄR�>x�)nml��D��0�_�����0�P4�u_ez�ٜ1�غ1�u����,��S��"��~�����	f����l�7��
���ߧ��g�dW�Pg��(hr��~s�����5
�lI�:�A�D,q��{��h�>��P0�X`"��YO��w4}N�GH[7����#�pN�0l׺���A�6�Z�P)t�9J��>������~)p�J�6�M��b��T�a��n�@�nuV��L�٤����?�G��K��7ס�� �O�4�(|������Vƪ����>/��vk~9Y�Z(�[�r^�[�$�Aʪ�a��f��O�hiK�֪��-���J��(M_�E��o���l����>͋��3����},#7>f�����t�򲓣'ǩ�0�0U��	C!�5TD�5$DW._q�x�9��c���#�圡�&F���������+̆*�jz�� *NqIo|��Vk���Џ��w�o`��P�\�K�dݍ��~�K�zO�#��Y�S	��ь�ĭ�!zة�?j���Ҋ�y�����������i�$C��v�YMK�[,��f��]K�=���ﯮ�7�#o���	�r�.�- ��L���.*�$��B�<�Rk��f�=f�Ss�y�2]�A]^��\�g�"��#W�oϊR®�&��?Q��^��x�^�>��
��S�#d�LY a��I����w!k+1LaS�`6�Q��
Ȑ�c2�M�lT����g1�6�c�E�˾�e�Y��S�� �jga����H K�D 5��[4�1�v��%7��eP��S��[�����1���5v��Y�u���>&s[X����~���C���G��1-�FPJ@'�J�Irw���I����d0���W�.^�?�ոY]�A~�tcw^Y�~���s��X�B��oݺŝN�玀�r/�?R��uɭ쉧[-Vڎ�3��L:#��&�@��Q I3/Xߢ������3�f���|�)1��]o�Z^�|c�W��V����Шj�������V�w�}�#,��+����uG@��!X����M
��dRL��:��A���+�s�H��ඹР��"'���}Gn)�@��	�6Kz,���B�NR0���]��ԄrH6��c9qN�6�pO?8ڍ��V/��PԢ�4�0|�����Bw��%�b��8�n&�0. �������[���������ΰC���`+�\�#w7�O�+r�Ȱҕr[#8��,Π�����Dzif���t��v�����i�t𧁆�S7���r��<���ˋ
8�#d��D�=����Z�i�	`ΘV{��Pv������߈?�#?s	Y�O�o*�ZL{��%���^�v|M�5����p[|�q��D�q�}�� ��^�3lIf���F��ge		#�y��n���_�Hk<�Oeai��O��w��F�m�4�[�T�.�D05���G�%��U3��z1��	x8���6�'�1����p�	�y�v�M�i����w^���?!����S���t�Q��i�b�N�m�b�������G���޷$��l%��r#(�XeYA��˻Z��4.�Q��hġΧtY����ý�tm�s0�P�~�� جu� Y���m���_Q�U�Jw��{D����!��4@ŵ�@Ic��ZI�$��tW �f���U��Ɵ^�3]��q4CI߯��[)�$�W��q1�:���G�:YiC���T4 1�5^�G:�qŏ�Y��4g��u^�;�&�L��UzR��C�?�H)�]�;���c���9��'�j3t=q΍���LM�*���F?����������P~8%��7���IȢ����#�f�|{��������=~� �� 壐��Bc�&^����0�pT}
���u����7��{�Z�=lؘ�I	�&v&B]67v80�,�YR}XD(~m[���1h(%G }�/��Q�%B�#]��n?bbe�)|/ӣUi�յze^�� �.�uO�� ���{L�$�J�\���K��'hC���� ��=��)�!�U��%f-�?��� X����$|ҫ.�d�ַ�ZNWY�۪4<����U������;$�>��##ƌ��P`"�i�.R�DO�Q�v`��	4����˛L��-���{�آ :����r��4(��y�Z0��Y�ɿ:#
9^�Q��!��{�nʒ�͐:�^�� %ba3���7�4F�J8 J� Yf��=����ޘ˃A�^Ց�~��y���(��=�lF�G
�Ӆ{�	���Iz���fn�|�^�L�vp:�H�D�E2cKS�t�*>�o|&����u�i
�,A�s�+�.P�f��.yw��	�Յ*��#���m-��[3@��`8��@�b�N�d���/�PU8������i@�Q�&O�y
i���.���Sg��.b�wb�5y�� ������Ҷ��A��+X�e��0��9ou.�>��N��~�!���AR_�Uc�s��B��Ł�z��s��kě��3^i)T��n���Zyx"Np��Ӌ��`�nOQ������¥7C�����g9!��Ӗ��)�6!��A��a��D��0��J���#An��x��/��ձ��Ԕr�L������ �Yc��E����U���Mm�E�x��_ʸΫ����:M�U�M����_��~�F�����@��#0�rث,�L��/��v��Ӥ��[!H�H�dbZ�q
ȩ�L��{P�~F�oB2K��.3̽,J] o�h�[��;|�P� A@�uS�E�T��h��"�".%f Th�?����u'(�	3FGB��a.U��܈�����b�%K����<(z�G�c�5�
^,�d7��[�@�\ј	�'��X\�ƀU�g�e��1h����}"�8�Eף�gۓ��X��࿤�gR��WYYMQ�e�NQ�g��tC�C��9�['H�zO}_�Ӵ}�VY�M��4Y	҃��<Y>��.�kٷA.����E6���܊�|�K�f^�G`m��3��Z����� �
)���	lV�q�79H�w�\I�s��+L�ٽ�}>]��{8wj)�F5�ړ�-p�L#:�d�0g��?,�]�A7�_�0HE�3����C�	X���;�!ˑ�`�L���,�im
��.��O��4M�Fx{�oM�˜[���y�Y�b$[���n>�Nߚ�����7���Pꐗ�f�1R�����7=3@��@\��P5<�6�.DZ��g~ݑ'�k��lɢώ�,9��o*��+pO�}/:h�h�XD}{�5{�)���P��K��#���I�l�r�b�<�X�������W^G�s��
(*�۫ځ5���BٞѤ
���s�`(:O���0����E;����5�7���l���?h�A�Pxde�G��2w�1v��c ��Mx�)E�4�a��nQ݂d��q�y���f���y��:VG�"+���Q��pK�v�f�4=mi�",�@O��H�l*m�we+`�a�:�$F&;���%۽����"vq�,�Rk�2�N	�z�
����<}�DPc����ZR��V� GW�Z�Y�-�03���Q=e�_���jR�����	��>�f'|���Vϖ!��8��Ԋ�ł��p<��K5�Y�[�l�!��#�(�$�Š�Y���m�;>w+x ���O"��7�$`����Q���,r��F:uL�f�{y�@�{ipB�˲r[�Bk����Іn��oX�6L��ٽ�I\�:	u4?���O�eIO�&��q���6�'�?�h�*�DFy�Z"�1���Ռ8��7�(�2���I��u��G�	�$S=��@�l�@S�l��`r#��G'!-��������F~ �P:�Vv ".
�/Xt]i�0灣����O(��0�IJ����AGv+������F����� ��b�nX�E���W>�C��Sc�nç��]�f����R��h�m]�����]���j��|��Z��ľ~�Q/j?z��TLx�<7s� |4�֏��:S4�������auˑn���D�2}PhE²�{ WQ��s(	��3 >=�fb�4E|�DXϐ�[j��÷�su��Uc�Fb8��c�*Q��X��q������#���x��G-���Kױ���7��n�u+��$�� ���Y�z��-�h#�O� 
��~��L�gP���U����5�� ��dY������ �l;GI�$��{"^��7*߄B�+�=�D(����]�����	,3;�\��T�@XV���f�!��d��8��*����4)}_5ޫ�/=|#��=�0���y*���X�;4��%��R$a f�*���v]�$�Zv�\�l��gVY����ʄFa��&$���*�~"��,��Ux.�r��O#b��:�˔N�))@U��'q�h�J�m�
�m�J�n�ǍF�w,�n�	%�f��&%Һ�f��9'_�xɻ�����Xt%�+,kx�f����hClr����nN�&��WS���`1��~Z�A}]�iE������OĿs7�9d��m�C����v�,���ǀ�����tsZ<�VX��1*��y��K��A��H��D�޾��=��R��1^!Z�%�j�a(W���|���;A)B���K��V��>�5��V�+�TW�H��.��g6E�8�FGa�`��������.D�^�*����øL���5E�u �QxZN�_����DWg�Z�z����͸�0J1�V��'l
p���q�ڂ_��"�9�y��k��cQ�Av�����j�N'~")7_��puf�a�!О-%���1 �k�cj*��A�&��F#��Os���3˳�1��6�~���N)�2�݃���������;���S|�=L{�q5��R�ߏ7����d��uS"���d<��ա�J�o/f�T��y��Ư̊���_��i�d����BqQ��\�H3O�3U�d�m�ϔ�-���	�K�,�T��*��L��d��|�p��*����k(����fTW~)����<k�P6���
i*go�}gj���SY�r��g��M�
>��(�Q�l�y-�uvw�k§e��D
��TR�=,��[�~�3��x9�j�����S�������L�ZΨ;�,:]�au~�K��(�"(,��W^�*]|�Z7
�_� ��s� ��]5�C��W��J�.�� ���N�\����h=��Mh�/ǝ�{��қ-(#G������Sk��Fĉ��I��sr����貚F(�+���)zC8�c�-_��펄ô�&L�/G�uӨ2�!�`���ir�{�}�Hq��b��
~j㴩W�n����9�s��&��F��汲�$�4��-�Ne��Ҕ�z��D�)t��
��T�3���YN���s���_��7 �陴��8i�a$���KˀUU�Am3��% ('��1{��(��_"��%L	��y�W���
��c*�K�Ջ\i��T��)�	e��l}������i<�i.	�8�Iu�_*,��wJLTrJ���4[��MM��9U�r}�d@*
�q���0Z�-z�E?���V_Jl�Bi����/����q�{G�8�c��3 Tqh;�����64�I#:�����,���J:�\[�)�����!�S-,�W���az��Uf5�	�uHĿ��"��ӡʟ)���ŗ�Oei�O��9uf*����'Yn�ԶB6�U��w+��*3c\8�;<&����d���|My�N��eu��	�����}PxE;a�l�1���Yh�3y�����o� �̰�8/V�a/��j�v�:���m�W�u�F%Cq$��n��A�x���Ҵѝ2`� }�~�M~{#��cj��x Y��ɂ�U�����-W�,���Hȝ�xM/"��K��|�ߍǾ���*1��$EM�6Fza����z��4Z�	V5c��Eoes?�jn�hĢ}Pd�ۼ���*�ԡ��������$�<+Fl�ǖ$����!��>1�����5>���0<EH��z
��f��m�O��X� ��`��5���!i��ut�P�pk���h(	�����~���Q�G��v}).�3��yO���h ���mj{��Pr�7����Fg��Of"�_tN٧��[2������-0t_��G�֢�CѵLj�������=�.��4�5����a� ������!���m�^i�rli���z?N�`v ϟ����w:����ݜ�28WV-��P0��&��Ѷ�]���\�R�ia�p!n����0WIY���H|V������n�>��!�o�ZAoY���K)lTqh@-��9{y�>���6����3 0�N�85"Ca+u�\l�E�5g�LZ��*o�_��Is8n��l��5֋�q1��i��Y��>RX���8O�-��Q�<�L���������@�j���CD�V�>x�|�_�˲�Mm��դs;�{��Ř~�#�8�.�� +#��~4}U�Ħ:�m7�WP�#1,k�mpu���H�����.����gtE�6�1LR��2��� �P��v��֗9{2	_���lH9����!g���n�ʡ��?��7�]�<���R6Cǵ �Ʀ���lQ����怂���j[-mO�&�!L�w�،n�҃�K�p�:�!)�a�#�m��7.'e&��EX=yr�P����.�����o՞�tD9�'簣����'>yz��V�e�h��6M;��Mֹ=Y�fНa+}ϩOxs_�}X�+ObYd&G֦R�������L�y��*��8H���s�jM�$aHeK��H�,�i���x���
_���D?�樷3�Iݼ2�h;��[Q��A�Hz	�6��#�fQV��ڡ;0<��h��m��rDP�0 �	s��LRr�-߬�j�p��պ_ӻ�4}4M!�sM�jxi�<���U}�����ƳZ=�j�uc&�56E��=?Wk<3�H˷r��k4E��'\�*ݠA�U���c��6������Q�ؑG��m���ѹ6UP�'�  �51�0�kϨ��T���	Q]���i@����Ih{�iʌ�{�)LI�m�U	S)�ǡ.�B$�g�ƫ �d�6�sQ�oHD`ʨWw����F�����h��Z�R��6͘���$P⓺�b��M{��w���6q������΢��2�-	X	��鞐a��-��f��ձ��巴�(�����#U���c��t�-����0�	�-\	R�~����z�Y-<[���!1�B�Xai�&.t ��#��u���O�>�O�?ISwe�4�� _��9L�0���"��m���u�5M!��m��U��0��7i	��)@�> �:6����0I����XS"I=#��*	�İ��ŋ�N�,?�B�1_Uq%�����N�����Y�[un�î��\5Q� f�ƹ�:���AY��+x��������L�hC�*&���8g���j�5�� �k[�Y{��ub��������'��I��f��+|K{д"�B��md�+`B�)F���j�����d񔓇 �q��gղ�>��&�a�P�[�C�����R)��;�)�Ͻo2yB��x���W���7'�4�{�K�ʚ$�(��S���h�::`�'���Э�i12���sU �*�[Xs��J��?@�t�]2"���.
n&�Ȫ;``�� a�Fd�v�Z�eEǵ���L� ��l?�;�'i�#�hX�D��f�rH ��@�CIJk�{Q�P>��	U<��aK#i�N�#��/�][K����6���}<�ĉ��z�z^�ʹ�O���ҏ(�Y�� �W��x��8��АFE�L�:bnS��>�B�9>5�kB����vT(�m�்��T�Z�Ϥ���U�T:��v�F�y<O�ʎ�$5#O@�j����w���l�3�La[�'�φbI�[���г#�h��wm�,���O,�ђܩ���ѕ��E[(a��=Oǧ<!�$�	T�h���y�=�/���u�Uq�3�2�l
8]��hǂ׵K�YHK�*m`4���Нν���5�v�J}X;�t��~jc>ŝ���a�3gO�W��3�r��3�t|Y��n�)����3t9���L�3Ͽ:�-���דt)[�E7�<�9�_�d�ݥ?_�|����yƗ*��LP�M��Qӑ���2��L�����R͎DU�������C1�#3UjeW����o��RpT�!� �hu�Ѡ2#y	2��I��&1�Kh}3�׈@Ǚ��o��L�e_/� ͟i��71�7�SH�tdρ��gJ����s�?	�H)é����1��|�K���Tkǽ���ۀ���
�! %����x۷���e ���Ie���S�*��x�_@"�aH+���O�����,���K�d~f䱙�;��)����s�����a���m[���<���=E�`r����J��O��5%l(�j:�h�M^�_�* ��p��t�kH��bКK����@!���W��PJ�K�X>
j͏C	���nC!��3`QkH0�a�����~���hԀUA"O�P��D��.�4��� �YCd�.���G��#�N�ߢ��<�&P�p�Ѥ@噳oD�
�6q��S)v/y�H\�u�ǱhCC7����o�|}ء��E�Į���(`R����(n�8�#����:hJ����,��7Te��Z6���Ĝ����#���P����VyԈ�q.��i��xb��'%�}�=����+�_�s���p�؟���b�����~x���r4�wSt�QUꝈ�'��Pgl|dqɈ�W�w{0Y��E)�VF�rRӆ�]�)k��ZA�u`>��]!d(��B۔�ͣ��T쬩�'#�q�0%.�:�(�ߑ�h�ޏ#�ҿ�C&�{ΐ���c��^�GG;�����V؋�F�;�)��<�7c@�}7�Π�-�
q�a�;ʯS���kG]��xj&��
��%Zv�p��h)�6�y}�/͘�į�л{����'ƚ�s���`��J�5Ýh���������kr:%��/�|��?�3؉�ŕ��u�ה6��j�h^h!tPkZ[ܸn|鹞0��lUp�����d�T�����8���� �v�����;�d*(G����j��z������2�f�ը��h��n'��r�<vh��}:q��F���ժn;�B|Xw�fv����5p>��a䕟z�`��̡�Pj�9��:#lC)����8���V�K��_��,ǐ�m�K�?��C��6�T���$�A`��=/gWd���?���Og�+lQȮ ���P��{�{�ab6}r�2�m($��{@TZ��"���A,��׈Tس�ٜT#Ov���Y9R��:9$\���%ܲ�	�P����{K�-3�D���h�?��,10��y�������wx��-�Z_�1!��/��+��li����|�3�څB�Y��[��Xʪ▹��ߵ�5����',NF�����^o"��j�����Qk
S2a�}/Tۑ�3	:�O��,C6�a+��ɑcZi*��UN���e������4�<CJ&�����,t?�2��:,�ܴ�Y|�-�����ϔ<��fܓ!�����k�Vq�@�������<��_'����on:6��^����c*�$�:�j�9�!�*��X��Z�p_n����Ś�z�.�qL�pi=oz���V{ޕ��=�u���%�ip���ni�	{i�Z6Q}]�X�[��	b��3ꀶ���e�ӥ�jk�8#lstZy(��Jsv�W������*���v���()rE_2�/y[nn�㨏:vc;-ߞ�̧W"�;�%��7%�]�
G�Gu�(�}���T�m����c��}��^3���`�L�l��%ް1aâ4?�_�H��h�u+�����8R��!�<3Bg��U^!�/�d�נ�%6Iv:jZz������`����}N3X�1�OX0j����R�Dݵ�;�x'[����;�)�^7|�|4�(B�FD�9�l�A��M���#�����"�+�Ɉ5\Qu��!e�q�a2�BQ!���(qA��Ca���.�
�X�Xz���_�1>�Ia�����Ϙ�N�)A�3�[� I|�������|v�� :MO��c��ȍ���g����]R�?���o��1]2�4����h��}�ɕ��T�����;7�`s臃Q����:�N��xwM*�V�+M�O��Jo��� u.���
;�n�A�ۅ�nz�J\&�f3h���L�(3jz�ww��[v���pW�(3`��c��B:	s�R��P��c�}���&�k0�Ff�Ŝ�o���g�5NkG����]CE��������sۥ�7�� ������w��?�Rf�C�P!
�^����Z��E7f�\��dD�Ie�f݇ـ���ԞqM���!ڪ���a��zP[>���v�����o����q�M�R����-������3PQ�8�-> ��Å{
���hٿ9��P��/�C�Џ�&܏C��4�J�)6�s�1�h�ɩ�VT�d��(%�v^ýrL���!
[�5��>�����sL��Y%q�:��\D�`<��OS*�rH=.Jc��&����6��	�o��^ʁ��������ۊ�+�� ��/',����y�Jsgs�u�MN-���v�v#�3��c|���OS@3���j���f�3���
��p'��ܱ>#��
1�����߼���ܹ����sq�g�
��$@hUSFsWF��W��a��NJк�q��	}�Et�c�j�.�e�p�[��P6*1��J�h2��𭢵�g��sP�
$r�jH25���	�?3���O�#�=��*���{�	'h�,�ob��7�n-.,�?��0%��o����v*���T�|}؃� � �;rBH�HnJi�iF�K�R�(���~ i�j2]�q��m�6!�$�"�c����g��<Î(O���n�L��D>�լ�}����\��,�s"���� �-�<�oҁ����y�#מ�R�u;(02�l?ɞM��?�Npn��2g��(t��=U����v%!2y#/#����d^�����7�!���'���~��Mv%Kџ�x�> �}�!����
�bQ���y<���媲�֐(&�b<�*���%�K�jU�-��~(�h���4�8���_L�K����M�p���8^�vA#&~�xH �m���$P?D]L	o#�6#��Oy"�f�GV@UAM'�T��Mb�ƹ�XX?DK ���pGJׇ�EE+���N�����=��X��g'���,���c���<�o��Hf�.�-B�5����x���6e,�<=��4�}�1�=��┨�G-h��@�V�?�/�����N2���SW<B�Q�e��:ڹnߊ�l���{l�	P׶�>@��E���ȃ���L��P�kr��ėx��B�V�S��f��J'�fe��Q<� [i�g	E����2/�&\|�!:�>��2o���}b���V��I�[˰�n'��Qt/q��T�f�۲���+)��î.��L҅|^rc 0�1�
w�_�N?t�E��MB��ֽv0v{}��灄�N3���	��Կx��'��5�i�O~ɲ���|�	����r���(�2�iQ�\�FǬ�� F��_ES��]�����tq�R�����5yj~F�*z�A����GWP7$5'o��¥8��<3 {�,�fZ_�v���O��9%�:(ٔn����z���X��΄c;dT
ߝ�X������u��gTH� ���	Յvv�S�nYv���H��o�z�U3���i�5�҉��7W�[+:����$A[�vǵ�'Et]���T����{R����E���Ko&r�Ϭ���&�p? �v��21��|J�i�g͞����F:.V_�����ABGQ��ol�a�*��'briQ��T%ٳy�7#F��؄���υ�ӱ��"୓$�;3�ż��7# �� L�_���d���S����XC\.x*}�&U��� ���)��Ҹ17�Et���ѽ�a��ݣZ+0D���<����T�?N���xK2q�s����ȴ~�gςm1n�������� �����1��eO�By��B��W�գ ��s�X�\Ղ~�k@�Ґ�SJ�~�gv>SJ�Q9�,O�_`��J�_���<���r!�.l>���F����g�l�l,�h���h)֠�
��&���W1�-&��=T�� B��]"�9�$s���&�"tuj�eD�a��H��BF�(�nM�s�6�3͑R��.��ܹ��կuаJ�̪�#Y���y��߿7$��Uy48&����6،����z:|W���9!�9�(���e��fAr�-�bhf�Ih�C�i�
3m�@��߬��a8p`wF,�]�5=�"���8�G�sn�2�Q�.mG�,���?8�c]�iチ�Ɲd����6`ӮW6}����(
��ƯOR� ��������D�]�0�@�G�@�6L��͌��R���ȎG����؃����W��" ���7��W��RB�:M�����"[�V��������h��@ D9+Qp�*e�s�# �S�/�W�A(�:�]��6����	���	���NyLZ�ڔ�u0��F�B&9��N�?��p��*�����'��ղ��f�k�/�Mm";b>���|��=����ج�,��J���Z�XY=��t��A<X��G�� ;�8��qj�윑�lEi���'*�d	���1,�������09��`jc��	N`�*!68Üm)�tu(��"f��i��e( ���H�p�zq����E����8�.ҙ~m�8$��T/#��ڈ��=s�U���q����S'�L��B9��؍D`|��ʰG�w��~׳����>�F�2�WC�lW�RGG�bҜ�E�dppq16�
�b��-�7��؋mY���M�'Q���jbV�Gt(;��X8���q��Z5x!�ߙp�?IPb�e�ԛ\_�.ե/s'���h���'�\}����Q���9��w����}L�"%��і&��>ԯ��l�����QA��j�c
w��&l�ʔ҉�Q,��W��pN3����G�^����A���ĸ�'�_ol!�۽��ZX��zRt�X1�h�z��q�F���p6�ʎɓF�~$ی]T�`1pr7��Ǜ�c��&w�������s�9��&��Ex���ks��%���u�҈ȱ'�_�d��pCL2$�N�s��'��F�,�/��l|(�HҢ8q�2�0���M������]r���da�����=Ǜ��6n',��,�dE9?��UI���X��x��"\��H���-O�-T������v��n]���ʵ�O�~ow&ж�����y���`%�L���1��S�����$x87���4���%|�m)u �IR�e��u�H�
�@n���Y�Wy+/䁰ڃ��V�B���օ!�ƌ��A�W;ˉ ݕ�k��aw�&�D�+'�'֕�[
��f�KPe$*g�\��Y%I�+7�j��K��"���}�NB6琱���I� ��0��S�(sXf�B� ��`����n�Y�p�r�RX�M�Ꞥ�Ҵ�RK��:)Sz�"�$���$o�h�=.�����9�d+N�"��:P��`Q9�Ky�b�����hL}��^���P�-|��"Ж��{/k�:f���QҞ�3��ؖ��p<m������Bz
���[��m�2�y]w@=��;7���p'3\
x��A�#I~�x���m�_�q�]Ib�爛��\p��7�"����������Y/ˊj���5	���(��o1DS��ͺ=c����e�-�A\�����f:��:�� ��,������-{tI��4	���{��,4KI&��1k)���͍Z�PT��H� p� ;���[fi.k��<��&"6��J���EE��(L���/^�t��;eU3��"�ai��5�G�\s��F��A�.w^���"C��BF�a��]QG�Fk�Z}�<?�W��m�҉�xJ�x,���+�p����gʖP�<"�n�"&ڟ_(BM�M���*��3�:+q �p 7�Q�Q�K�?*�n8kVM�G$��e�@���?�.B
)�\7}�^BK�B�[r����
��4����k�L�.B^��"щ �/0��^Э�ow������$���u] UZuМMHO�WGv6�%EKx8�Z8���ej;���f���qݯs�|��g֕�eV�m��<PI2wƕy�a�h �R��ZO����+�v�����W� �0v~[��̔K����r�xg�M���k6������D#���
���G l���Y�o�ڷrA�LO3ҵS;�H�et�P+:��4{/vh/E���(�HH1�/ܩ��П��.VB]n8��=uɋq���2�v�zUݭ���V�xv˛�^�<>P�b�~�0=!O�Fa�������<x��8��J���&B]0ΓG�o�۟�=�,%�V� T�{-N�S_A\~;�2�wэ�pT:\v1�LLY��מJ?�o�Z&�(��r��}�L�$��%*���1�n�>�2�^��a��.j��$��f�1�N6GD�ӆJ�Qh	ը��%R�_����2�p*��هB�5B?Ҍ��@zT�
=�x9W�o��-r�Y�@�Y��Z�H�x߂m�kq�l@�*r���Ȼ.`WB�B��� ,���}"��=����}v{��Gɛ�4��3�U��"b\����� +9��8�%��L�:$i���5���'R��4�W�o ��q�0��. ��4�Z:ъ�SM�}j�,�1��K�E^G��6�S���0�I����k@�Y�4�T��k�f�����?�4j�Z��p�_U=�ެLD�EB|����k�&k�VҊ�:�1f�6fr��=���S��In�Cbz��*�q��2*ڬ��y\���]b�p&+AmEs�����i#�&@U��"��ǜ�V����Ti��#B��r8>e�d8=�[�%�CM��AT��ܒ�b ���s��~I�j'���( R0�U{}*(I�+t
�7i�g��lwL�J�h9=fO��ի-��:ډNY����fDq{��Bd_B��#
T4Z��:�������9\R���l��MV�I��ۇC!3ݼFq�����ֶ�AZ��n,v�&�'+����o\	��Lf��X������R�=����{��gn��E	-��K�yb��%�E��}�D}�D�݊�-�d�\5��};ש��sșӲ��p3�۔N�t����A2�O�@j?���T��sSARYΚ�D'Yʖ�6'�i���W:�����[���4�+A�j�hX`�� |}x�7@2jMn���� Q+ǣ���
�ؖ��R������u�B��=����3��,���j:��>.�uG�n�f�[�xVI�����I
Ӊ�C��h����m�(q��"TF�J"��3�wC���"d0�Bx{�������;ϱ݅���Y���!zRC{�?� g���_�G�ӓ�U�}�T3ӵ75D��g6�V��������3��U3~��O�,��l��+tʸb�b��k������k��5��Z����Kc���ˠ,����e�#D�`�5��
�/ЈYK�-u��3��(�0}E�_Su�EL��ipG�*�HVY�C|;��s�Ň)�w����������S��?>Ƒ<ih�o䐨4�1���U��q�0������wI!�'� ��l�1U�:�ؾ>�K�2�H;�A�]Re�+QnD	�m]@q������w�aU'�4F��s#�~������B;�\�/U�xrAqd�x�=��Ed��
r����Uԋ�"7Np�(�&_�	t��BQ����<�P{'����|%�Z��o�t4X��U�<�?"��J#��<P."JŒ��,(k���-hG?�-�G��S	\�|��챐�]�C�: �i�G�� UKq��쓵�]��g\���U:�<һ:/=�?_�}BUh����Yo̳O�댱T�������s�����t6 �P�UK��a����R�G��=�p��`d
�F�Vrs��С23w���A���1��ݚ�����R/�0��j(���Ӧ��r6�G��/Q�Ȳ*���Sh*��C�ޅ»5�A��'�%��?�I�QQ7z-Per7�fn�8u �$C�|:��Z�pWŬ�A(sn9�8zweګ��ׂ�'�~�vT�����|��`%�?ά$B���P^�5#�9Rd��M�ĉ<���.e]8I]L+�!w�Pkȼ�����I� $o��r���/���@��6c�(�l���Ĝ�b�9\O���L�vK�!Č�:Z	(��kf� w���?�9S��a�K��)4�� ´G̿ߩ������J�ϲ2�8�d���W��������h!�g?@��I�g��fE�Mt%N	�e��y>�Z-���(�W���4'�|8�LI�,M�߻�Ʈ4ŝ/�="ql��U��G�8	~��dۥ*m�vM���s�����KYc��Ef:N��F=��5�R@���nբ(�+���⾴��l8�N�{r��9i\��X�3��ޙ�]��_���0Ҭ'9�
�gS�~��l�g{Q�9)�@E��TM�O��-�}�k��n��FJYN��!��/��*"�|����^�S�v�EZ>�L �g+��������Z�H�3#�
@���;4��	�,���q���������I��>�Q���y�P��N�9�.�G!�Er�$o_�3�S����u���O�6��/]P�S�MdR���d��su)y��ν��0��%R�� M�ӟ�F6�ڢ�n.�u�S�9<3쿋��y�C��5�*�jK�$����l�����#B��cu�3(�W;��\���i�3� SO�Q?
�ү�dMb���ѧ��|X�杻1R�F wp�raA�let�E�i��q�ʁ�C�i��q���F�YD�2�:2c�"N~s�Ϊ\Xv�K������|�;�!X����4���2 �s��sm�ƹ˻d��9Ϛ[\�^������p��(p�����}޿ ��Z�>u�C����bDA�W�6�C5Qel�݃����?馩^;��>�ި�,��Q���
$O��p�{�c��^n��j�~�b�RY-�DGz㤷t�CO+��:W����V�>�$N�py��㷲�(#X#�h��+�~�~bQ�JB���!E�;Ӛ�R�@f���Sw\Al�%����w�>�\�
�5_����0�4 �v25�م2��(��čY;���)2L��vo�`&�^v�\,�7�m*��aQ�(��V���Mm���Ҋ%�1�?IV�a	��|j�M�FW�
��>��S)�v�6�A	8�f�m���n��VG�L����9�!|�ܡ:���n/{��wRpʃ��D֜^R��(Vt�A��?\1m�"�-7��YB7��ˮ��V�\"K��3|�~�]^ioʧ��7��&�*k#�<W�w���-~�����!�̚�>C����:J�%O7^&rN2́׷�;�����UС�[��$�7 ������eX���(s`�&0�Miz���f�� h)��8'��H��{@��8�NK{�{���\��M-�dtT9P1�#��&5�����ӻ�����S����2�����!�����7����O��ډ$���"#���7l����oSsz`!y
~��k��kF�5`��,��=�o51�uLօ��R�G;a|K��,��o��ͮ=������6�K�o! ��_A/c��aSΛ�1���k�a���v�D��G;�P�1.{-�n8�}���i���Z��!�y�=���V�Қ�����9�d�7[l��$,s�����C;5s���9�/�C^����Z��LR�$ڙ@U"����g�`�n�?
P�N۔�^n�U��&��Y�\��?�2z'"�+�b�9eHC�9�X�0��r��B	X�B6�����"���)�ç����$	Q�Tp>��1�=�h���8*.,Ƙz�j��T]A�.x&c�ݲ^�b?��x����|)����]%�	�@�o�7~���K��ʟ��fzyE�uz������bb��I�xfh[�П��tT��gcYȹ:�䦅�צ��e��hR:�taR�ë흴0��e7\���'�pZ�[T�����t�I�M\�,�#J�c���Ȝ҅�¯�&(�7��'����:�_(B��ȓ���]�&7��l��D�?b�;�k/!t/K"W�s��x��/���7�A����UZ?W���(;�Z�5�S��Z��L��Cn����E����B@D�s���6db��}f���c����!3{GyD�?�CN�z���eS�7퉆g���߀�M�v�$�7 �#N'��.n���M+�X�V8I��3~�K��M�x���J���{�w-�P4S�A,>��B�n���5����K��0㓛,'6�uD��ϭ��,~��_&ҧ��u.)�y���Uc��o��Ħ�NyL�i��2a�J-���m.���~�ԩ������&��其���G�꣩v%�t�~�O6���O
�
J�u�Qm�@����*=�]�I�5����� l�,�.SZ-�b^���9����=J��{*$��f[�&��"��$\'�M��ey$�@�=r�q��?~�-�FM)+P���8��DE���ټY��@K4G�l�(Qr���I�
��I_�V��yX��B��V�R�q�P �[�A77Tc�I��	�w�-���$�
������|�[z�ε��r�3)8��b,H��7d��0i��3|A��~]��?�mMZlwjh���1մ	����^iϏ=�����+�	�\�����?Y��a&�A�?Cjꗕ���.{�熯�kfC����a��ܠ�u>�����0�J�vL��w/dF����r�5��LCdx��������4_�7P^Q����q5e	^���"K�|���|Ҫ���N���7��,�-�PL'U+:��%sd��Kd��n��݇�n~�6����f|����}c�4��]&�Z��;���.z��]~�.��Ss����N3�>	��s5���Z��J�E_�����������|��) Fy�������g�/F2ާ.X�5�
���w��P�/�$lbHq���a�L����"&����#���Y�>0Gh~�v�NHOw�����D�{~���-��*��Q3�f�F./�XQ���,S�x�[<��7�Q�w�Ҫ^�%���f_ֶ��h���Jcڴ1�ﮜ1_ "N̮2b��A�3m�o\<a�ě�[�;���%��ͷ�C��H�1M 4]��P	�@�� a�x.��'?����h�����p(�0
�����]0&�lǄFr�F�����%m��V�&��TF��%;>���"�>P��p9�`H�k��g���� ��Ȝ�n+���'�P�)	�D�
!�؊�Ȱ�9K�X�^y��ۋ�co��������΁�T���'��tDu����a39�m�
ѥ�������RÍ a$,2ГiC�0/���^�E4��^X���)l78-�V#Y�����u�9�0��*4u���4��k��d����LK �45LtT�5�Fb{o��\��x��� �P�v��o!ɗ �M;?���IQ
q���Tj4�H�OȮ����a��\5�	�ic����/�[�ϥ�".�Y�ޞj��Q�(j�g�#�Yq�̬�2�p5�&��Q���G�@޷���q��$�e�t���f�*�e�8����c�<�|����aG�pA��1l'|h�E`/���`{}�f��D���<�T�&��N���. �sD���o���}���9�U^7�.+�zd��t^�(r�H� �\�'	�����+)��֐��혻����-u�6aq�a��!O�J���p����a���(�nm�p:$�X+N�#:�9P���D��#��}����Ǜ���7%���&�̸�7��]�Ec�1��7��YvqvQFN$�Ώ��<Hc� �r�<TXk�����Y��G�/�0q)��(� � B�LV)�a��-S�]@�~�7*�{y:i������:�d�C���ʵ��@
����	"����*IxI��	FA���^�?χM0���c'��ϑ���4���H���x}%<[���n�G}n>�հY�B�:��d/5��!�zX4غ5 ���tL�N�?IT��1��;Z�)�&�Ą��,��Kz�H5�*"I#iy�N�h�5��i_���,�G�!4?�U�[��/V�q����:��:��{��8�\搝^%�
�t!�b��S^�3�.�<W���D7Hc)7��ZI�?]�t���e]�B����a-!�:?(���d�.�껧G�锵R��H�x��
k�/�^���[��?hN^U�t������ �\~�A�̶CQ[,��b���lS:D Dy]��w�^c7�u��~����/��@UmRC�Y�ru�j��clb��ЈN�r ��M�A_`���֣VM�����O@
�����j#��k/%�\��A&A��x^�e�fQU�J��&j0>X����D*�?٥�A�n�-�n��˿F��(�	?EH�Y}��&wE�UÀkI��f~ZQ�b��_ {()�"����P5=>[���B�J��Ni�ت������%���
���o	t^��oyc��>�^�_�\pqZR0���-?��0�"�N�6�_M@W[���[��6���_�,}�-
�B��%F�=�G��ZɣK���z�!r(?������~)��Q\V�>(�����jO~4C�s�S�4�u��ʋq.p_�9�^��l8Pq��Lqɀ����a�Ӱ�כ�ʟoP$<���u�))
e��m�~�,���w�$w�ߒ�\ǆ�(3��j�p4�$ԊAC���E$8���R�KȵE�Q�q)��x9�DYf���#0�fAl'�'�Y@���q��mj^r�Ϳ���A��y���1�����]���*j�D��L��<�F�ks�.�b�H��e��ً#p
*���=/iD�'+V�Z,^�2E�%)��G%)������s�T�����b*��ѯe��)q1G���ܓ��l�,�?�)1ce��0������޶X�+U�! �LR�έ���Z��e�3��q*1��6*bߜt�zR�����pٞ.��kl={�!�o�ώ�$ԁ��f��{�IՄ�,�m���e��̛��+���k�2�&�9L���
��+��sN/b�9G���>~-��f*!�1���Zni��@[iQ5
S��NK�i'n!ϸY�QX��E�?��N2`���r�KNZ\R��x���-0��8a8^Ua0|=K����a�7TV�����o��&�G��ԣ��y���!v%��N�[.r�(�N�`�b],EP�'H��>M*��1ۛw��5E�������=���O%br��>w�ʭ/�qZ��)��oe4�K�]�SoO�+c��o��d;,^�r3����-E7�����V��J&(�,����'��o�*Wp�.|;v��.�F9�A�,�Jm����&���C�w�\]7�d=J[��.�S����VX��Sĉ����C�^�{�xo�a*�얄��E}�^ݰ��U�3��6��w��5�\'j�(���;0�&�gO���S��x@E�A7Z��2`��H���	:*�8��פ0Z8	+.�fo��X!�N�Kx����N��I3��Up��<�~��[/~��?)�}�D	Pu�V&ZD�G����42��T�����w�}ŋ��>�]�*��E��=����]�j��g�nwY2�z�+o���`�!2��o��<��o�"��4vg�Uړ���ɐ��C�f�k��^IbMwF]y��;$:���fB�lY�ISuns��u��R�[��-V��s���Ϥ�d�ӭ�(2�'�K�FQ�X�T�)�+n� Z0~�p��z8꧋=ޱ�=��P����H,K�ͮC���0�DҴ�2��Y���W��f�!ѵV7�2�Ђi,�
S���L�-$�xG;��#�Lb�p|�A��i~Y]l�H��MpM��Ttd$���1�����]{���5hv��$���a���w����U%R��}#����[q���V��G�A-P3��n4�PtP���c!,6��$<���<�E�O���,8�� GDU�#S "��v��bg�hZB�um����.���^iQov��%�~�T��w�x8�8C��M�C2?�R�3K�� I&~���h/A����C�_h`kj�f����� z�r���@	�گ� �L�g$CU�@��քj���<�O�Z��,1��r���-(Pc�ծR��|�4�0�k��j�k���ǖ����ͮ��p��X@�0J���F�O�k�,�J���;���iQ�b"؁)	������d��Aԟr�EX�`I�����xkv��oU�%���N��W��D��1)�1�6����F���)��V��1^���3�	�%;��$bSR�Zs��� ��2��s�Gծ��jea@[
��$^�~��h �k�ei�����fdَD|��8�EX�|5���?)W��T��K�;���p]�69��L��۱&�������E7�a�H����^���W4�IX�>2��(����;t�����a �~u�g��JL�5�}ZԱ	����2�<7�������n�@"nQ� \�� >�!��1�3��cUh�Y������,�$%��X��W0�A���~�l���������QrsDN=���@}�]���/�~<�.=�W�{�`O3ȩ������y�(u�����Ta!<&ak����<縻<�$O��)� �Ǆ9��"�u�4M��B�T�i�1�%#KL�ށ�
"�!��X�ȁ�{�x����G��t�ؙ�-y�/��@R/���3�3Pӣrc#��p1�!`�US�+�d����RX���qP�1���O�^2*[`/N6����؃����"冈��MrD�Q�\6�2	'�[dDv�$mV����A�¼�;�!;N$)�(�,v���7������Ӕ>����(u���f,yXB8�z�~�k8�a��q.|��F�g)\��Hὧ�dE��V�V�tL�5+"Q4z��\���N˚LT�=�ٗ��=�#Zb�H���=�$�L��/H�����r(������w�@Tj�Ӑw���1��H���1@*=e�������WS&�R�"�;b�ѱU5�I:ЇL��G���W���6�X��M
1a&pQ�G��S�v�����n��%���m�f�
s���{�X1�����M��i��#�ho��F��[1��nI2d�tP�K63��X8Pp�Y�U��t�0�Q�k`Ӿ�Yiࣕ��%V=bD8�ɫ�_$D���v���t)
*�e+�����ų@݋#F^����d�e}��va�;e7�D8������{�_��][�eO��nRsQ6GDr�;;�\��f��|;=�����{�qŖ���*����?F�1�KD����l��؄s��7�Y(��u�q�79L��lw��ki#l�2��	����6�k+�.W{�ҥˠ����训����:,�PV�]BO����c#�ݟ>!��� O��N1o����:n4�����cZQ+`�w���PNlJ�"��,���~�v`�5��"���
���<$�)_)X���Y�׆�iټ��Sk�0���e;�����d��`����iO�҆_\_h4�s^�U�s�B>�.	(�T61I��n�P����t�!h bJ[z����[T�"�(��9QH�'hH�\*��xo�`��"3��ܦ*<=pۖ����HG�'��ĒTJ���@�p�t�I�@�C(��z ��q�1��!أ���:*�+ ˝Ф�-ayrwT��o��:��H��-}ޠJ�M����CqϾLR����a�c8������a��
���mm~!855$Z
���N/�S�8 �!�h6�!d��S��]&^`,�KS�O��<��tQ��O���s��S$��[&o�4/޹{	�E>h0(ϐ�I��I�2��YR�O���Ve�n� \Q�GWFX�,�R��ʫE ɳk�_��z��m=-*X���G�B5�Dy�E�<%�[#��vV�%�P���s���ݮ��ˠ:o����a�A��]ʊYQ@�I:�m#���ͬ���8] <����spc�)�4^ξF��>Zy��ԗ��P��Er?���H��Z��IEx�oˢ�6HZ���!���H�����|�/�OQ����ޜ���Tu�A.�p3)�ja��/
���O��Ɋ$)L��9�u�d|`�5#�K�Bm�x�M��Ƃ]V��N�4���3��A����
���� �"���b���i�k#�T�g0���}����q��0���-��r�e ���YR��Q�7Cꮮ��JI�\� �^�>LN�M'2�)�-�q��S��S����6CE��~90TDP(���	�zI_�lXǎ��]�V����l�W�}��c���ygMӴ��*��� ����+�:.�}
f����@���`���a�ל^��r�W�-��k�U� ��f��M��xi���p?�bmu�9V�|�~IV�,����s8r�?n�.���?��+��Kά�;u֠�J_S����?��=�ź[����WC}�����]V��UÝZ���+YꝀխ1��_��e�@Vv!ڄ�P�\h�B���+w�J�=и4`-���w�ec�9����@�z|����=#p���l�m���ݝ��=ëa�Ӗ���iG����ЙK<%�a����M@�~�
6���G3��u���ֶ��U����ʾ����`�7�-�p�YRfq��jp�Y��4x�+��kЉ���0�����ܑh��:�e����ʯI���&��Hpq�h�rl箋�\�X��.gr������ipK���D Sm�乒��qho�h�e��K��u���H'hW(��P�tx�c����wI_=xB=�[R�<n�C$+#�������~���ɗ%�hJ�{}��_�*B�\�V<�鼩wkჼ��^'���!Q'Q���~���\�A��F�G0�)bK��:f	�3P<fc�0@�蟲�'<��{��qV��W�����nMV�1���V����U2�^�����F�Zg�ɿ�u}��&+���W�8����F�%ĿJ/������j�v��0Q�z���A�WC���ӎh�7�s�CԹ=��@�7���#C��;k��h��:}]�c�����Bfm��WP���v>F��煎��/���K�?W�\#!p��
���`*3i!��O�����)�H��N��sޔ�rK�;9#ʤh�C�W OhJ���/�D�+N\����T����0�h�(
u�Ytz�@�q����V%� �v|�����8	�`�Nb�Tf�*��t$�)1�g��.�M]��],�wk�a���R���zb�ċ������'�����4}|�	
����#p�ln��Q?�d���*(Ɩn�4>�[�Y����롘:�}�:����m�6'[����N=�q�S�A���24bv8b}�
B���p9�Y%�g������?�a�T^�� � �c/�K�;����d��48��f&��'/��}�W�؇;�ȥ�M����h�T�/�&����o��.�,hn�P���p�:��<��_dL�����Y�-�Q<�vK�KD������>$4@����Q�=��Y��K�Du�}��1���6y�3��k��ښ���4,M.��x焄�sA?�@�n	�C1��RY�]-!\�tP�uf���;�*��7wO�#��Ut���c��E�|[���l�oI��Z[JL��u �4_�s�����N���d��{�ϱ�hO2U����ǖ8.��I��+��'g���Z�>S�tF3�T���Z�[��ZK@��h1���Fϡm3��k�6�i��T\T��1��U��x�P8#�l_,	�32�\�L��"��ZLcI���O.uY�9Q���yV�g[].�X.��Ɖ��XI!6YU�bd����R�r�P@�N�e�U-©��������~(�f��Z6q�>1B��͸�U�#�L��9�nu�Ƙu��=�m���}�����L�0��H�xy]^s[���i���_UL�8<���T�źʱ�/�P5=9�%����1�`��ߣ�j���P�5ί6��8���V�Sp��cU�W�8������U�!lG�NuO#�K�tI�2N��:��,���4��5���!y�s]���/�t��^Bx]�/�x~y�ΒP��H� �ϣ�K�G�c[,$��,Q��?�@�L�sD�h<��\ZZ�4z��Д����q�~
v���~-�vqa�lU8Vb��Rel�ŋ<,.�Xdr>�FK۫NJ�����^x��8C�?���6Xm�~i���w�n���;p��c��-6����u�u�Z�]�n��W��������J��p�u��l+����%��#avw�5�|�t�*R����
�����aJ�#<-�t7�Ut0��_����A������:��,|�޹4�)�'Y`�P!Y�>�^�$�Uq��*`z-���շůӺ}��WO*�+��`��q"�]��ƕ��Pw���R�j'���w�D��">V����� ;����/����*�=P7�S����Aa�;��]Fr��<	h�E�č=�g"�W<�*�՚Z8Ț!����yQ���k)0��P�V��Dsa������Щ٩��L>	���2�Q�tk���Iw~�q1�斑a˧��u�	��M�8����ֿ�%���ǡ��Ɔ�`�1�KA>7�2��Z���b���fa�K�~7b�MjDt{0/��(<�0��������BH1�z7�� ʢg�@`x�9B��/� �<.�?m/���.��]|/&���o6=-�y�j����#f�����v(����ٱû�o��n��t��t�}$��T�V�$yue���UԘ���8���x.;�3�&��m���r���Ek>88��Q�ы'��f�9cO�Ӹzʖ���e�Z�N&[�Epf^���goS�Rx*�Ş���y�2��Bh��7A\0 ��2�����k�R��J#���Y�C=���W��B�A��(���5ײi#�+c½3q؝�=��&�$s�z�(I$���*D�G"�//�Z���O;
�7��j�O�8�3�mY-2��#d���V�*�7)�pͧ����{��°D�&O�`@�.���b��m�HQ�xڟl�t�p���n@Ҹ�$���
 ����S���v�����1����?�!�&s�ʉ3ר�F�Y4���xz}���$�zJi��Y�h�JȅH���Xb��u6E��KY�)$�)<��6��\����s��@OY���c2��p+�<��x�G��6��}2�. �M���Ǐ�j�<���Bȿx��@:��b��Dd����W<�Z�筄����Ƌ&ȏ��&"�&:��1�/�{%�آv"�;K��Xj�_�ģ!L�J\�MH�7�+��C�ns%�@���/a�0�W���|��V]	A(CS����VJy���1�>���>e�V�ۆ�L.���b��3��Bf���vD��ʎ���Ӟ�v�B73# T!t��T,�y;����ܶ���H�`	SHx.tg���-����Z�*����s���p)���lLU���_�f�Վ�ff���mq8�"�$���ms�2�=������j��L3L�ݕ	n�\Dc��bvD�T�'���#d��=F��,��ٞ�0S�k�`K�r��u%��4R�tm�x�Ri%LN��#0�mlRp;��<Jj�}c�5sY��3W���u���FU�Y����
9��R�@E�5�V^]n�e�Sw<�	O���b�gسj-o���"#d��6�=t�W3�di�nd%�W?B���y2�R�/a��P��}��.3�?�H)�ӹ^إv�<�����~H
e�|�Y���Qc8N���D�2�}_��9���d!�EB�_��ω�7���
t"��0�aJ2b5�f�1��"�r�>��.<]��{���x��Taό"7^�|A�u+ ��A�be�6�jcb���; ��!w��"JB�8{��\ι���s�+?.iw�J��0��F��}����a�2^���3_R����8��&&�T��LT������|��=�۝�"7J{.bH���(u5��*��kF@����B>Y7��	�Zu>I�l�n�$pv]k��m�]{e�O���Q�=�����V�Ry#c��	<�7Ts_W��D�t�����n��7�aP�Dp�9��(��ĶD϶d��X��@��vY�����N$��G�2�-��ť�BG0j"(�J!�l(������ګ��ȤÊfe��+!7��r�)���_���'ITSv��(|�n�
�9���x5RѢ!��(:��v9c_!�G��A�qϬ����M򾞬}�+АoE%���� a�m|�����9Q��&h}$�5��L��K�r�B-]+���\&�*��RY���q�8A���.i�N�c�͘����:0W1C��.��&��dWy�=�p�7l�t��*�Ԙ���_�p��]��3��"1��<��Q��uUf����V�F`�Z6�ƍy�D� L�|�穃�!��H�����POX�	��[�]���4��>���ٱ�� �qR��;��A�7�6y�o(_�PV��C�9�}���KĨ[\�p��#� 	��ʋ��!�����<;	(�c$3̤���g�B_]u�� �p�zIs0'NH8�V�9/w�3Q��at
`@
Y-3)��+3��od����~�� �)
�R�\l����/ܟ.>Y��k����X�[�q��)yg|�^��X�m-HC5w� �R�$�-3]3ؑ� ���fj��|	h�?V�0o�Ae��L/��"������6k@�Bm����.(}�ފ��,��	
��c�y��XX�Z��F#��6K}���]Z��;��V���{1��,� =�x����W8�Kj\�N�jfQ�KĿ�]���eZaQ���I�2�0u��˴u��7��܃H���M.�U�Nr,��(Gɐ�\��ȣQf	ΘƋsz`6�9*�CыҬOJTKK�q�)��\�9+]ʖ�vL:�>	�'t�6cU��+��.����Y+����*���Us	Q���K�bϽG�U��]e�7��1ؘ��	�y����+/z���Tz�-���MO?h�T��9nᢚ}ôc� ������~H6n01�ҳ���x���$���z7����X���g��зU
=̯F�?�:��]�W�{;����*`c�@����XtU+M�qTM�d>�j2�2�;1��XzReC�Eԕ��+��K���-�k��vT[���q�o.RlP��6+(o۞��� $ы�XCS���PnHt@���yRLT����X�����+CU jQ����n	#&�e+��a�\=ĐJ_*T��G!1	�r@KB�p����U=�t��Aޒ��N�$Y�d�ո2��� ����,��b�Y���aDۈ�S�].%�*Vl��P 2�E ~� Ϻ�,lh�.w��ޗ
u]h�Uۼ��E���F�B�4�ܟ��PJ��Fr[���ݼ�0]�-?�ޑF�o�Ɔ�kС�[|��UL_��=�lD�h�h������Iл�2�����/�*ed�;!]���x�ȃ�74�6F ���G�U�~�����E�pTA��Rv5CnI#f�g��5'�x;�m���-�=���M�r���C����ig��k����z�uuL��m^�8(ՠ��@��' OMwk�~G˃��z#j9���O��7�
�݇���I�¶ J�l�E�R���܌+z�F��D9��%v�A�a�$��Nӱvm-�/H>/��|���\"����n2�<��Y�����^)`�F:>����R��/�fk�M�]R�� �(UP�z���(V#��.ȩo�yL�9+x����d�uf{H�e��@��Nz�a^�t`M�x�xm�eӵ�J_��#��3@ƣ�6z�k�K|mꐝ!�� ���^��/��p�>&@
U��$4#9��G~����Y�ߋ\���)įd۾�;v�+�"#���e�+* �L:x���P��/��d�҆3u�>;�v��Gd�{7\��(��~��tN|X�� B�74@�ZRs�~:M�ﯴu�ht]�8�r��5��PFwǒSUZ� 8�����+l�i$�t�)��Nf"�98������+7�
7�}�)h��%C�(�M��}-��Ǟ�y?�N�8���ک�`$' �$��>������p�_��
RD�M�Zt����H�Y?Ϊ��ز�ɲ4�s!i�<6�=��E�$�ЀRO�w0�hJG���P�&oA: ��z��G��ctՏ��O��̘�"�f�����d��w��3}ZtJ��2�ޤϗ���R9�]$������`�(3\g�Ӕ-�	WԢ���z���48)"ZA���WZ�y?�g���T�TgZ� P�}�.�4C�_E~�.f�
�P�&AC땓X�z�;���«o����F��`B�L�K��1En��Yɱ���a9dX�s/��tڗ?�|$�[�٦��b�=*��4��AF-mH�D��Pkv�C(Z��;r��)�)%'�� ϵ(F��6�m�-���ܤ��M�G�>�\w�V{����8�M��q���х���i8E��8�r��_��#7Q��YO�V��7������^bW�X'�Nf�a��a�_��$2������ �Z��o+P�?D�;ɉAU7��P?��ʎ`���Γ�`�Fݖ��^�j��b����S�����n�H���oy�!t��>L�7BU<�i�I��єk�k��Uv�����J�
l�L3��=[�x:��{״t��դ���%��*u�FT��G�u�|S�X�����k���.����%yP�C:Xyt��l?]�PGar�
�w��Kl�L�}h
�Z	ƭ\��V~�n�ҟS%6r�}�D���Ay���}F�=�hu}��c��7��+F�"���S((u�M��(�YJ6�u6�š�//���ũ����G|������g��P����'e�,T���A��59��"����8�V���M]��4샒�9�?���L��T:�`�w��:����~�v�.�����B![|B�Ԃ]ʸ���L{��N��J�7���;��J��h1XO�\��*;.���e�R'�`�١�`���CGc�}�s-���gQ�YO�g�����;a[��hՌ}6��vJyA�BEm�2d}�$�+ԍm��V{6j��MQ� )"���
%J@�: �B�D�aGv��7
&w�·$t�RT�\
h�Y��9J0�}��.���s�Y���=�p/�ֆg�9AahD����ac2&���_&���#�i�yǙ����AZ���2%)��LiJ��~�P�78�lr݋��/i�������i���[��ۋ��տ��.��=3��R�֕�m�����	aN0ِ�ig�ǯ��epy���j�Z��t�<�=-[�\�<�%����dk#ٺ����1y�ز/�m}��VBw�@��"VH0 ��!�
ҋ�ɛ�<mާξė�T��ڄ�7q����X��;>����g� ������H�ا��������A���k�;�h�f�bgU�Ʌ�? �3��Ӡj�?�Z�� �9C�cl�c�N�NMu��6�5�@1+	l����뫦�f�go{��п�iӱ���7����j���y���j��y�F9�<��/���Wl�Q��g�U9d��W���ssH��;�Q9�[�R����Z�W#�R�?&Q�jxśє��+�����	ظyO�|ի��Md�f4�� l&%��'G�ҳi ��ܨ�{�b{��>c�O�M��D;�~�?8�a2?�g�-98U�{#c �[p�N=Ȇ�/�fl��DŦ����@g0�?Iא2~R�; b�y�5��6�j���!��Ǭ� �6��e��v%��fjovx��T��4t]|�$������A�7�`X߲��?�~�ȏ��� k����^�8�ك�me��2|�EcZ@%Z���y�@��O.���ɜ�[t[ʟ�MĽ�Cl'����i�r7A�]h<4�f��*�?FJ�5�]�z��[l֐b�Ā�bX�Y���w�*����b)D?/�P}
�1�*_**��g���2W���N'���4\#@pۜ���F��;�@1 ��k$I���ul����d�g x%)K;upޮ�����n�}yO��io��\�[�5r��3�ś&�[�2"%2uKܖ%�]���-@'�+^wg��w�/��\�_�˪տ'�p�6+�?����"~��IV������m �D��M!G8]��	���3�]KYqڟ{yP��O��UW�� J����:�bqo^�&y��V��C
d�@�-Jr�Yd']Z ��B۷񔿕�\-�͏��)H�P$�O	=�P���_�#%�@yiG�F�@�����,�lʯU �(���f��n64�cJ#k_͘���%z�����7j'�V���aw��N>_�p���
�g�����q�Q��xN|4���2�����{/��w�nV�6;�G�;U���V�:hΕ���.'"��D4��xZp0DF���I{�$���n.	Ŝ�:�G��U���+�I��NV@)�����Z@���Q��8���"6��Τ?�]C�|Y<��-�8R�`oп�⊐~��Y�*��Je�u>��u��nX��*q���*ʶ<�F��R{�c"ku�ګ|_���#Y���<jw�a��<��o=`:{�e�!��fe�>! �@����v-�?fN��V�7�@��N�b-�EhXhj�+��2/���[Yl�W���;��#�}��C��f�G*\X��0�ŕt}��Ye�:\*F��I���"�͏I_e���u����ذ��gC�9W�]�g�%m<�"eG��^�V�e"��/�~�@/P<;z�^t��jP�)r�4B��|
f��q��2KR�W����@rM>O��We?�
����U�	��k�#-E��j�*kk�TXQ>�$π�'�0=�̽�[����\s�_�D��
8�|dqt,o�QvmZR�ZB�]�(��k hpj �II�ж^��?K���]4?����9Wo敲<d�E�Sfw�3�'���~���Փ�`������N�z�t<X��$aQU3�����d����>E��E���$��O[��IQt��(���$(��,<~J;t��Ք�o�1((�y���:��'r��2�;d-�-�p���f�)��	���H6����>l�gU"a?�d&�U|H@�1��g���_픲.?�_��x;Bg��J@"�h���[��|��4MX,i�%�H�T	���'�H���;�1b/�_��0��@�A���B��[a�BH���D0\I@0�q�~}
�9H�nǬ�(�ح��%����nq�'��^fFL��;���#^�=��˟�R�VhীĮ% �ݠ>5�oW�7:ɕ�G�]�xg�7&�^+�?bV�U�ѭ��P������5�]��ͻ��xF���k�_n�	}9���U�>�A�d5�m���dշp���p�\q��4SЫ+���B%���ɘ�'v������ʹ�x�����H.	���G��ʠEsɸ���쌔�E|n�f�Ӫ�Mq����ȲGBi����~�ۓ{�h9k�'�V#�o�ο��������r�L]��Z���,�,�g_T�]3Ⱥ���"��v������Km�*���$�l2}kV0�����d���:o� �$����6�V�h*$s�k��!߁�,���_���s_ip,L?DE�`�ɤ#�x�c�A� �;?��c�	?y ؓM�	��I0ꠈ�H��PǑX�7��	�����ll�ϐ����E@����
��Hk� I*�7`@#ʒg� ��7�S�� U�ǎ��e���n.��'F�;{l��N�U�MN���� ��H��[{��YC�-���� Ni�Y٦�uu���JyԒV�)��A8UN����^'��q�@�T�kj����`�g���
��;��>��vU�������X��9�_qp���\Fx�A?�Nh3��CH����|i��A�⠃F�o�o*'r;eUN������q;�����4���V�H�m��1��kmQ' w3�vg�������3�;���(�@V�0�~�RU�<��7�Z���� T�K��\���r�h��m%�u��XH-���.M���]||`x���k�T9����Ml��j�@��oX�A�8����<��UQ�l�i�ҍ�#)>ۅ��A0�V�ВAKG���pG|�����Q�L@�Yw��gZ��9��=8Գߑq�S.!��^sA���ܬ?�Ү�!�4��_��g���m����y���:G�2P1��IE�y��C�i�&*��q\��A�͓%NAN+�X�x�����Yp���Hj�¤X�ɴw登a��;Mиǆz|3q�Q-�'[kv!ԧ��Ɣ��B@,WF�7am����M��b�����7�����4n��1�ǘiw�uP�=�&�3�����x�4��H�pn����2֋t���
Đ���ޯW���xӁ]"���ĵt7��3崬�c_��y���;%��=ʳ������9ia�Ϝ���8m+�p_�@ɕ�o����³I 8=H��.;KyR�\�E��;<LxF�<"�8�H��D�ϏS���!�q���#iV��/��M�ȧ�cMv~r+���[�V������1(T�mM�%�Veq���@d ��*�}�O��X�rS3�I���k3w����38B;���h��$��J�����9G��
���p1O�V�@�(m=�&���)��E�e�T�d�NҜ�"
ǬN����� ���@�ୄ�U�Q���M�ր(�����ϼ���fL�2%��w�P�ɒd���P��MT;&�UFp��@��n��qi�m�E��ET��@�PܞC�g3� �-���sH��r��5Ӝ#P���l�4��gy�*�Y�֛�;�����_�ގ��,��0}�w�E��ON�t��;�p��H3���*r>T���")nGwJ.7��W��P��_1�kD��6�Ю�q*��2��<��%�k���|�2�T%{.���]�KdK0�Q�@2<���f�T������߿	��7��~�sB(�����nW�D)(��1ޗ7�o[1���
��l�U�V�A]J�4��o ��r|���SJ�{�(�y¾CI�e�L�2�c򳲲��@��*�~WϠ,*��&�%���l7� ��.2�Y�v|��m�<��=�A�aOA^���!q�9�M����wܦ[;�F�fސ���tf�\8I���Z}��8T	�@������i�d�:Z�FfxY�y��Avx6���i�	+0�Is��F4S���1���s^R�����r�;7�����e�j��N)O� ��Ɇ��Pw���b�o��8y�w�Fqn$�W�q�lk^j����t @�
s��I�Hx�	4�C���f��A#�4ܷ�a��}�??#�\f?
%3����)�-��$ύ)ب����/�l�h���y@�E�|�$��}�����P��N�w"sĠhg��d�J��7"I�����n�d��n՘�1}���%��{E�π���c-�þ�tB��8 �$5'0Wa�*;��M��ڴ�{��*�����1`��{.Mf�����h6�^���'ߦ4��$o��� B�C!��K�G�.��{�)`���PR�Nav��4�S�=���<��J�M%P�HނB������^��D,�g{R���P��0X=�b"�F�H�,��xp����5?T��Y���H��Ż�<��|X�Fi\��%d��/\��էj*��l!���V
W��q8$!����Rtkz�O9�/V��	b7��	���9�I�~���o�.��CK\+��ſ���nל�UG#ϧ�Dn�݁�&R���������/�H!�c��5V�a\Dxi�r������ya����'�~$������{/�Y+Ay�|?&�ɸ}���qe�D�Q�-6G�Q"!7+�Vbl��&�^3:�1�<Y/����:>�T�z��ĸ&�v���5�t6:
aɣr��٬�*qT�b[��#��L�"��k����o� و�:>u��������#X+��=��k=}�qP�U]�,��W����W�Kt�c�$~"k�.�[H���-b�#��'�BY�������Ɂٽ�6��Pa�t�~�1�uq�Uʩ�go�`^�}"���X�n�ё���7~�MC��x�C�P%�!����:���J:�'|32j{��kqэ����=߳�ij,��;�0/?���pW��S�Rk��BZg����ߥQ9r�Z歼����U4��W���U�ɹ�;7BJ�y��U1J�m|5������U��T�~�x�C�S(��7.R��lI�/��?8tr���JY�!�����^5�gA/M�8K5������z���P/�w����x Lw����������n4��ܵ-�D�m����߁]K��O4���n����#�-�tqRLWhP��z�<E�Ȭ�X0{/�l�x�/QżOP@i�ĩ�ݡ�~r7��m���cB���r�nL;4��� c�h��VZ��ճ�j��Q1�]�_��&[Zl��C�a!�e+�"������x�}�v�_��1�e.8j���0$���_�m��~[�!��r�!�!t���@�M���Ipk�$�?gj -�(����ۣ��m$ c�ʎs�����HV���'j��I&��H^�a����SS��B�>�h^6��WH��mzW���gĴ⯆�J�Zo������&�f��]��瑹a��/H�e^E�!��}��y�kd�z�~6��%^�<��M�z��.L��\pQ�1��5��QJz�g��+�Pmo�-��d(���-ؽ&��	�_�����6�@��5ʓ�ku��S߀A Ul��62{.Z�j! ��`m�7o������TI����a��7�O<7���������
1z�J�R3�̐�i'F��9���|�����\k�'c�1�����x��T�A?��R"�eD��7g�J�\ʎ�3e�u���o�#����bSv�蛫i�N��l9Oxꖐ���49���Q��B���<�/�^P|[漳z�I��)8��p��΁��P��anaA�_��M�m����{o2�D��B�N�d�8.oaoN'��1k�l~���Q��A��}kLT�P�<MiX �����W��\b�� 0X��8�P��B�>FNt����-��߅� ���zj��?lM��<lj|��v��)Gxj̿�*IT�o"f����y��8Y����&��'��o7��i?$qۑXa>ƨxld��,3�4b�M����&��Y����Y6�?�����Ό��P	�*2;�N5s<�h'4�z��_)z�o�����ޔ3�>$�n�>����0�{I�[I���>X�5$-PZ�{xb��E��-��U;%�!%}K%&�]>?Di���R�k�ۚ3?W��D����:0�'3��eO�l�$U����
 Shڿ��˺�W�V���fApa�4ZNo����4�PJM�Y�]!RV����F)�bq�nW����p���!�C�u�J��z���jW��GY
n�؄�l�anV�����>c�n<�י���d9���p�k�{��j�J�Mj�l�,@-,Gz���$�����"�23�vm:x��#7�tNei���(�
sO��K~�>}4�!�٘й�ʡ��t�\��r����Ȼ���:�6C�Qڳ+��*��`�3n3%^qv���a���W�Da��V`�/5][d��z�mr][~��"|_��}�p�����*��ջ��M��u��EAV8N�l�|M%�WLu^g�;���X�_���'j��]�y ����˓�k��Mdf��Pe=)�v#8W\z�L:�:[2�w�.��=��қs�f�I���k�]�'Pkb�f�8c��i����~I	p���6$e1+���;ݡ�"��c��4Y<��-=��Ep�����,��ō�QjMŸL�Bg7��'����9Hr��].����=��K���/�f����p.�rHb�̸�h�l�[z&�l����_��K���ډ��ܩ���g�Z�BȌ�e&�]�5&�St��mH��)�8��46����VEIO|K�jϺB�(9��C����e�pE' ��#�9�@J�X���M�Wle���Q��80lM3X��7ظ�����v��&���-K׾7�!O���¾_U�3�@xX<�zn���)�7��^"����g�������[<OT�;��U�P _�W��D$����2��i���,��Y��Cuv ���{d�e���)2�A��"o��+yl�fj0�-����GBH�j��Q���y ���g������	�؋(��.s��_Y$���cBMނ��X��(�Le��~��hV6t�ۂ�?������5����c��H+f�. S��y�Zl�iׯ$^�?@*VOÝ�oe��]Uc���Я�=}��3����9�H�v�D��F����_!��=�T�<߇~�����1�X3�>���%�k]~`�`��
JC�
 ��B����X�C�P,���,&˱j+��(�a�V������:u#I�B��Q��A��;v* ��~W6�_h�)���27�4۝�(���=|ny� 0�_F�*�	^�����`��\��~����ЌSr�ɚ��������~JŰ ���Ԇ��h2[c� l#[��!�Ȥ�w �w&��M�f��^"C,�"�=�w��?r��3D��C��H�sL�c�y�ߓ�^��r-�UY=X����G����3$:XEQߋ�w&�s��v䥸`oR�D6a�E��q�0��Y��`����˵%�L�_mF��o+Ą��Æ�k.�e��e�6K6�;0I�kx���1��k�F[�����*Gʭ1�!cJ���y���x�6s\��2#cP�PG},)�D���{sS=�6�_鰒�q�n�I[ϘB���ǅh���5��Cȑ����eGOh(Zδ�������y�l���DN�ƽk���+���Jz��@ဦ�9S�o�&�N�x@�],Bf{�V_�;v.*9t��Yn����\AA�g�ib���|��8�I�koM3���5d��P�o�V�θ�����M崲/�%�3����-e�9Lm� f�$J�j�o�i&�s���Q��C��7G�����S�4ޗ"b�U�N-ԁ#qF�h�h���f%��%�h0e�"͑��gv�����o��6�d�Ɔtf���Ea����_��ud5��OM��6��U�OͣApvU�yW��*�ܗ�������åZl�5n3��N�ĤW��|*N��Kv�,Sg��EZ���Q�H�V^��0Mi�Ҋ*g�-���0��>��kk  6����&1}�e�T�_q^��>2i�;wz������J/��M��pG?a��&�)�$��ұ�ӎ��Ї]>w�GǮ�ri�<�����=L�#��~Rd����<@���*�R�D;aW'��c��3������σ;����m�gǾ^�˓QڨW����e��R�LO`��K6!��Gc�)���@H���{��E��,�cq�g*�@��u%	M�y��x5D��慎��M~����Rֱ��꿿d1g��*��p���*�`����]�U�W9��k�?8i��
�:g����
`0Z���c��EE�B5��b��AB���Mߒd� ��Ku/T����J`�?�#϶gg�ya��$�F!ܛ"����Q^st%w3{g}���ޑ����k�)��l�����p��%DVh�R3��mC�I�U��=&�CA���J��/[4�T���Z�k����"5���s�|��7,tt�~�G���q�7�Hɏ����~���5�[A�'�Ii�$L�k㇬&���(4��<[��$����ܶ�ɹ�r���}tHl�(�����F�]��Q�^�y�6��������N��l� �a��Z������o�ԭxCc*#6�e��(��Q��p��U
���y}�8h��2A�[d�q��N� ڔV�5���@��_�����-����e��B��C16Ϋ�QiXx�f�4p��:��M���{, ��W���Ӏ�o=�Ew����A��͋ԩ��Y-�Ⱥ�Ǹ���Oy�����Ls?����asb�;���i-]�K���"ȅ�u�aۍ����6�~X��5�%k�P�=ͼ�05�j�p��k��=���!���]�J��
�0����l9)&ͬ��zO��+�uU's뫆s����ߠ���́׸���g����#�GN���`K�X�ч�����OAWRl�3�L��#�Z�W-D$��7򬭸�RVJ�W�_�U֗��v|@Gծ��'�eQQb�*��7a�b�fl�j���6��
Z����`q��zC��G-�u�uk�������n��|5���<�:$}AT)=�6��sE�:H� ��3���O������ʡ�͞�.'��}�r5M�����1�ᙝ�����9I�������8_�1{��<�'�s�XG�k�E�������0ƃ �6��M��sK�HKߛ��^S,�"<��q���4�H�g
N��X���*��xbLC=,�/�����/����+nw�׋�C�2�\[X%q���)L~�E���0��=&�4�?�Ƭl[�鱢BĵT㵰�TN�	�H5��f�o<�ڼ�s�g(�2Y�,ֶ���!�Y]�����#�����j*�_3��쿂	�fk�e��"�W����W���5O���O���>6	uI���B�pR̬I��G���6��j�8��S�z�ݝ�V41p�rƠBo��o=(k�t���mȭ�
3�,�xZ|�6S�O�_:�;"@{9U]Pu�^r�w3��>��.N4o�Ǳ���̍@�	}��j�G'Y���l��]bνք�e{��G�{q�f� (kZ�ݦ�� ��3����H4 R�K���Z���W��|]� ����N��V� ���N�N<�UG�ЫE����3�������" ���6��:�~�6뎹���;��B����۱���|�r�@j5��JN���C���J��<Sq��h~���h��H��!y�RϡǢn�W��^9c�����8�������,��͖��D�-ٍe�)+V��`eP�_%L^ L��w�۰�ܶ빇�܏|ĳ��M��;G�6��G�K+e.!�v�o����n�b���b����E��p!l1)Y$��y���m/m�V�sU0�@��i '#څ����I��?>�RD�v_����8AS��������u���S��c�ĝ.x_~K�G�O,�ҏ���}۶VCU��ĉZ�hq��;�d"�!�5��?N
��9_�l��t+>/�*��;o��Zu�I�0�񰴖��[�R�3>��ȇ�V��$���r��x���'3���@3� [J��$<ԋ-� ~[%;�,U��*���ݏ2[t��o�8S��S�v���p7�+ɶ�/0��ѡQ��&�P�'4���k1�5��@V�{{�k��\})#d���o���+9��d[�8aau}��'S�C�ؐҌo���ܓ�6+S�v�yUЯ���鰱�!v{�J�*M�V$<�%A�p3ať"�����ó7���ߦ⟃���Tb��'���v5�D�>:fB�l�*�݀����#~��{rI��Ȓ{�!��S.�H	�f[��`�p�i2Z���CLv��y�f���nyb���/%����i]�ƒ��^Q��e�;Zl���>Ԑ���n���=6Q�W����h��N�kƠ���%%k�����`k��.�� ���n���W����1}�b�C��Y�{Թ$��
�<K�4�86�>�ڗ��H���٤�ߑW�����������|GM
;���e�;�kj%=�O��Ha���i>�2i�@�${���-ph�V�X�VPA���są+F[��a>� �Ru��[S�|��Pwk�;8�sGV��.J�1�B�bu��`M�w���P��Q� �ğ�����+�QJ�4-)F����,��@���l3Z�%0��z��BK�����]�J�4��[��T� >%_Qr:/�BZg8�k�(/6�䙔2C"G��t��at�|'u]ֱ,�6����f�Y�b������fd ��ƪ~/��e#�*��5o$�E,�xjeV��y���yߨ|��m���v�F��Ң�cJ ���E����4ީW�l'Oj�ʵv𥈊7�c&���Hw�6Y���m�ɉ���]���y`uP7��w](�j����t���yڨs#*r�Oi�DHV�x��@j[����L%��4��0���az�wh_��_��(��*��5���۶J�վ��?��G���R�;㽮��[o�Vo6>7�K���NP�h�)�}���7l��g��r�s�N |��o�<�V=��/Ov����|���\���ni4��߿�yI������m�|L۳zc��"����}e�"FIU�>����o�j��0�mQ	ē!wr�+ǇyspuީSɮ8͌d�S�0BO��/𑼰|�,ag4}dc�b�y�J�@5/{&}��Cch�����	�y�Aj��,/��=��R�gL�7��~tN�}�펼Z�<F ���L�VJ��+��C��H�L���w�f�>�zܛm���}���;zy�v���b������ӔVK�Rh�E��^ܡ�דi�L��6�K�JVV�v=�Ὗz���1�ܯ(���_�a���'��� �=�ٷJ�Ei���2��+�rȗud`=ˁ�W2�'�AK������b���?�	r*��T������'0[0(�^�<��b�uHg9��+4?� 1�0?�^3x=e��{mc�Z�\zh��a��A��`ڣߡ��/b�"��H"���Ӝ�t$�N��Ī���r9�ǥ�w�Ƿ����3����2�����s1W�I�6�A�Ѯ<�&�OR�|����Y��8��-*aU�-��D��{�s�u�Ɵ��di�&�����F8���٧H�poڊ�7��{v_3�^�E5d����ry�o<��#��>�L'��l}gL��m爎^w_԰{�@x�#����o�_�NdnJ�����9���q�`��օ�wW{�m��'�d�˼�6��Z4��0�|QC|��0s�H/�2��/���S�^r<�Gw	��Ʒ��S��(ʡ��O�+4����--T�Ne��i_�L�Ma	m��o[��D���(�y�}��-Ah�A�]���6 D(��s@J$>!{����?ؚ���X��Co��0\{�}�^���(�\Ea��gL�d������#�O[~n��W��=�Ig��	fpN�ݓ�t���J{* |5̓����b������z�H�|���8��De,���?��oc����� x&�
T�֩�KE���6����%���>�p�"��6r��l֤:	���*><gG�lߪg�����]�Mob
�4��tF6���k R��m*���٬v��o���t]9s}Ηnd�����㢺��t��(�-Ұm�/
}%�7�?ZF�۟�� ��BW�`eO����Y����� �-�����!��$r!2��<�ܠ]M�Y �/���K�
ڴ�����u�B���� ��Q	3�"��f��� ���\�D��fތB~�B�  Hfnlȉ��W�bﲀ|kt�	 C���@���x��uA|f�ɦB��H���[�q�'�ƴ��`\_�����ݶ���'O` E�$��7�7� �e'��2��Ge�f�"�:s4S�Fc���(nxi����R�Xڅ�O�,�v�TJON�D5���+���[P��!Eh�řN-E��nE��n���[����懺��ך�)&���0��ȁ���K�,�U�2@gz����w&Q�T?8;}�?+ƶ�
���ǧZ���ڌ�:����.��]���]B�hm���\C �z�K�@�Z }�d^����X	�*Z���׸1~��,��n���ۜ�����
oG9���%mC#�Le�a��v�9y����gG�1ڣo��fQ��`�?g�A)�	l�S3�`V;�gƾR�%�Ԥ���s;�[��>MF�R|�����n��=��ձ�S��.k�L$Y������M���ӆh�bq :��.?�3��7Uq�R/|���d��&Ŋ�@%]w$���<�������"��g�K�c}IM��3�
@�u�,��n�[7�o�|����e��38���������c@��r�z6z�?
ܚ$��:��=�`�2��ɡ�ǖtZ�R�s-f�?S-'�j�� e �3��MΫ78fC����?ux;zU��h�1*�!��hl�
��ꊈ1�5�Ŕ�����d���#::[,���J	��[J�AP�t(��b��n/ ���H�쿬��mc��!^�'�@��G��YX�>L�F���[�b5����+����}��k�G�~5FIs���B�}&�,���ʺ
�Ǻ�0�C��(��������V��7?��<��m^�6�����v[@�j<z� ����\��f�RG��ӆ-4e��|�֘�au�)X�����[5Q�U�3ʨ
���]mT�g��|ҫQ�������0������S �l;˞�E��W��R�4U蘆m8��n�H��.�<�޻�>��ݔz�h��'z��=�;0�K(�!�+	#	ٽ5��R����g^���c3fy�X��a���(K1aB��V�
<s���pۥƼ��;��������	��Xm����'��8wՏ�;a��6�e�hp~�	��Z��h���������b�j��R�[W�'�H�F������8&$����x�w��3��� �^U��p�-5�X�/�	�9'�%�A�C�}��9F=?�7��F_�Sft^uԦ�06�s6�tѢ��0��b�;�j��e:r�gPD1���2��D��xn�l��^&ƃ}8�w� O� �.��Cv����(7��A�C#��(S� �p���F��Li,4�:%���ᦝFS�gYX�0�`��Edy�L�{���ex��k���sQѥT?�q���Z?�I�y�1���C_j�v��;Қ�F[p��Y�NٲA�ϑu+*QBӳri����>	�r�K��*��|r�%rPQkOٍ/}/��ɮ8)V5��V���?�YjŁ[*P܀���֚�}����O��pz6��z#T���۬y����2Jb��K i0_�������:�4+���l����ٮū�-G���5�j8���x0d�nk�ɟGh�����4Z3L�m��S'����׮��y:��Д������G�_�H_��Rw].���{���>�$?R��v��V����ak��s��6�.����ƦE}y�{���T�Ђs=+S�0���Thɾa0�Z��DM�s"z��U��o	)�n_����k��}�=����,�0��'�(��
�\=4�I[ݕ�I��*�T\��È�`j��Ht�,a���)�_����V�I���S�0Vb)�q�"c�1���p�DX.
2�{�ޮ��h�h�U@]Y+>��(:{.5.Lr$w�
Nu���������[{�X�f~D#T�ē�D|��H�kD1^q���_���_�L����mw�GǰK����t�E��
�^���r@��1J��V;4���������Ή������+� ���=SS�v��V���m1'6Wq��@�� �h���c#�G����|�C��Y�S�P9��-8���l�ۧZW�:�����dh:���zQ����`\�à�8��mO?!k
���oK�ؾ��8�a�Y��vzq���a��v�<�|�9����wi�~�.gZq[9'���.6zQ[����������E�'(u�*{*�X��l)ꖂʆ"���v�i_�4eb�sԬ��统��i����bͱ6��e��=���ꡋP��Y0a�(�6�&�أ�!��ϑ�%_�>9D����aDpq�(�򍈁mmy.(�9M3��L��� ���7;��k�su�])���(�V@8E�M�3���d��2�50��^����@����d$����c� �#=�J�k�2�`rB�[X?�XMy{����u�����Q8������\9��XG�!����e��Ki��� ���PB9��5�����H�&�̘ܗR���>^n�\Q~��Cf ɱj���u��W@��X�c9ˁ�4<�#Ⱦ��k��A��I �@�8ޏ���8�{?vg���᳞���]�ť�;%h��E\c��(�%���IiYH�+��$��WV��]E�jo}�k�s���*���MkMS蹵o��pߠTx�3ƞ��9�d�g+1����됥S��=-߻1VCy�m�0��W�����SӾ�X/S�����n
��Ch$��RTZ��|�)����v��H�$v��Y�|�5k�/D�`����h^'t�,�A�e;]�3�C���왺5�s��C���'v2zN2��L:��T۪�*��$O��?�@���0J�1�b���bv`}����v;F�|z���(�����5��p7��Pu�	�ՙ0�9����]'�Y.5A���L��h�p^}����o�Ur�=#�����#�r�`d���\x?B^Lq��qy#̵N^����:8:��$��	C+��r4H�}0�Y�V���S���@�>eϧ~�9��~4Ts���$8�H�"	�,E�zw-t6�$���H��Z�,¦��-;g��nKE ��OG&�G�Z2�� �Z�d��x��Ĥ �l0�$�݉C�I�.��=F�v�c+枆$���h��z���-	R����|�Ƕ��p�!_]z�Ҝ��̴
�Mw�<�0�����쳻�=5z`�1����r�5ahwXN���crr5E���S�IcX�6���?���oZ��m���,'֏9�u��~l+/����L���_Xj�$k'�oJ��Q�m?n��DJׇ$^�`2^�#v��[�����BC:H�>-����J@��U+NN���;��I0�A@���+��e4z-�,��nT����DMa�dE�+�,�|1��UV�p���d��QΒ�����f���H�9�$KBP��+uxK|�c��(��pB���EA��2�]L�}O�z���؅���;�N�-"MA=6׊�l�.ٹ����+r��kc�}�Z���Y�x�l
Q']&�3����n�\�MÄxVM�Dz׹�鰠D�U��S���A�e�@̇�VGmS�s��wMکG�+�M �qG��v����[�^�΂��֪D��_��L�21>�c���l7�ʣ��s{�Gw��7\R�֎2���Cp���'6��H�z�_F�=؀�E�h�f2�S���[�{zT����]x�x���',"�:)���&g�.X�}Xa�����"{�q�K·���B.�8�fɒ�K@+��|_�k��|x0VΪh%��GE�1�ߡ�'n����I7�t�� ���)5���C�19�p�:�_�~�K��0*'�0l}�f�Xdu�yD���Ws2K�����]��� ���u*�:�0C��$ ��v�PHKlN���O�Ys��|n����HH�ȃNr]�m9ǜ�3{�RV6�#u�b��>l�%~���K�+m��'���~��X�ܘ(_��Xf�G�������FH�4�jL~_+����]s����K��+i$,-���5��Z(�e�ǋ%ҹ�i/��y? ��*:v'�ɐ�d��{�')��f3o���Fcؑ�+�z�~3��>+n �⮼x�ҠXo���Vd]\C w[a�X4㵐!YDk����	/�ܻ�Jwx߾��%���E��ԣ_�'��YǶ`s\-��+l��__��=�y�l�z$�Ds�CmAR)�(�2�'D}��#�7�����|3�U�u���B&Yj���Z~7E��E�^,��MV�MH�F&N�l��X������͕�Ɇ�i�����`M�.W��t[�g�>� �uA:�t2��.)7��!_�)��BC���=ۑ��M��/�Cp\�������NxZ���(b�A�D�󍓁��������EV��1�y�9�'q����4�b�@�_  ��bF�Dd|�u49��vNd�����c�O˚��14<L�T��N8��h��`F�ta8j���j�G�����ȺB&�>?
�ʁ�;�N����(hQ��T^n�Xz.q�
S�$��]�s6 ��+��t�<=����sE�Nb�肮*�E���i��g���ø�|����^1�p���|��̹�O`Rs+[�c;�����g�p��k%2�ĝI�n-����v�HN/_8`�O`m��G?��B�92��zc:+��".�[�:�q�yR����.vq����0åo����YJ�g_=���!`�i/�ki0,i(1b6�&���^r���J�~V�3��y0MjQ=��z�!9�LG�'ʚ�ys����g%�Ճ������e~�p�1��k�8�\�%~r�� 3gs�" ��lE����*�Q�":�F���1A.�LB�c״��������pe�7JK�0x]�%���YY^𼴲RCi5#�ɴhbZ��``�zڗ�H^�sfC���r?{�#�k_�и��D�5��kU��ݠ9�J�e��ӻ0�#w�^��竖�T�0�1���F	�8;��]=�r �V�S
�y���v ;����=X�E2�}<ìC�V��n�ڰtA�!�Y.@D�bmw���|�{�F��*I8�B0�9��3)6��,�6f�[����;���A3H�#�s�X'}��	��w��ɭ$��"�"��zܚ�}�-4�o�e�8��Т����f�o�O��	=�#]��C����o��/�1ן�x8 Q�0:��"��FلJ��q[�;ۆ��dhh1���������@�Y��<>�ȵMz(�Y>p�U�Tӫ��,F��T�p������u�!��i��RF�6U�-� �g����kϙ"\�Jƌ��ņ��J������J}�+��*�����x���"`3p�X5�[���n2��8��� ��b`ooe���[Z�i��>U-�z}� �*�uڴ�MJ�߱̏)�C������K�(�����&g' +�zшKƫ����	�#)l�}T��)@b�YH���ӌ 敏�@�t�ga�;�`m3fa|o�#��;H��P�~%LN�D�ς��\ل�C�aY!�_��!a�=vU�!m̍����9B���D��h��f9A���n�(�ݡ���0��H�"�J����TL[�S���R�����$d�p����W|�Y�K8�^'�����_0v6�\��9��OD�k� ��ca�)�1Pn�-�{���o��:���Vl�:Aʶ}Y���ٿ���<_M�DB�Y��k��v��]9j?_?ې�����
l��K\c�~�sW�b�F7�c�yf�� =�=���fX<4H��� ��"3븱-=ݒ����K�����)�W�k���oi
�5|���E{K��+��kW�T������}2J�w���g'Q���7R�,Ky@Ag�I����D F-I	�m�<nF��%x4Jg��ʯ�� S<]/D�G�F���Ë�
�u��Z���\�6|?��� 4��tp��H@��r�:ňfvC�R��<�"�)nz|a��7��NJ;��q��>�s�gd������X�w@�l/�(����O껞"��x��stXL4�Pr���b��$��ζ���-�f!���2$�,��<�a-[�m�Obr�E�ތ�%˰��h����4�fQhB�m��oN�S�!>��М��@����0�T	�@��]ÐaX'M��PU9��wx�y
ң�Qk�����!���zջ�Mq�\#TsB�������j�[��Zx�L
����S G�R�:� ~?ȹ�����BK�մ&C�����j%�?�F�7a�hP�l�<'��ۉ@��H���M܋���ɯ�J/����
�w���a��?���G~ٌ5�����i58]$N%�C���;b|�+�C$0-����	~�<��/���f:�)C�n��4�K{����G[,v�b���U�^����x�8�f
��e!&ez�N�	E��=gs��nZ�,S�f���(�z�U��7��4��Zh[ղ*��\���C��ż��v��x��&D���ؒ�n��V��Lr���q�>T��f
��:��_g� ��"@8�j{Ӽ̃;|O5�2�ؘ�/�D`���HVN�\Ca�� �	.����6'�.K0}��@��@���_^~y~������O������e�_��:�Jo���ʣx��)IL�\�1�'&�$+��n��P��i�n��W����bu8��݈��7�%x �A1���l�������N��� �ۣg��E-�pX�z� Ahȯ�����!X��O�gw"0�������/�1S?t�f`}��O���k"�vY�j���	�i�,G�Jߣ��h"|%$y����}�͎[��L�m�J�o{�;G��W�a�bÔ�����|��ơ�-c�3zHdޛ�9� +���	��;�3�&�g�n�9�b!�v�3!6y�GC�&_FQ���ǘ��@���z}��TG��>L�t^pt�	Wnt �߽ų�p۰�0f���Htv$n۫�	�g�»��IJ�<X��-����X�ѡAԊN����ǹ{��Z$���ǂ�'6��Fv~c�:.eI*,�ʯk�Ӌ&��Q��U5!�]�U�H�|�e v��7������|�Ta����p�EV	�+o�)�;c���Υ ̊��w�Vr�f�[0��*���rFW����L/���v��Β`T��M��T��0�"�[��[�3�wc��s�)�]��o[�\T�߯�å�f�B��!����/܍s,-������]r��*�Q�jq3S���y�`����ڢ�~�JGL�>z���X�IN�� �Ok�@%�2��Y���o�n�3)�@_����z��+�U�C9\��G�&)J�Ra;y����њ��zԐ1G7��
�|�i�@&�oܝ��f�����GiH��D�n,R�~�\�M=s�_	+'ř�²^�BO�׼���+�+�XMGVQ����rʁ�W����P(�lz�q�QI�=�W*$�9�P�1�)ĀK��yC�U�D�I�X�q1��{Mt������I�>F�q%�����~o&�u��_�M�O��'���
h��5[ $/6	�=�R��D����mhs�����D@��'A ���,حO.��B�M�?u�a����S"��i����	M,ޥ�XG�����sB' o'�07�K
�3Ia��.�4< ,ŖFKv��t�̥�-�G<�D��>��#��m��KI�bwBIڅ�{q5L�K��i�=���!�������������Z�����J��t��5B���aŎ�r�(���:*�<L�?ETD�8I}Q+)_��JzЖ��tQ|DZ�#�X��-E�bǃ<�LF��)��		��f>�)�'2�r�-m�ܖN���������m�R|a����|����շ��P0}2?3�03ܹ�+�h�;=ކ�=��wp��ϓ�?*e�09����%Q��0?Ehx�ֵ5�����Y��AâU@�_�xgk��,�����h��L?P���`���5<x̓��TD�Wc	��j�/��KJ���	diTD���Sp�&W��ğ:^'�Ϭ��o��p��M�JS.�c��m���j�(���cS��� wP	���1��Om��:��j�>t�A� ��+_��ӊ[�=M�|��8�3:/l�Ƴ 7���R�lZƪ�P��_ޅ͟�l�����c��@��P�f�����0�f`?��� �| Ųɱ]T0m��C�:-`p$�m��oJ�q݅=b�|���_��A1�0�Y(���iCٌo��g4�;U&v�+O��4C�M���0��A�ݎ�;���+�I3:�XAk�+F��ld]�yL���T�r��N�R��3����h�K���κ�����14u�$=>HQB�EU�+!�X���u�����J�A��D��9s<������#v�g���@�˸9*�f�"qkg3�k��k�/Ń�a�\0�A�w}l��[&(�`5�90ܬ�&N�\��9M�X)��5��j��í�{$K<㐖 վ��<��L4���7���L @4y�k�[Z!�| �0[g���块�N+�g�Kꍩ����?@��Q����	c�n��5�����Y�cxr[6�����Og	w��׺q}�#��j�+}@u]����01��
/��ժ#�Ҁ7�;�9���C\�Bs-1	���ÍF��B���'5���_�^��ֶ�h������]������n�y(�$|G<���ʙ�~���*HV�'�R(G5��)���t����E�U7���Z&�V,J�a�H�%1 ~]N�"Vcz��[rU˭����|nd�f�H�wl;�PF����|}�<Y���iB��l�80��m{�7��n������2$R�!�a�תc+��C���v.��:��9<����YB���i��>�ɶ��N��(�w�y����b?�>�gl '�C���]$��f�z���C�S�\K����i ��+��$�q��Я@�'��F�Q���[��'i�0;��U�5;Cc�o�ݙ�-�A�N����b���mt1C���-v� �w����c����+cLe��{�l�$�����cYx��Cҙ�;��~��R�^�VBolT1� �WVK$UA�2�ȃ�Ԇ`�;v�����$+0�7l��2�0��ȋ���,U
\�x�[G�XR~F���0��щ�|�^Mr����H��E���� �T��'��ѽ���iq�.�(U�P�W��ށ��q�%U��9o�$DGI� I&ź��*�*߷��xβ�s)�����[ђ|��fy�b浰׬���aCcG4�5m�F*���IAI���{:��@���7C�v������ޙ���̥Tv�?I\�2;�9֋X'���@�����ɱ�'r�+׫$�� X�X��*9��dF:M$��|�k�2gD	��Jc"%����
�eb��R�z_K?������JPJ�������l��q$<p�0s]L:&*	r�ƃ�r��gj�@K��u)�#E���	\��(1�C�M�d�9��{��i½���S�I�H�wr�8?>u�y�Ob�1��x���ps%���P��-���C��m���ev�\	��ܦ*'�5)����/�-����������ŇD�5|�#�e��� �T�5���ű�?���7���YyD����F�/��˥�티����8nI�O8}�T(�oc��Q�Q�Kʄ����R	���oA�}+����7<�~������l����u<�~y���oĈ?qH@8{m��	�}���i�:9hr��<F\�-_A��~b�'�R�Z��BtyGC���B_�~v+]�51���LZ376�����5%`Kv8u"m/Wz�׽������D�ǈ�s��uȲ���z��n�\���t�j�a� ���!�vw��j���wLL��4���K��ĸ�ƙL���`T3�`��Fe�r�������҇�0
!���<h��cx��R�n��"G��q�"��S?��6t���,qȹ]��X�ј^�\Sp?���;�;�2��4���|,��X��q���#	�;#� �V���o��)�Z�W��y@y��M��^���;�S��-����q�졤��ND[5�⿕�SO���07��� {2�]�R�|���[~4�c�FWbi�3z��l��ҵa�P���V�|.�����HX��E<:V�����}�z������-`�6.���Ы�y���E�6O2 �!t+T�
���{�#ڍz���dP�Aԙ�6G�d\H^�H$����Ǻw��g�0�l���)WJ���n&G�����ܠ�1개��N�/Wmdn3����G,�pG��'_��o
X�f��
�h�s��?��Jg)㧯K��vc� ���b�q|Gg���2�.J��0�؆b�F"�+�j��N߂��^:�h������\֝�Z(�|�b�0xPDPSc��+�+`������%OMڏ;�������BP5P��~~w�OfG*��k����:���L���l�~JwTl��}k�+G�#>��}� �E�UW�'����U�b[	969�7��狒��rxo�i��&Go��x�qr��F�'7����@Q��K����t��������U�Q��A��ʸ ���.��=8�h� f��[Fw���$�c�����8!牕���0�ۣ.�Y��Z9y�[���ٕ��&
�N�0��,��M)��H��ǋ�Ԙ+�]�)�bu +L�S�zq=A�� ��\-�g���.��ݒ��Ya:Eh�5�#�Bj�Q���4��)�fO����3'gՇF>�ZC�p9�Rl�3��b��̌Ȟ����Wt�3L̤M�x>r��"�>?!r�w�~�?��q�~|�>��QRƺ:|�S�*P�~��3����oI;�L#�t�M�&�nJL~��VU�+��"XI55�~�)AI �fX�=��@w���D�w��x��4�7ƪ�g�����:*��:X�c�$ �_���|�*O��G�alK��*5��Ef�#�АF��K���ܰ��N�2�d�b��BĔ� '�����+�/��1ӣ��}ÍNx�B��iG�(�8�����[�ݔ�B����S��G!\��(�0C�`��쟲���jo�&b��̙�@��0JG�̓�Tʴ홴;��T���E.��vH�&��0�7�b��1}}�YG&��+��Q�u��[���������nAW*NI`cW�<�-i[�75�A$n����@�n뛒ZN�bIܘ������o���ʓ�M�� V�b���އ�Mo����ϝ~!Р8�D��i����l����`�#�Dm��� �?��Bk�.�u�2�������g����gxru���g̵�QfE��je��HF�f|Q0�\��̅#��JN ���J)���C�&r��'	+gC�ۖ�HQ�;w;��ѱ����'���8�S��tg�tlKX_J���(��5���qx�i��r;T�$99�o32BTj��=��A��Z�/��t1H,n�>��������%��&�E�˛w��΢L�O�fOetI"Z'�Q�tp�V3@>�o��Aߩ�?�����:�TeY)AHůȾ��)����ا�&�1*[e����Uz~}�n)����^�IO}�����W0���Tl�Ʋ���x�r������?i,�s��xx�`5��#ǒ�8�ߝ�@0���g%R���ܑ�e9
�Flz�2�D�/�S:�$,A8����b�=�Y���7{�:�)G�"�gC�㵬f��SN�ӌȏ�p�׫)y�d���l�7.�g_��z�D������,������T_�J���i.@4� �{��Š$C�1R�?�K���=7'ۡ�߂H��O���aZh}G���l��������n�y�q�r61Rn����C2�X$8���)W�VT�r-��ȳ�L6����'���PŃl3WG�j��S��N����oL�OmU�읋C$H�n4=����]��B�+��}1s�xE<��M�&[��6Y\ۚ�Z�J\�r���S������Hx#g3���X6 s'��iw����dcJ��������
qҿ����:^(�v�bx�8Ĺu�h/I���zE��`��;L����+F���4<ͦ��T�ܻO�_�f�찖���԰�@�XU��Ih�q�`�D�D��j�W+ݮɗ��P�ZhyEq�V�Y���xo�	�M��0;�S3� ��6�<�Ei	��c[m��o�|���A��Lǆ�{�#@��H�����q��0ދ��{F|-@�@�D�(��b���*���U��Q���]��g
��O8l���!]���x|Kj��M ��&�x[9�I���m|�>K�L1�"}�sJw���[o��'0ɮţqE�Xa@p��>���lu-���%Q�@�M>K1�L�v<+�6�v�}>�G9`�g�+S�\*j������ѵ�!����Xkϫ"�ߍE__�O�V�I��;c,��$S''L�J�����oK��v������x8�п�,�w���i�L<���3�!�tSj��/7B㞕�̩�N���exL&�/VYB
�&���x���Q�#iot�@���; j���8���k/Ra���8m�' ��E0��I����DA��d}���J��݌�q��j�A�����s�C ��xߚ�{|�+�̓�M��Kt�eMМ;٭�E����p8w'��_N�اo�����;��7W��E��@�o�X�P5,��Ṍ���44&��F�g����ʶy2�I�o=A����B�MrGco��9�G��J�s���A$�� �+��R�Za};?��<5����>�1A__*V������<�F�o�*�șُL�Ϙ'j}� nC|�vrD��o�#��r�������k��]��_��:0�X���c�<�$�I���/S��e��}�p�<�_���Ҳ��4WrF�-1��}���|�W�8j�$�ˈ�tdkly9QK�N��35(�r1��ކ�a�i�T���fƺn�U���8_�)-�w6��~W�X�v�E5oz)W=I4���2�jgk*?�;��$��i�E"a�N�|y�.+��%{��Ԑ�����P�f�x�������L�W��7�����a�~01��Ս���F��;��mO�ْ����DlG�!��u9�z�̙�dٺ�7ҥ��r����Л�s�{�FN� /i)�;�n�Xu8c�l���lPZ�Fe�I^�Š��򼗸�'b��.%���.aK7*j���qJ�:;��ӹs��|5KS�$�+�ϟ�4(�$e{�=QVՒ�9jȾ<f��N�����qE��y�w:��};�8 �#���Ona�n&!S��M�i.���0�L��f\T�7@�� �����I�v
��(��c>E7�n�	%]��%E��2�#�G���:�JU��9�x��8���Tƾi�bD�1�Bh�=x����Mb�RT5m$k`���B4b���/�3��[���C�O�]���mb�Η��3G[.���ו�:�=1��:����ȫ�Y�1�l�> -�/|x�t���Y�W����Y��]�ߍ2jF�d%��]�ϧ84�V�s�S��b=c�۩1���Y�)4T�uN��9|]��[�������r�.�uzʸ*2��6|V��B�**�v\d4=���3����4|�Z�#A�"���z-�3�C��Q	�Y��W\�إ�$@�*�؞�@�����X�h:��{t����D]�x���U�_�8��Yo#�T+^���䝁G�D���'�ܞ�j�)Z4�3vՕ���X�`riߥ���m�[�Y�4�u�����>���V~H��G�$�r�>��a�0-��D��~{k::���!��S>߇�L�C9&�eV��4�7�X|���m��hpj��AM��I��mh�a�ρ��d�xwH3�����8Z����˶�p�a=�4�)�"�EEG"An'�0�\go�	�5�N�x��L ��Z�w�k�ҽ�+9e���9�w�^u�c�s����<)�HS
P��G��s��>�PZ7o����1N�����w�o"�W�gn�OS�K;ϖ�g~�p��vx�cm�π ��X���V���G
�����{��&�W�(�uϏK���xq.����������
���$�;ype��u �������0�R���k��t*<�;����fjn��c�\�Ò���E���/�`�s�fS�*�����J�_��,�+�!�*4gi��T�j�`�o���u!Jk��Ԏ�����ϋ�!T���g�q�j�@�ʻH �I$��� ��W� �%��Dv�M;+�a����z:;�g��N3�rN���֝�����:gBr	�4�H