��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��V�^�Zð5-{=�8p؍� �]I$�/L=���|�+'B�����c�*wZ}z:m��G�WJW�0cYb(+i��{�3%Dp�$=灆#����3�E���5/,�.��F�� �A�u�@�/5OA�E�o7skeEp`��1��a��4y�����HUK������Ɖ[ft��ۼ>�1ڼ�K�Ir5�����p�b>�֦Z�/U���1v����T�Ί�Ҙ�sg�%;Q��Z��C:TW՘�\Qѯ�p�m��ơB@.�C�[�(e,��X�%�ϖ]����%���T�eJh�0�&G��Cm��r�i��6-��{�zx
�Ý��Bf�d�z�o�Q�7N��}mݾ��G���O��;�Q����!%j�`{�!�{��4��3�=��巴Hn�LD<�B	[��x�\sR.��{�i_�ro���;���&��	w��}�d�2�nK3*�{���D�b�+�D��vz?����R�>���J}��� �h���)Hg���e^���~##��/i����7?n��r��hV�VT�����Ny�2�j%�E(|$�P�V�5�j�7�|�Ox}g���&�-�p���^*�
H�1�[N"$��:��
����3����nZ�K���;�~�d�s�HDnvf�,SpMW�x��vD4^�s��B[U&�aQH)����mc"����XjM궯H�����]k�F���:قݼ�Rథ66J�<�p�`�y%W�b���-VT�@��ڋ��t��RS�c2��*̝�3�Ӫ��u�/sO��Hf�m���p���!ŵc�"4�����@���|��J,�ꟗ� 5�L�s�-٬��OY���O_~�`?*���݁>�����Nޏ�LكY�#�p���A��Oi���H�q���Qv�����Z,���jP�R�fcB����zY	��ϡ���G��5�(�?E�<�죽3ѳ���Qg��yv�ź�9�6�R�n�q��|]��IJ4�v�vC�A���[V痱�}��V�'��w��Ḇ0da��pb����KO
5QV/��b�9+�-1M���*C�׶��D����&R��n�
�E�x2�:,���$�(�Rg&\^T����#٬��
u�T��t&�[�eA���9īk��U.�Y�½�\��N#��·�{���͡_���y����w���-�����I�(���hz�a�pi���;��\ʑ�i�M�@��.F��2>�K�I��7A����۞�(-<܄��QO2�E�!�`3���E}��[�}ގ£Z���[��ɳ�z�+]|qg�Fe �z�db8�X�=�;�1!�"���0"���q8C�~��U@�7��vf�(�`z؋[M�OM��u�D:Pލ��F8)�"���	97ɢ^�
B���(�6^Qj5��Jv�w>9n �@|�c���c[��ol�����h�`�.'��5�3�S�	%)}?�5w���8�,�&�bN'@w�9�XO�%�~"���gi��չ�����W�����3�M�N8Ѩ�Dj�"%%V>�L���Pɽ��	l�4O"M��7���;�OuM�P%�R(|h�@����
լ�b�y�
����往��N�t�[��w���&"�=��s�d�X��o����z���Q����,f��@�E�����e��Kǘ�6�{�J�Pf~ط+��`���_������B��l�lp��4�u0��I�Bi6��'ȜDF��+�4��Ʊr���GjkbP�v�sn&��ފsw��r"��$_��
a"�ez(��+����<��,M2�1\����(+�+���0K]�Ϝ���%�?`8�c�}̞��g�^K1:��H�p��Bf��r�8
�J>�)�-��1���*��?�����hiv,[�<�ݗx�S#��2?���/�wT�i���a�]뤖^�}��������x�w휉���̛�.^m9i���'+�?�-{��Cس�b���3@����T	����u{�������!.���}�K�H7ݒ��f�h��GM�v�A�`ٓ��`͏l�9�8��Oa��ok�����!9��Đ�C��h��s�皧bo���B[oUE:���R/��F3��hi�~D�4�[�I��(y����M@-���}�`]���,x�q�C>���Rы�h ��N�O�O���^^:�M���qeXYg�mz'�I���#���g���?���K�8u����u�(��� �9��\4�������J	y;l��ڛre 5�����{���5$fdi+T�����Fc�@ǍV㚞�e��t�iҽ ��ѡ�y�J+==��=kH�M]g40<�����%Y��0�}M{1rI���5 ��ߖ�Km���]F�*2K�}��ݱg���F���i���F�9�m�b���E��S1�<Y�3H͠�U|\@��6��$Ӕ*h+���z1�����$h݌sv4��c�X� |��8�)�1	e�gA�H<�z���PP��X��z?�wc���Wxo��D~����_Y9�],���-v�g�� &h<���Lm��J����T1.u�[An	�w36ƪw2���^(���c��5�7�V%�7-y�py1.�vޗ��x�RRv �*7�||8�͂X���j�w�(m�@S]���ezB����݌�o�.S�������r��c���r��'C�,s�`��M��А��t|���x�θ���6b���g�Fa��(�����J&��Yق�������/SR;��ϭ��6&��0�1�I���P+�<��DӴ^�%��9\��v��7:�1����ώR6wHq��Ѻ%���-d�^9�
AM����'�c/(��bA�,� Ds�O����+�!��8!��i��z �c���Q"�z�m����qK�O'm���u��;,�L��������Gq����q���1H1���z�`�O�[{&훁U��%(l*R��,q�-<�wN����j�<��j�I��ԉ�*_5��n?�/d>mr	��GѤA<B�e�%V�9�3���� �]� ��^�p:-�����[_�ܜ��0�D��%�kSM��eA��k���fy�N��We?�E��@�\��z�l��?��~�����Pu�EL��k�H�t��#�`��j�t��c��"n���meHTG��a��9,��%��������� ��o#;�h��5^�wqE���``6|�_3�]6��0a 1�#3��K�>�{=Hsh�Hʋ�Y��v��!��T�*��e����|���w��~@�%��Z���@F:�O�R߲��1h~댚#s�w��n�I����IU\sH��~�Q���M��|������jkt;dПN��EeUI����;K>v$�D��Z�i����[���O���71J��F���T����R��tc�K���R�����Բ
�fC�)���p��U�g��:"3ةڇs�N��R���ʙI�N��%����ȁ�_P���#1f��$D�e�-�8C�(�!UF��^��&�H�^^sJoݱi�'r�'ﾀ�bq-���d9OZ�r,hUSR���JCVӜC���{�P,����>����ٚ�ؘ�t&^4ٶ�[*�fj��p�<ɹ\\�5ϋ�z�#L5O��5���׹�eS>�����̼d�f��.E|�鏟U�
V��=>�ި� ũg�����+w���̞�pLQ˨Y�_�	lʍX���1���
]�d��ޏn���a�}=�9��Y�+*�|T�PJ��2J�;s�Kͱׁ�2�N�����b�{�hD�x���Z�{)�;��]�BV<8�ip�V(~�"D|��$���N�e>����%S�,����Y� TMrr��w��Íq�K���S���ӉN��J~B�Q�Gg�4u?��c@؂�((E*�,��i�[�v[�%����0/���>% �ti�����V�$�UQ5<y���+$Ǭ�!
Â�`b�0����@���� ��`ͼ��=;�SD�A�m�;���zcd�59)���-_��F���a=ٞ���\�v	��bp��y�*�I�HA�B��鍗��D����;�#��|��~ocp�2dd��~���P�{�܇*�Y�Ty	���|)��p ,fI�
j���Cpt~��J�,���z�X!r-:�TJ��u���^� � $#��D�g3��<W�U�� ɷw�L�M[yVj!��D+�� ��A��B=���}�c�፰3Tko�2.ύn��T�
�bB?�<!<1o�H�q$���H��\��es�������4W� aΖ���ȓO�\z���ďB���!����p*���s(��/q&�%8R��˄��3�����F��=�e^+�����:��넄�d3h�՘CFF����=�͞k���n�#:�J���Β��I���0��&Ӗ���X,Hc~_�J��M��Dq � g��"��t�<d�M��&��M������U�q>��L_��$�a���搘���}��x���_���B��I�0�7��k2����+آ�%F�"L����A||�͝4���
%����S����Q���ĳ��b�^�iw�w��$'�%��s�M����/qQc����,���?ol0��H QJ���O���ݫ�|�Z$��]���ty퓤;�u�G�?@D���r2����i#�%��[�7	9w�v�^��v떸LiL��L���x%�Ģ`I��D?>�d�2�<�l�k[�Q|Q�d���|�QO��/笵s��}��L}π��9����Z<�]Ҁ��}^�9�;�.ӌ��s����Ŕ1�T����!m�o�6׾]cC��3��L{���]2�`_�v���T�&h �A[���5 �����x�Fs����`ETe�����q�̆]5�1cv&�C��h��[����İ)}�A�fE��/H=�v�;�q��&����mtu��`�#�4!���a;'��0>��N�� ;�j#�L$0��Bwo47Q���I8U%V��ƙ�u��6��/]�7�*+����6�0���=Gջ+������ �x_�=�n_�ꄖ8�A�!��ܞ�M[�K=��o�?j�T��T֪�H3���
,��^Z1�T����3!Ǝ�MqTqz�E�G˼���G�p�N0pi4n��ZD�('�z�8���=t}E��y�Q![Q���Ȭ��F0���Z��2�������}^%i�1��?�o�BC$׹6~uf+-�4�#�ۄ���"���U�ٶ٪�Z����a����"�VY1�gv��S��,]*�ª�\VyIj������*�'t�L�O
�����yl�מ ����$kGe����O�{2�
[%�Bꂔ�+�}���R�%`����5��L�̀��VEt�ޘS�Mo�D,Do�6�x��&�i~׹-L >Qe��t���pr_�7�YѰ��ziy9�3�KxDy���K�LE�ֿ��66��F�U��V�WSB��īBMҔ�w+�ԋ8%����G��E�+�撨�Ρ��T����dmK}�C�y�M�*�f�J�v�H�����m���j�$ڸ���)���>��Ƒ5���{r�mHg
�z-�΁��iy�K|@�>c�"�cj�m�3h-�$�h}���f�W(���Zi�o��W�e�E{�'��Q(��	��CE�4��*��:[Zˮ���,x�J�I>lO8��v0���jx�Gm֝�Ae���)q2N�/�T��wUct�)�̼3ȱ@Lq����!�R1��3!N2M`,�އ$cv�ʃ�q|�-�f>Wc��]o�R`7�9sg��Ee�γ�n�f�ɂ>X�!�&�0i����`�p��K��@?7іp�7%�39RP�~��hF:�&�0�g
�_^!0.A�ʽ��]>}&>��S
T"���<w��~�U�@?D͕a"]��@�s�`% ��1�+������`Ї�G18����,��^>��2��lt�yN�X���ɋ��N�T�=Z�̱��#ʊء��nֵ�@B= ����i����<�HD�9*�coT�_�>����r���q�m��f]�NzJ߁��(�a.��g���65N���t��M^��ђ$��!��>�K!$RK���x;4�1��Td�r�;/����{l�5F#)�j���˪�A�勻$<���f�V���{[L�e��r��{���A���8��6�!�Z��WT~]ߛ���L�����DS�D 
��o�f�Bؑ�oծcZ��B�Z>(�ʁ�5�d�;�q�E�+&o�tX�G%�ɦ�أǆ��)_�ŭ���3��5ӛh�T��A�JT�eIl�2���>B�S����+ɻ�A�k���׷�h��o�H��b���Ӏ^�m&�^��8H���@�,���5t� ��!�A�Ȗ�����0�J����[tz�c�%ݷ�<�S>f�dd����ׂ&����nl�Q�'�3�a��6",�Nn�Dk�O�$d�?�5N������-z�R���+���^_�R����6��SX���*5�wME�ƥg�Sı�Ӫ|.)/�*&+B��o��m���sq�S`��7������v7���1�]��\�..BǦ/��vŜO��� �	%��*�X���7�?��c�i=
�ʎ�Q�V�ݿ�z�/�1,r�ɽ�
��67&��)Q�%TB�`�9��ٟE��`��T��1�2 <��2wm������R!J�-�_�I�)[q����m��� ��#��>���@g&.���T�l��V,�7k2�֠Q���q���w���a�F���*nkjג��+�/-VU�H�d��P� ֡7L.U��d|yX��z&\ֺґ�Y�T$�0p`�9Vlz��/��O# n��63���*�9��k��-������t���I3�8��S��S˼�oof��R�X���LY��c�)S�4�׵AR,��g�
O�o}�J�^p��ۃ#ϋ�$|Ko�`gV���4��C�S���wRێ%U����W���p'��m�C�q����X�9G�Β�}�l�o���,圇����BF��#@�d
�T\Z�vM�,_����`BA��x�{�%?�/0K�[���sc���S~\�������ͩK�ɶM`�cPD�ZN��ٔ�j}�ܴ&H�'�K+�U[��ҙn9Y�$ߪ ��_����V�0�d9e����|��"�����
rV�r�S�<�L���C�_�'J�?�\�"3Y0��~în*4hW�"T�镻.|��l�M�J��#���#	�'��dQ�B�yK����� F�n f�@�[X��c�Y�W�\�эw����w���"�7iH��_8�r�[ɑ��8�Gб�Z���\(�S�,36��>[��w/��i�s���e�e0Y(>'�zQBi��1�����/=�U�.�̃�61����b�2WO#�uy��yJ4;0�`�-��N�S�&�������2OM0X�3�`2Ԛ�Gs�z%����_��' ��%|n�AS�A�-�L� {�PR���x�%�cGG��"�����lބd�����LΙ��WK���.P�%U�)]Z�7TV[4�v�_�E��$5n`�sJ><�f�>7���h��4�3�y�
Ƀ6��b�U�ޞ�G��q��k�zI.2g~4���0�nC��	�f��D�P*WH���sY#3��*��