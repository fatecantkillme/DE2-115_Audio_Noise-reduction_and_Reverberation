��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|p�n�U�_�e أ�w�T�)Ѡ$M��_�ES�3�� �����æ��c�5c��cc��N5��d��L\�b���{
��v�0	�ݫ�*��HgZ���B޿B��������X*�;3����Tsʠ���`�ߞ)X��vJb����x��ؽ�Fz�OTB{�ѻnRd���z��4��rg�6�������,7i�Ab��_S1��r�?Q��ز�>��ю��[��/�R����`�像�Iߊ����I�2�,��3yU�p�U�b��%[��`M����cH�Ecf9#J��ҎZ�X��ݟ�L� �}�=�`��&q׏=�>�MJ�4����I�o.^;z2����E&'��!3�~B��$�z�[_�FyF�:`Nec��S��c���t@WN� 0�*T@���G����󌮉J���/ʹ�'�¯jL��l%f�Pd���DJƣ�~R��\l/���e95��ݔצZ9֮��}d,�=�M���lM�^��r6h{_ؽb)pHK��P�Mh���È����j�L�}�ލ�5!�I��F��D|j�.$����D ?Ֆ�J�--���J�VP�j�	Jxg?S��'�;��Q�q�-����� ��
@����:�[F[�c�(�zy�Y��֓y��[�	�|���K2s�cwXeq{�*�?�W|�s*�I��py�N?H�Q��ii�9��$���^J�zd�'`a~���x+�\��\��MX.��9.x!?�pB_�oȼ(�\���Ɉ�����{nB��H"aZ�b@G=Ô���t���^�y%�6�쓢�.:
Ho ����sbܔ�0yh@Bj�����W:��+Q���&]��!y.�j4��q[��Z� #>�1c��, Z�ވmD~CIZ0ώ�$D&@�k@0�0��U:�����d]��v� �*�Mr��)7�m;����M�X��taԞgpO��;g�5Av�e�ܪ��P�!o�����7q_j ��*��}6�?�x�J���Я���E ��ɎN�HQ�JlRaJ4{�Ž�z�c?�hl8��2!m�O"��|cO�>��@�m@��Bl��_��a�>���	$:D�c��^�:�@,?��cg��y4$i�a�0Fg���E��J�X��ma�w��ܭ���[w�x/9�G׹S��a��T�v�e��ղ���\"x=t>w�VF'��R�OeKhs�?N��4�0����l|� q��R��I���3�~~�I>��A�<���ͽϧ��I5�گM��T���w��a*v� >�.��DȌ�l�P��|}��x4Ũ��L�l�1E��
��az0�&�pD؄�m8�с���W��j,���$<�ݝZ�����(E�f���.X��M����Rm���Я�ܠq\��m���K�%�Ē�dӝ��k`֔s�b<�K��{=}�Cƞ�l���)=��կr���o>��L�{�����J���b��ِ�1�v �����"˂�)daG45z'�%�����'o�%��Y[��J�=}T��ݧ�_�P�P��j��*x���Sv�����#���Tj(�B�yN��d�0w1���ag����x$�H�P��ʔ��ڙ���t����Ƽ�<P��,c�jL7pTم|!�[a��t("f��K`��8`)n0.�AΥ��?y����r�������CH��o�OܾNkV�#����U��~Pu�HI�
�!��6�&�A`Zva�WTjO��(��%1o|QҾG
�Pq4$�CKf�X'����˛p��'.\9Tٷ��0Ŝ��֘(\Rv}�y�t��k�
^`��4�w��"�e����x@ׯ`*�v��t��³�ua���^���e����^!�;�r٘SY>F#!6Ԥ��أr��"r^�5]v��S��B�s�^@6�w���!�4�a�S�mBc����J�R��
��͐�)�b��O��O��� �����-"}�g�#�^8Yp���*��hi�|%9� �zRN�<:�z]y��.��L��=z*����o�TP[�ll�\<�,X4>�j2��'C�À픣 qsFڗ��2�$���H�ҾP6$ʋ�5�wQ?^�Y��v���T֝�.���XN���G&��5Q?�1��!��y�^�8��~C����}D��[m�a��S���I�U\�EKN"��6E�񶹽�.4�>�"Y��
f@��xˌ�B��m]B\����R�)��U���W?�k���A5�{we1�],�c(Q�������@��%3�4�"����Jݥ�uH���DVx�!�(�KuCr�N8z¶�q��Gr��"$K�ehSj�L�\��g�ZPFU��Ύ�>;���kwt�:�fb���Rgs���WB
V��'�8Gy�j)&���se��5��]�8g<��7v���n:��w���T����JR��W���F<��d��
z20)���5d� be��q�%������ߙ�v��)N��(��U�:?*��UmV��?�7B��ģN�܆��<a[���">�٦�N/WǺNn�֡h
9���X��w���5�M���M PP�x��y�M��]}�y���-�q��$�YM���Ϗ���
�V�����g"+b�0%�I��C"pH/c���M�Ч������6���$�Q]p{��#��o	���J�[!�h����4O�����[��"��f�}Ks��P���m�;��$[_�2��V������F�ߥ�]��z��R����+X�����'����
���һ�2�k������@�]�/t�\]���a��y�@�`�[�f�N��:WWL.��%}+K�Wƅ7��J�d@����<�ɍ�6c�O��?��"@�K��_��ب�UXvu�2�z|�)\�ܙ���0l��?�ܹ��l{c��-%�S�J��R���O������mZ���H������7/��UQ�$V!�������P�/�rс��,�
����q���(��3 ��3?��<P���6+���sbT�b���x��6.�	4i�� g�h���6_�i�]e$+�t�yՄ"DavW��.�~��ȩ'�x����Ż�u Zo�
���7zq+�Ϣ��I�l�7��U��&�����y�|��)m�q]�!`'_��ʒ����Esȴo	�}���~�vVHc�x����M��q�xj��S�^�]" #�,�%)Y���������S���LK_����m�eT<�C2� ��{�]GW��(ۃU���P5RG	yO�R�TM�Arpd+�#,J!�+"�V�˰X�����*��[��#�#0lR�(C���֍��O��һ�q�.�?�9E���������T>�����z�'�}8bk��r�m6>���-&A���j�fZ��~�N/��T1ϥ.��O�9��O�����n�F���a�k�����j"v�S"�hH+fec��d¬��:%&��)ڱ$�P)������İ���E��pc����?� �GpG�|�>ba6�n��_����Ol��kV�{ٸZ	c���$��I4�}U�E�xBi��L�YF�(+���ϸ2h��գ]�:�F�}��+����=�����)w���4�Ulz�P��b��,q�w���G����Z�-��w���-�at����+ݲ~<\��պX�+vqS��ݻa_߭-���3`����4F�=
t������Uˁk�����v?	>xԥ��r�%%�X��s�� k>|�BED�P����>�J�$S������!��79�0C�I:8�mk/	�� ����� �[���;�)���9�ݓU��!��=�D�+�!�T:ɒ��j5�]�J���ׅ۽&U�]9�Pj����`MJ�9|�*�<"sZR��o�we):��CRFH���������\�cy���0��憎gl�'I�=��EK��N�GE|ƭ�t5��My仌��Ü�oŀ�.ԘĂ��2}��x�w���$��דXE����!?iV�kM�E�r�[��{�qI؎�u���-�)3�����I0�>ݏ
F3ݝS��Y�����p�C�*,�(MY�QE��+���<�.=���̬8��.ZV��Z��K0y�G�}���	ij<���$���w�R.j�����[1
�۷&�ɧ�/�kH��ہ�}\������A���r��L��R*�/�ˡc��&�2�\���Mk5��Y�C[=aj�4��2}�>_������Ʊ��e��f��HW�S�h�g���dϥ�/�+N���i�|���fI,�E��wFٜ�H.;@$F�!�/D�t,]��x(���!���� 5�|
 �C]m��(l�-6/�T�x������ =-~̔^W�w��5yF�ݣ����YkN�,�V�HI���/��*�>A�����LP�l_�.:���#<)b���7G��%�:"���^�D.��)��i�S�䊇Š�E|�*�X1*ѥR��@����Y�=��
�^_���u�f��Ä��d���0�ݞ�{[�bv� ��>FG�0��]�UGHb^���A۳�iG��.<��-�g7��dt<n`��O���'��Z�@[��l�]��i۬����I�� �2=�.@��՞G�<Fs� �O�������-�\,@rϽ��^8�����,�>P�g�$��u)j��T2��@Ug��j�<%�5pn@��f�iv�z@��c�gV�3�6 P\��Hr��t�E��=W��?�R���!����bm}6]>�N��}�V�' 9ӠJ$���e��q|�J�y�7˅d[��.2ǆD ���칓t���V׏��'���^���Ɋ�H�vp�\�F>&�����1~��泪�G�im��Y�w/�s3�����[~k�+�;�w�I��t$�J���mgr�tc,�c���PRx]60v�����=�m�~��?���������\g��|�\F�_`��5t�wжO�qHj�pA�y�����	���qZ#=�+;=;	]�M�ފ���$0W��}����k�5�OU+�<B�zN��!M	"�0W���*1��A"����c���<�h/ׇ�|_ s�����u[�B��k�N(e��wus�td��m�L_J&h:]�4�0[^b����pg�6��c�+��G�Y�s�2�7���=�����{ޥq��Y��C�#�F}r�2�ƺYXA��ǆ����e�ֳK<�￧�qy�l�|�)2,�!3�Mq�M.�q��a�(�F���^���j ����Xh&I�T�����_xM����H�Auj(�O�}܍������!t)�w�2�W��>z Pd;Ie�=�e3������~}*�2p�i�O�M�*(�`a+]��I�r��&Q?&�Haܨ"K��ڮ��5-HA�E�#�{�iv�A~d0�9H�ޭ���2i�W+8a�b����v
���$}(�;�/��kS�'\�{ms��d"�isg�O+�9��I��]w��Ԟ�?ɤ�à�)5��6��լ��O��!<,�B�ӫ��0�4��9V�����\ͩ���Rw��u�rg6N��p�ȅL�h�sm4��/�J�/=��4'��~;���R�xP��ڡy*�I��׀�:����x/�S���bS�������7�Ty�`R��U¤�%BA�;Dg�gCl��M�KT�=l|97!&��������2����أ��X�k���\��'�gј'�&�lc��~�3�5� [�O�#�.u��V��C�a�n�f(�<�1l���.$0�N#A����@7��_�r~1���d��SnD*9I��ߪ� �I
�V�1���g� tBQ����I��XT�w�E�I�����kg,ǂ���+�BA�GH�&���twTR�r^W��w�?_u>��Q�	�
�zS4XF�݄������Z��;c�E��A槳W���D&�e�񋶺�xPN���W�֦Ae$㉝��źG�M�p�Q���86=�k
a��-[�s��A�PxK~�e�zj��,f8% g��v'i@��Ruʼ��i �J�4�����ur+��Hb�-ȑ��|Q�K�7i�Uf*���j�#$�fw�Fa�vk^b��x'c�1�L4i�굹#{;��_�(�-z�ժk4칯����{�ƢE2��ķ�AX7�/V����N�P�2p�ߊ2�?��M>C#I�뿌�Em����
�Cp"�-q��رOiS,���%�q8%�E@�������g���Az�nVw�����ݛ**����Òs*���,�{d�ũ0�����0������*�~c��X�=�����;��Z٢&�O��dY�v� +���z��.�LmM@uy��7�$T�%��hm-=Hy6�C�B�D��p��30r�6���<��W��5fp�+]|0&�q�M�z���ё؜��~��a,�%�N�<���/�"���ǳ��!t]�w��8Nf��A)3����v21H1(���;����ڀ�n>��!�WgJ�A�4��Q�N��~��LV�R��3ru2�2�J"Y�*��L,8t!n�ȱ�H��n�����B�4�E%�����V��ͭeh+�!�>��X*��ɛ���	�Уr��:�]7��s;eS�\֠_�9�$���Qc���ar�u��1�^[66��֟��!�8���b�'��/W�RjV�o#\�OJ:<&NH�����ƥ���P+����h�EBҰX����g=�>CO�h{{wm�Ed$�m�Źq�=�t��'kY4L>��yeWvn)��ku�amJs����S�#!ڞ��~��a��!�	��݃I�UPH#�&�ZI�v�u�#Կ�-��Sb�4G�C*sܐ�R;�r=|��/JtK��f��a�R���g0���l��dje��t�4�ŒH�+��L����zy�tp&ðl:<��þ���70*�dP�fBBhq��:���3_����6r6���k8��-Ю�dϜS��|8#o}$x�@���9�۸U�+!�Ě0Q:�[,�낀h����`�K��,<���M��8Idq�Ah"*5-V��No|6d�Ӟ�BQK�ԏ�[;���+��:s����	���^ W�?\�<�
��F���@R����B��i�6 @��^ߤY�V(��2�����tdB�y_�4'�򛟅>cg͔5!��=��k���Ml����=�w�,se}�N��5��w?�6Z)W>ܷ��Qwd�ƛn��Σ���A����]���@�n��
!�'�3s>))�q��ȱ����%�$[@b�o��=�ٱ
�nu3$�"0���!ٌ���{j�ޠTY ��PP�����`�_\����Lf�i�1��%"���iG���a�_���}RZ=0}�k��~�=�8'|��NDK��	��h'&M��zL���DO��%�Ѿ����ۖ#�Z��\���EC���L��Hf�̒�	�Cn.0@5t~�O�nk���`!j� %�׺��Q�֑�)�'&9����ń��(Ze�F�^����@O�Li`ڷ��۷9�LƝeϒB�G:R��kɩo����i�?<5����(��\����i�W�	Q~���^���'�|�ZH���m��qO�/�Ã��~#e��eYQ�k��
�?����#�r����;��	��_(�|)'�
˿��v.�#RM�loq�������zjټ�!�_@����������r�ǅ&��!-��*۽.!��A�g3������%��9I�����
1��6���-z�s��\i2x?W�
���oY���'���������?��")�z `A��n����
^ʴ�-�,�(�P�,К���~́�+ԶH��������_���7"5����q���ϯ�̉ދ5��Vu���6�l	��4�:�,hl)_��EwQpo��Xl
��������2h���R̝�|�s��B�&�ե'8?lB�ɠ(`�*ʔ��C��}�m�����g�St�p���[�y���HW�o�m��J*��{	8l�⥱�a�\z��n$�{%Z�k�j��@ˌ���?�&�MU9=����KT�di�+��?3�[�r/AK�st�F3S�׷�N2�gt �<����y~lD� ڤ�����\0E�L�l�%y���8�����A�q���[{$Uh�kR���*��R0�����Jl��9T5��!�=^aHc��y�OV�_Л��p�m�A��B$����EwRb��p�'3;Z7n��?��ګ��OHUX�a��5$����}��Ҭo��<	,� P�����^�g�cw({hNΘ�N�{zX��7n�-���k�Vk��+^�ZI����;UѼ��u��5��r�S+q?�^aˈ�T�d��9��t�(t�$�ϝ��������Z�����n�^�x�k��]�;'�r)oF�'�JO�Q�Y�%��������N��N�{*���d�1;�y���z<��1~ܹG��� ����ü;��~k��ښ�'�C���h������5��&|���׊'oō�pN�3�ĳ�s}hV�$b�����d{��j�sP����tYW�p:�Y��C�;�W���aQk���"�{�fֵ�~�i���(��笣3�������j�/��s{���^O����"�n�hz��������7x�2�7ks��҇^� ��e��Ǉ1�y�Da�5�+�KR�V5v)�+}��!N�[l[3�U!�k ����ꅼ�jbd3+M�@���`��'}�K���m9�ǖ�O]�����;�+���3�;��{E�i��w(k݌��s~��6����I���@O��j�j5,!Fցʮ�H��IX )Z�As��J�͑�Gb��������)��U��R�{$˂�
ct�2�"b4�|qI����0�	%e�˩gl����_8h�LO�ψŏpy���B'ԇO�FwiH!R���"^+G'�K�)G��/��]V L-Yˀ��tV;�x��+n��Pǘjlw�N��?������;*n1k�X�S�+xO[�4�~ω|7�?�NQy���p�E]�vf��K�T]�Ff>X}����_�ec�`/��Ifuvy4���l���R]���%�Q��.�I���r�Y>���K'���3��P@�������|���.u��0>8
�2���h���[��C*t������v�[��}=R���')��Q��>L�A5ʵ�EPte ����P{�˃�O���U���Q�O�ޗ�]����C`�1�"�Sh�\��*���5����$!�����-�d��d �L�5䘫��ȷ����ɇ(?xY��}E��QLD*����Z/v;a%E�D���&	��i�2�J��dO����]�i9����3�گr6�[f,���k�ba�>�˔S(}|y2؇�3�C�j��Z�]�JJnO~�[���e��s�?^����;MŠ3����Y�3�5��|B�)���q�X^�.��|��J?/�CL+H�!1������׉��3e��|�G�EWXL�ԡ�a}6�󘓞l ZUl[ ��b��aԜ6�VTP@������ePu��i���Ի^;n��2o$���	Kl���9h��bb=���i�Y8����<�A��G�1�µz�ڑ�4K�
�bh%G!D��RDx��}*߹=~���g�#ߡ,��}�m)o�ߙW*�k�ko����+��C�Q�N��D����Hm���z�l{6�#��$p�2��Ԛ�� �O
E��y�b1	R峒B��(h�6]uk���kZ�q�ϊ��=^鐷o�GD*�ƚ�?m ��9(����f������R�s)�6�S�Py�ΐGP�'� ݧ�_ ;��p���6w�\�d��>Z��"�|�Ԭy�ߴ�^;�`��{|F���L�$Nђʽ�Kc����%]�6�G�Z��S���՗��F��<ɾ�0H����ct�f)*��#�E��wq�	-�uXa�=��0k	�����b
:n�c,�X�)��ԡ�8�����J�����))_;\.)b�������ꇥ��RM�/62?ոx.x2=C?��ا��ζ���/��Y�r�����$wt����h >�e�#�[��r�vȠ���SQ�P�Z�4�ҏc�h��$��NKi�Wgy�[6�i�iBY/Ykʔ3;�c���\w��3�qr��Z���œt�M�!���v!�0 aN���xH��HR��$���$�?��}(3Cm���薽�d���"
8�eM��5z�S�V<��`�I�)�o0����JUU���2��`�(#�Dvwa��uM���,����\{@�9On(�g���F�&���}�@�q� |;����H��R�䌥W`)Rw��G+ǃ}:c*�WZ
��o/��.��5	s�/c��f4��v�lR��B$�Ɲi��k��"J3n:�$ދ�a����\�q���{�&�(�*B	)-��YeT��r���n��D���3�>�ѻ��@��e錝�`��if�N�X�����;����s��$�>�]�"�zʹ��}�D�;����8Ck��i��\ �\���x.�
�*H�[��i@�y���_�]5���m
.E�v�K�
�WLJ�AE�����.'�̰2�@�\����m�.�XIJ\jGk��>t&O��7ݪ]������hS���g��`��S0j�kzީV�<�(��4*�'cO]7����9��C'��ư*�NGY�@���$T�@>L�ʞ@i6��@��;"�	a1�����y�c]4�_���ž�6�Ns]K�Ʃ�#~�v�9�E~K�����Cd��ᔴ��UK�<W����D�6�eU6��=�"%v�[A�����_:���R �{�3��r����^��ـ��V���.f!�,2�FwkB�8��[�2�ŭ��X�r}��'<dd-�Uk�m�B0�+d��-��A�:��.|�i`��?����9=3 1f�b浲�3Aj�2�w����?�����:��Hc#z��|��iI�����4�����a�_]b�ޘ��M{�t�-E1�%�>�v���*L�Q�ix0��<-��M�=5���#^���TK�7��)��j��$pj>]� (��Ox���i +T��:���ǳ-=�09�j<���#OT�&מ�l�!���ϫ���!WJHa�z� ��F~��!�Ssn:�9���]��bf�g�6Rl�u�#�����^�i���4��͡�������<92��Z����b�B�:~�sa�\��{��j,�S%�$7Mda�BS$Tg�b�$�q��4��'��B���������@Dqb�*~�\��B��Zj�&��|l���ys�����xO�>�^(�7�,E����eB�ʟ���w&�#�e������W�����|���ʦg��j��Dѷ��E�_C�g<l-�gF~�a�~`4j���	�:�������@��&�QIjߨ���6�+J�zs���j\�@��O$��@eMk��w3�Oc����*J�������4������^+�-�SAUB&9���Di
�k�!<��;l���'텇�폗���X�!��JU�����%��(t-�9S�"�XlĈ#�66}��;sC�k�2XW�ȉb�v>E <I�s��*���ė�Ҭd�Ա�O,_W���e׵a��3Y/v�O�
�3��c�'��!n�y�0\ye��*"
������td.��I�v�a�����A�P�SA������7A���I�k�?��2�q�n��C��-5���U!��d<b_�ִ���#ieN�]�>�F��0*�=ڹ�Q��eܶ���|>?�"%������]L���.�2"�ػ�n��g���#����-��� �u�8��ݓU��v13W���I�줫^:e*r����ٳ�@^V�Y0[�¢搛ޮR6J�r7��T�ڏ�G�4��x�)g�,7��] c����.��\�=$�L�H�I��7�.��7������%��Qi;|g�^�<�d��2����'�|I
J�w����l�C��T����N��V�TL}pS"ݻ��X�� T6��D
\j�.U��;�|�^"'!������G�Ŭ�'��J*�m�֬f�V�9���	�x��ۆ�ma��TR�B�Ü{�G���-s0_�|ڦ�<#2A�1�8��(X�Og⃎���1�D%�x�䴎�\����I�cK�
�d�7�OM#�GS�@>rK�Z:�h̒�/26�h�ƿ�iU�J�)�Ѿ�+5,��i��f�����~���Ӯ
���ƴ'$��m#��3;J'�l����b���g��X����u�|Ҵb9.c��71�^���5ᑓ��T�1����Y�yBB�N�K�~TÅO���f��u�-���hf=dj�5�Y��>L�������ضL�Q�l|���;���`��sS��+p-�]�%Pk���vYx��B���lx}���_F����G��'��3����ϔ�sdg��-/�N���/e#���b�����5���S/�r��8���G���W��_��V�a�O� n�!,JMQ��|�O��'�;6�YZn�1%�>��G��H[�*�Ѭ��{����?�@���m�g�a�|�h�Af��9Oʼ�n�`B�!OW[���}�`D��_/۽��;����U���>���}I�f������G �D����U{�{A��� #I���������ݴ��UȦ�{X���B�mKr���U�X��6���?Pi{�r뷙ƿP��N6A�w���qC���� �N��2hM"_��$�$�Q�$��׵�q� \�ePa������lLAv�D��`a?���B���\3��Mg'9����0ƕ���4��F�J��4{J����2�-Ix�!�#��:o�~�@tJ{��T��������ίm}���P/�)ȓs?[��.K�
�����2�N����a����4�\N)՛C
p��E�X��=y'�װ���N{+aNg�z��ɰ�}�>,ǩO�L#�r+K.���+����&�o�%�\�D�򌺟��a�����*UBL�$��h��%�6XL_vV*����x
���E��ОjV���u(�h���VE�
�����ά�}w��Z�pM�+�t�����,�3�I7J3C���ShÆu..wu�5�UO���N�=HꆋaW�_V�L�g*Ѳs��%��f̄x9��l=,~�`�r Ǒn�ɋ*�%o/�x���Y���Ҷ�L/?��r�9
jz)��[���f��R�����(�g_R?8�`�2B����O����2_����ָ�,2� ������݊�	n(�����#�+��A�RK�	u�gju�溺��#�a$�G򩿿�K<m�:���b�,'����W�A�J2G1IH�Փ�BG���N ����ڊq��U��&>w��6��k�ʆ�K��f�x���{����_t�9��@b��C?h�Ǌ�+FJ�7�
��ݸ�@���D�.�n[�Ġ��z��t#��8�r 2Cy<���Y����_��M9�w����c;�G�i9;�b�ۿh(�	�줼��N8O/��}�%Df���"��@��g곪�)���+��ЧK�q/+�� ��K6�N���� �f�S�f-��t�T� kgZ�i� �%^����}y����Ey~F׃�c�z�N�\��}��O��^��Y�R�2m:	��e?1�ޱ;�^(�����F�����*6d�M~��sF�<M픜0���"��T�1��*��Go�!�����W5Q'c�C8l�Doi�d��1=��QD���{��+H���Ib��Fϝ\!�
��I�A�x[����&��I<_X���<�ti�cp",�Z�X��wWA��8\\--�2����kv��qʇ��"wm/��8��X�.>���SQl���S���kp[�DIr�x�a<�Ө#n&��_YЕ���^�������\���uO����6��Rr ��aJZ1�|�4�1?ؼLz�9Kc3�e�¤y��A�7���G����8,
�1s��!�t�p=q�p'=%n���#�A��G���}�|'�ƪ�f���,�:̙f������J,�g?{86/���2<3�*���(P��(
����Nݎd%`�� $	s��&�\�]�����V���kzasV���/���@�	�����I���s��]��2��m�b�߂Řzr�A��od+�'0�%HcB�+Q:����|ܺ�K���h߄9}�T�y�$b�{�e)2��5��,��^Z����B�0|�J��.��`����6�.��;ֵ��q�����g��R�gLlB�Vv;���a��3������,����o%���W򤿠��@4��9��̾m��d�l�NJ4w��@��kC�)����x�|4転� ���4�w�p�`ɴ脖/#M���A��+Y��E�f����}~'�q֥�V�ұ��,���3�P���,��\`�(Y�&�g�c�~r�u;Ja�zꖶ��a�3�T��P4�V��fc�X=�)�HTp�<�d�6B��6�X����a�$�Y��&k�MV���<V
]u�ˇT?"ـ(DڰbP�y�,>���_=� �F�BZ�\��c ]�A��<������O
D�$D��]Jkn��`�&��cgJ��N����3��*�{[��xbAQD����� � kp����~��7��s����o�A!j4g+"P�^�����E�T�d	>m��h���4�� -t�ԙ�c�&���r�d�F����F�>qb�[�t޳b}�5G�8��߿��i^́�sX�s'�QcP�������eؓG6�B5��1@A��s3^�38.U���x���=Yÿ��(�,�	��6�M�~`��\�"B��LE@;`[��cYM=����5j���ߔO��1ڿ!���T������4������D2�I�!F� x�����X�±��Hf� ��6�J�C��u$���
K"'�r��-N����P6�iZF�w�\RX���m���0O���r#��3Yqv P]�u��P�N4��ss���W]��fX� �ܩE7q/��������'�c�b����yߋ�
7z��$}�Z�.�C++����di������:P�����$�	��+E=�YF;�e\�ٱ�"4jBR��$+��9����!%��U���j��R9��7;���;�C5�3"q��?ǬC[�>��G� �j9H���O&4���?�O�|���PO�xkb�	Qa���%��>%�i�T=�8(hA$eQ�zۢ���d�n7�"|�"	6ή4S7+�����(l����U7`0D�vo���z�0�Iq�0+�dO�n�� �%��*�<�
��W�ง�_�sE�<c���F��7��
{NP�in>�@�!S�Bu.gR�,eQ��kKz�aC��n�N~Ɖ�}=��Z$���	���X���N�%�w�*%��0��.��>��iC���١Vp��QШ�,v6^����9�C�	�('���kk�94tMF3�$�>�12M�L��+9L��*�J�l�3h'�| �4�m��-@��t05�ѬU���ʓ������Le�pH�8ɹe"8�+��)prP�b��T�]���P���iF��"�܇������[���aD(z)+~"���n`[�1��g�8*��*�_?��-���g��~Rof�髓�0�q73C�\%'M���Q3��N��QO�{�A����A[*:�ɁϨD5��ɣ.�?�W�F��4�.����Q�اQ�@ŌL��ѝԁ��^yR��q�����5�kh��񖴫qu���"�'��ϧ̵ '�T�Ήc�M��\���Ȱ�I��zFl��%� (�����>�htW�.8��5co=OV	M���s�9����{��`!���2��QR��W�5����/혣����P�DPA�?"�7�b�����Jn y���O���;�+d����J@`s!��㱓��t�g���Mn��Z���3���?ņ]62zj�)�[	y�!s�,d���tqyg���0���Q�I�i���.tx%]:�߷�����)Ǵ���:�(�u09���6�O��ae�v�C�{6jE���f��\�O�]�Jy�ސ��ʶ	�j��� E�l�����x��5;�*-K������`޲l��:l_����h���=�|�is)�7<�`��Z��iWU��"��7�d�����V�[��q���xۉ[��( ���!pm��Gq����8U�]�S�UfI�4� �= ��ϸ��2�uLp�Ίm?��IA����������{ǈ��~\�RO��^����^�P�`��=�96>0�Tr.+\��*����B�sO*W�b�9�|o���4�j{���Qa ��	�������b��;�1��F��ӛP��[/=q����G�wԣdS��~N`vwɔꁾ���'���%yB@m �_}�h�52�h(�Z+���oLts��k�*VG�Ť��]e���8��:����L���Ղ�(V�$~�Zz�NֹP_���aE���H�)�z�Ũ�ߣP���4Q��︊�N��"
�2�����ҶH�2bCᭊ����:���X�-��A����y/2��҃u(�ā��k�M ɰ�z�!|Z��Wt���P�Iz��0�b`T���{�*�L���ڵ������rk�m��(x���n����)+�e"&�Eh��~Jym�q�5a5�*�h���'Ï9�Y����)<������|�	�x�|^hj� �r��sBq�������t�a� @��Y���E���9E�z��Q<��k��1����J�P/@9��Cy.�<xG����?��??F�<g=×����7�����}�fZ�k.�=�S���[`����љ�)�@RQD����j���E�={c�NQ�� ���s��aT\�b�����7��
r�����
@1��sXљى�&��x��2hQ~�6�1�h#�N�	Y��L�!S��04�
x�7ȅ�𣔌�,�?>�U*y-"����sou��h'�Z��1�S�G�`��9��f	���b=#�7^�-鹱ï�p�� �$�c�+h;���<�{�H�m��ӫ@��-����~��(e�q+���#`�c3�����81���R$�� 3�-7dx^̋�꟤���V�S��O�t�!�������N\|�pK��&��d��T<�$�<�~�ҵk��L��� �^��I�BRYG���5A^�jWRU(������K C�$Fp�j+��������>$XMnrf�,/��T�4�_�8mLQ"���J��9�t3"��a��*Ō���"�Ckӻ��S�q�o{���l���D�����2|HR��ƪ�nZ"�&��������sLo�M�0�H��>���*TVl���`E!p_��J�Αn3+���³"����/Y�\X��1Rn�U�h;7�=Lf-՜](����5g��_V+:�IYk<h3�I��En�\�vp�v�#$;I?�[��$�KȢ<�T�ܚ�Ux�	z�KK�~��y����$?�]�s\w�HѪ���˟_ީ���7�S�.%�?=���s�0��~l���m~hܞ�8˄A����v���%���[�8\�5ٻL�oJ"����??R�L���r��]��ؙ�T=�$������\G�� ���^r�ipz��&Ь2_�����t޸)hO0�5�Y{�Ш���X�d�ʐ���bh����N������'����V�(���E���I��q�=��'����1f�E�$7$�2����JI��cX��,�|�h����&��1�f�D�i̳A�2�ɀ�%h�<^��<[�.�l�/�>x�hL��0�[��[�$�7�W�.��s��qyq{�	 ��h�?kP�U��*/cn|�ǡ9��OKl�{�?g�@jp~�l�TO:a���w����x�6ؕ�Ue>�:UC>7���:C��Q�ö.�#�n}��>g],�j[�I�{̺&�HF�6�����4Ė}D�!��]+��A�!&y�餄�Hv��j��>�m�q�P[���(�@�=��׳]m_�� �(g��Fr��"���Qr'�e����gg���/�,.��>+7�X���.��V]�	�s�w��c#$�����?]ΩG7W�p"{^�ԅL����UJtX�yn��Kd��Q�	�]����p�*R����u��H-�����,i���G�F�uI�
�u�6e���O��7���/��H��e��֝��z�~�������ea钓S-���O����p��?J��k��A<R����Zd"�2����0M��!�g2�S0�9�10���d:ш��"❹V�dv�KI�bj�Q!�`8X��K��ty�
��αod1x�}�{V��š�Y���p��/�{1uOT~S	�	�qb8�~zRD�������nP�>p��Ի�A��,��w1i'��'�hi�ك�a^L��*�M;~"�� �sP-���
�~
?b��|�n3��F�f���rrY�bg�õ��YC�xd���PhTJ�F��b���( ��s�a;�Z
Nߍ7�J��O�MF'��CƑG�����q�\��3_��O*c��Эln�HqJ���Q0���u�}��<mU����Ą�2Y�/�R�]� �Z*�,{�Щ�L���0�����s��:�p�I��2x�s95�P�K7'�|��VyA�U<�ԑw{��̈����E���i��iؼ0�G���3>D��g�YO�ڡ��W�����2����H�����9��s�;�?u#�PK� %�MZXC�;���V;�m�@�u�I��5S#�=���z�)Z�a��@K�R3�m����8�����&�h�*O��q��2bnG��d�Cd'��4M�?^I��g��0�Rw�hX���F��Y�����ӌT�� ���0"ia�Etd�؝�6y�֏h����,5���X�3燔�D׬5�$����O"F"�T2���H�)�ʵ���.�SΝtn.VbS$�Y�A��\�j��u���|�e%
�^vt��dy��V]+� ���]��)��&��$ �W3�0g��E��LC�ȹ�	����
�KD��
^��8`�{�R���4�H�o��~u���܌���H��zܗ�_ʎ���~��n$l\"��V��dg� ���c�e @�eQEb�:��RT0���/[���/;т�V�
Д��\4���5���	����N������Db�����S��*�l�pr��Ĥ���ڋ'm^�=۹ػذu��#�G����<q<N9%����-W<��z
.�I�Q�WR�q���U���#�1�~���rvq��8.���4Ib�,��U�i_~���
���īt����[-��G�S���* ��[�m�ٴ�����s��I�7B8�d����6�AH�Z��_�Q�Kz԰�{z�M�m	x�H-�^yA3+�g��f�C:c�՝^����[X����t��\�E�ٛô[�%�c�]I�#e�1X�<*b�g8�kqH�j��t�f�$�o�V�!��(�rIk�9ԎB���W_X
�(��}=F)�*n�)�>&��wn���9��&A<�ANz��hg"�=�7fkX��[yi����a��H�SUU��G�Ĳ�"���o��e0�ר5	D�ok�����:i~�����?���f0�;v)կh8��O���$��wж�<o��X���-N�����N��;��|�"��4��$���"+Dw3�}X�}TA�q����􆊒��'�
��[dZ���sd]K"∘\������(忩�čc�y�ŀ[P��g������\ټ��Z�����A��{��
�.����&�����I�m2��U�l�:��f²�@����q��x#I�w��`eE�ȡ�E'�bx�M/;-�,}��q\4�F�0 ^���{s�b���%�L� >�걶�c�Rn2d�f�-�%�.�t��l����V�59�.�cx�
�U�f�]h(]O����!S���M)'툭f�Oy��mSU�3B������J�8��g�͵^���-�y$8Y��b�݋���kd�ɐKO�JR1JXl���r3��py�Χz,T�3˚�}ߧCO��@%�w�h?��%�O�D7��: ]��j��a�p��'sE����N�Y!\C������*�\d:=� ���|�5�@a+���dt�1=�A��:�Ӱ�Av�mm�&??B6?��� #��������M�/ôR�e���g�L����N��s]L�:\�{�eWI�F�rܠ��4Xo���|�q��罷�߷�٦ +Y����C&��-�4�j������6���.���'|����q4����6������?��k%�	Q�f�=��?u����b!��Y��B�WRonI�P��qhD�:�	m����I���(�:?���Ѭx�;�Z�E���/�I��WB�~��N��9^��.4^�J,�=�b*���)�"`M/���������L0y~�ll:�h]��j�@�L	�ߊ��mY+#;dj D��DM'�-����HhW�F���n���= ��le��J-��-�k4�cCO�Z�F� F@j2]
�ǁomTD��}o��W�4������Qu6�c�[j�9V�.��U�i�:��s�훜�3RC$�xͺ���k�v��
�:�{67�W�i}H��O:l���O�րϗQ|R��`͒�9א��Ĕp`q�ʿ�0��:�TM�;�����3q`?�����m��*��6z!���I+g�F���v5�=Q�w��Z�Z} }�[����2	����!ҸUۈ����gL|�	��+�0����+�Г���3	��u�F!8�jVU�y�w������\�]��'���W��X�3��̀6w}19��k1`i�����c5���+ OJ���=�D��sK����X�a���n�M����צ��Nv�ኒc�0E�M��:%U�yXJ������z�T��B+�gX�ЉJ�>�R���u���̑fH�O4����j���EW���.��Kb=��|����dI��s�
>���8iq�2�h��Y���gU��ףZ@m{�DI�hD��N	aIǁ�MU$WQ����Hi����U��2��'�����b��.�b�D^�?W���>�{~>�:�!�J���`:,.xM/�-�9�V���Rx��K,��'~`E�ѝ�C���^�� WBt:����ܗ�JD�
���zY4�F�����,��U�C>�^�fe�|t��I����/
Gtn*^���� ��wL$��x�ŭ��Gq�����[`8ֳ��*{�W�D��ψ��_h�?��$)^�S�4�m�)pxJqH5&�~���ۜ��D;�C {�������~t.b�u2]H����Y%��
�˹i�L満_c�1����(q,��8c.��]�7�x=�3ƈ|
��k�����g����[��¹(�Mk�}$�����^Ǳ�zKt��װJ�nrnx�jM*�h��#��bg�{f���8F�` 6O����Qi
�M��냴ը_����l9�����ǘ#L9�-���W�����QL_u/�^C���NE�a��6�~ ��Q�x<��t����b�k$�\Ŏ�����L�X���t�V����	EC�F/�w��c�і��d5�"	�� �<����2� fȦ0��X9����{����^L�fyH1co���D+��+Ԡ��[5��	<;]��h$��*z|a/�(����_�0ܶ� �����kkg��Y��VI��^��Rg�"��x��p��P����V���\���G��U*e�BdT�"�1�@[QF��SxL��o��n�C=��ԂJ��߈��R�_��i�Z���GO�rݝ�j������)gҋcT�5�W
�D�X�:�JWQ,�O2���+ځ.�4|F���'\��Vz��yPDN�a^lvP���4�ڟ�G���`	�\�Q����:��8��k�W�������t����
;�
1*�����5���Y���$3�|Zݽ�JM�A���;V�t�ll�8��γ�	i��`��a�H��hT�#oyt�'t0�=�Ut��H�-p8��\q]�Ɲ��i�e�+�6],}���0�R��x#���Y0����T��	a�����tj�
��G�|��m��$f��u�a#��.!��H�`��p�/���R<uk��!ύG�X ۆѭ��K��-[u� 2y�^�`	�QH�o[Y��#@&����?͗�H�-�H�kr�T��Æc|e�z��%���ꏉ(&YH�.Uw@���b�����Ӻ/�
뿉�0}�&5r6n�e9�J�j�������ݕ/0�_W��K�c�xI�x����̃�j��R�-�.����ſ�J�"��.�FR��Ŧ/LQ.�մA�.�Q4�~Fv�1.����<��3�GN���-	�5}��\�a�8ϣ�h,�V��.��n��u�:�a0��y���g�^��N1�I�r��ճ@�s���K��"�Z���A�dmɤfĢ����է=d�J���$'�O/�JuN��XRdd>���{�O+®�)��ùrV|�.�t��y�L��VLX�b��h�g*WqZ�5�q��;�Z#�G�ټ}�X����f�m�\�e+���9=p�P��
Z�HR����0�X����b�zUĸž���C�_�y��C��j�Δ�1�H����x�T���@�TT�Y/���Ђ�X���6�����Z�/����%L� �;s�q�M���5�E�AFz�ɹ�L���~�>N��]��"�=�h}��ɺf����s0+��CH�?F�*^�q*7ҳ�����z�#�'��71�F:�{:϶�V_[�rҹ'��J�d�(�>��Nu}Ų=�?���i>M�^�
����H|�XL�H�B���-H6�%H���L[հ�n҄�=�r�RXy]5օ��Y}�eIN=��+6n�P�w^2�(�?���%�o�],L&���,� 4zR��(3������I�LR��$�UO�f �(7,|�����e�BT$���a/�����7��Ѓ�>�ʰ��D��Lo*�.�IX�isNg�ts�À+,�/y0�[i���X�T���0~ܶ~;�dq6���8:�Y-	�&w�B�����?�3	�j;j�+�g��ѯߜ�y�})����U-�@���Q��+�[Ղ��qt�s�D�$#g�Xµ�5V���3��7��Ag$}����|W���B��ݹ�+�C���|�nb��Z?)Ξң��g�o6*`����0�/+q��?����M��1v1z��q�6�BG�j|%'<e>�E�+��w+��4%�'0ͮ�����~�%�O�$���;c���N��j����Sm�E^ ԗ�