��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<��魁�7��V���%.��bn�֚�^\O�Q ���ԍ}��ց'������쎨gH6*ލuM��u�>k�D�WvD��eKNY4� �D=\)L�U�eA��A��z�S�h^kk�������Bu��2�5D����~|�5��n�ti79�g�J�>�)�'&������w���/Q�O�4!��p�P����I6 @�!��1��k`���Ҋ����-p�[���>�B��,w�V<�Z�x5~F_r��c���+�bl�?�뿱��S�ټ.2�EB26�\q:J�|���l��G���{C3�ѷY�k| *�H�}�i��T���v��[�����ÓK\�����C0H�I6r��ބ���P-��ضW���h/Բ�]H�J���lGD%�s�S R�:�����q₊��P䔞q��uܵM}���,p���ۧL����$�^%Yp�I7>��{Yċ�A��9m���)u�X�N'�MQW��h�䶙����"����!�{��1���(���F�O���(��Ȭ��U��A�e�i~AT�d���1��A�s$�O�L�=1�ڲ/C�!JiI�W�noK�%G����"�/v!�VLj2�V(zP܂>��Ӹ�y��{��mp����y)Ը�%b�����5�ȼ�i�)�0I���,�	M����y��f�Y-�bthZn$f�h����8m�Ë�d�A�� {��P�X��n����<�R%��W⍉�/�d��ߑ���'�=��IY�I��g:!/���fiil����qR���wA	�t7�]E	CGp�ٟ����ލ7�s:�r��o����4�s����S�+fcT-�Hm�;�
MøpK=g�$C=D�TT՛>�h�m������x��*���>� ��c���ϗ�6�CP ����yŶ���F6`�>9ǹ��W �t��8�n�e�*�^2�#�+	�01ɢ[OQ��,A>8�v�L)C�ԉ�>��2��`�9�a�1dwy-n6�VLR>�S���0b��k1��ڑa���(�L��H�c����2CAm�5�7g���j_�u_<,��1�ٓY��4q��jV��R@�^V��@��\���V�:!LhN�m�rV�
�0�_a������|���Fc��ٽ��W�eCB �C�i v\)��j�n����M��?�gɀ���}"`G��c�*~��/�_�̡�������~Y������h�4�� 1a"��7j
02��(V���\u��P�D����3�{(�6�����G;�_��5Y�:����xG��0�ն��x.����w��%����	l�z��Xb���y�͌GC�z�S�Di��u���3��k�_\-�*Πt��%��f=;μ{0�9:��!{
qW�-[����{��3�f���4�Ts���Cu�TI�W��SL"�)����ª�S�j�M+�:sA�}4�8?���
A2"��a�#�Z������}�P��WM�M���r�F��(t�>.%���
Ƽ��q