��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|�&���ڴzk^�2�\����糿|!��g���!aXZ���s����?�.����
��NT.��}	?���-�$�a�G��m���E�E71hx^���x׏D���!���N�� ����H5*_X{����e�hCD�C�1�B�@g��3��;Z�T��M�fU��S1��P�W�>���w͕|�s�y���3mAݜ�'��R�u�/��*�>3\{�۸�6W��&L_�_��Cr��!����x�X{*��c����K�b%�Ё�p��D����X1.ǂ�.�բO�hG��HV�C��>�`)��>�j�A�>��%��3�y���ֲ���܎Oe�s*�ߏڂ9��/i|!�Nsi7�Μ��Ӌ��Z��T������_�v���u���
���k�B3�]E�}���H���Mg�db続�`�������X�ci"p�#�����1DJ�3i�bz6/��˅L�ݵ���ūG'84�Y&Yv�=��_&o��"&�Q��H��݇ڸX��3=<�Y >(M��=��F��Г��K��͹jU���x�x�7�C��:P�}����賓��h���
YީF��� M����6��XD��a�B��B\j���Z�D��2�(�B| �)�qn + �n�7#T���|��;>u�"f��. gW�
�����J1��*pM4��%�ҳ���g΁��e�\��P���+k6����5׮ͿJ��gf�����5Q�a	���>:�v*^9ca��QRj��N��R�X����
z�d���[!��o�#j�4�;'�3~�?��n�$��`�"��{�7f�o�8�A���@�i��8l�hXvv$?��|�
��JĔ�`�#������|��A�8����:���kN���Tx�T?f+�h��-=��3�[ϝZYI[�C$CP��Bj��@�+/.[ ����6���1�l�	4^��*8S���!�N�'����P��vf����U���pGM2�&p��F:��A�m`
�5#�`���(��G�:�_)��S1A]�+�Dlo��J;��{�U�b��5��=;N��Í��ѹ�-U^K�uҧ����)���;�\*���OEYn*D���n^Jy���x��ݠ9RX�[Uor�W7�[�Z�f�	��n�2=z]p�w�z1�4�v������	���D�M1����,-�6@�?Hz6�7d�Jҏ6���
㽿�s�Y@��cgӓ*W�{�Ә�]2��Sr������m��Ͻ�$�p�{e������
�f���	�z�
��r������?�'5jTo�2��k��T�8�B�C��b��I,`�Sv=��gU�=Āv����K��I[�&{~����V7u��MIB�+{��@�;%�k�X"D������+�2��'�㌢{��ё6�B��u��E�ZXAo�/�=�3%����Mޫ�+�y�o9� � ;}↱\�8�C�'݄fW��$=K��̾SA�{hf������@}��ա�W	w�
�Թ�nfǄ�_���=�������gu�fZSޘ�_�q��Z+�D%��M�O��MQ�N����s��i�i@�|�[v�m��>�V�Ϝ�Ѷ���+�e�� d�K��ُ��MݔwY�d·�"ElX���<	�Z|P�f
C8�	�9��"�E	�M>8���ǣ[�4��yuޠ����P��~f5����H/$4%i���#�%���QG>�p�~�,��lvw�'p���E�e�M�����&xQ_$N3d"���.\�>��$���(�p�`�p�<�s�=�j)�>�\zu2ɦ�+V����(�F�u���W3/��"��PҨ���ىE����;�ר�!�<M�2JĞx��e��z(kHx�V+;k���§|��@�׻�L�X��U��YFVP��C����������US���;�-�!s����	B6P�����w�P.�~��M=�6����/`��\V�"��O>-��&$ᄄz��$�)�\;M�p	?�ٶ�F��		tӤX�[E�����R{�E:��E�%�:�P�������j�"���X��ׂ.�Q�z$�bv;5~��&�I/E@��T�F��j�:̐�q%%��+>���U.1FA(դ���-��Hn�L�擈WK-���<i�)x|�: z��T�b�C�Y3뢕��B�.�=�R�M�ֿ���r�Ɲm�i���`�(� D�=d�nk!0"{��|V�@"oH��������(�R�J��������'������) ���})�}��d��bӯ�M�k�>h9q$�����p��8�ꕊ�O��F�G>�$��q'|�p�,݉f��J>i�(dƥ��هL�3;�[F!8LŒ�΅`�R�?@a�zP����	c@�_��0�"N���K��y����������Ga���:&R*ȾE����E�zQ��I{>
,B,w�Ŕ(��n�N�!�X;5n�m�N8*F�-g�9� X����n�N�����wt�Q�b�ېW?p/� ���r��,(�D�L`�*�͍˗��Ũ|��_��p_�p�2�o�=���Y���~vo����_YP[4.�d�Z>�@�-�i���ni��`��5K+�Y-d+�Z���������Ո3^���ʂ���pE-A
~J&n3"�A((Jq��\o�R���fޛc2Iq�x�*�~�t�E(��`g�U�T�:��Q63�mj5�V;N�3w;|�J�-i�h�.�5���.~���r��wIG���������L� �Ġ��(�)wDd&���@��Ε5�)	��^� ����C���)N�Hcx9{�񋙰�\��G����X����N�DP0��B4*4�j���	�����Z�xW��|f���pW��޾c�FjgF>�
 �]l�I��p.�k����p�����M�/hYI0�vv浮�Yɜ;�29�1�I�kl����r������F,so?_Q�%������|�*�4�?4����ZlM�>X������}����sg9oځ^���c]$�#H?���
Abo�nYr	wL\BW�$}C� �N�(~��2;�.��,��3E1���g7:{���K�>��	�`�>�d0�-0A�1F���4�9R�x�;$^ȇx�'O(t��u"������,mWO��6!�AJ�=՛�4ie�3z;n�fN��`4���}U�tA��Iդ�g�|ծ�Ι�&aԑ����flH��y\�Ss�2R&�-����s����_Ws�'HN�"I�'eąU��.cx`��M}� �v9�Ը��|i�3|P	J�c׽�W�=)'��А�lN�wUf�c�NـJ����R��F�����<��&q��|��Ƹ�6��r.u��N8�˩�g
�ca��F��AڄH\o"aO�/�k�1��[�ϓ��~�QI�K$���d\�)vh�z�D����W��g ~C�����!lx?HxNh��o�#L�����Y2���P
4u`br�n�
s 7��kɚ^�γYt������]q�1��K�U��$i�*ޠ'\�U�A+<߰$M�h ԯ6�"2�7� <9��x��깄#��6Cj)c��"�����E`xk)k��D(�tѵ"3�4���x�wڅ�w�4�~ǩv&�����\�?�ԗ�5�����77k��x1,4��8b�秡f���+���q^�:�����	�<w�'w�*�QQs/Ó��n>B�'"��u{e_[�ՀH�R%{y$�z�j;� {c�Ő�k����8Dj�&6��6�(̉A��	���Y4� 7b4�s��ܢf�"sЕ�s�˸��]�M^f0릶���P1G������v�8�9c���O�C+8���_g}冕�Ͼm� ��Τ�'a��8:��y{�}�(E�ir8��Q_w�����T����Z/�mZ�s�.�0خ��sNg�	��uB�z\d�-�a �vx[�\.�B^F�,�Ɨ�OW���ğ�9��e0�d�<�1�_J�[�p����H|��4R)�H��4��q�n����=�dg� r�G��ٽ̈́: BNh��c�����]�&�;�>�r.y�!��]��檖`'"�9Jlw�+�6n���,��9���ܷ'ͳt1���1�	J���$�h)�.j���������)5c�PRvp
�Φ�7U̪W��[��zm5�X��y�D��B�ф[|K�;z���|�O��c����r�v1�(��c7X81~xBy#;r���'�x	�748)1N��.��+�����Jg+��N�M�7�d� M`��WP�� �[�̣W������k��,I��j��3��u�9�fz;����N|���Y���rpP���Z�
����:�R0Ux"����e��)ЇP�9h����O^�iNcA���O�ǁ�_?�`˵�j1���k�vx�(7T^'�܇R*d<-��E+��"&���֕�8�~��b�	wF܋����y�]c�V2i�)��GP�N���������x8�ƷD��aԿ�1���a��i�"n(�R~]�!Q����{�cj��O;V�Q���j[C��Ȫ� Fަ34ǝw��5?��5P-"��EV/���!z�)��X��l�*�H�ӆ�#l�À��{�r����[��m&	.��-k��{0]@v������2Unx���5�ͻb����)�.�1?�pI�)�GE��gd�z�R p�UxV�V~�F�ܛ���$N�6P���"D����SV�v�h5ic0��	��4��#����G�kZ�g�iU�J�l��E�*�؀��C��VZe�����13�m,<�6�_�t�]	��#7ث�Y����Vyb����RI�m��I,؊��]��Tί�A���+�VP�b���$�B����8�|DX}Y����pY��$��C��&4�4��@
��'W���pۨM�q�~�˷$����ye����-S����]SS}��]2@��/���$���˃{ �M��ܕ��ax��)�kˈQSk�l�Xaw�[w� �x5-�_���j Ϩ��n)��L����oG�ډ�� C':n��Y�����R�f����O�%�GԄ��x�':�</��(�D^ˣ���:+ţ�D]�A1��{U�:�,'��E��O���n�%4ϊ}n#�s\�v%������,����Ѱ���_��34
�Z+��Ի�~�<�tT|XVFl�ݳq`QFzZ�kؕ��j/}E\с�(��ߛ�y[ϝ&�ھ ��I��R6 ��`�RF��L�lt�F�~dĶV:�Cif���m����9��H�O�
�lJ��<J\�,+B����8�P��~��W?��q}N�N��mx��������[�z��%��' Qk�y*��[�
��_�DI�Á󀡆�����t�r��
J�_B��)������������Y��h���F����I�,�G �o�l���f�mLrݔ��U6�z���U^%�O��ة2�{.�ͬ�X~D.��`�� 4./�[�q����8��m���v!�V ���9θ�>(��"g��EG��	Sܢo��8� y{�0��l��Ω�O��gCs��	�t�:SZ��SŮ"-7h���唞!�'�
cl'��#Ȃ��o 
#�t�� �4��/u<9��'���3�ω������n��-�ɌZ/��nU)�P�����q�`�$���r���9���5�Cգ�o�J�O��Qz�hzv)�s\:e�E�������/<{߫--�17pY�����k��o�o�,0*�U6qX��?���0�qQ%w� ��y[���iw�T]>G�Z*I�,�?�Q��on��|�8t%Q!xޤSIL<����V5��̹��f�y�e[9=�@u�5��pcmG<�8:��>��%o�X<��i��\�U��11�w���~��B�aW`7������B��4� ~�nP�����/WHx��?5�3���=3�h��Q�j����R<���la�o0�� �9���şNH��kGT�"8�??�l
]I	R�q�6�D�#�,K�����K���4�oɡ������Tń��"]�R����̙t��Y��k�Dy���c��<2 �uǙh��;~j�ss�3����`�fB���'n�Pfb���-�:�WP���kh$�:��E��*]$�oP�hIe���W