��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<�\5e�)���������Y�Y­��i��=�����,�N����K���ëb��<{ڼ|=�~���kѼ�?=����=ئV��|e��J"�d�~Z��d���*�:��S��q�ɲڗ\v�*���dR��S����gG�/"���L�[߰j��+�b7`����.�x�Z%o�#��ɾ�*�*���<^��D���C��(��^�g�.Ȣ�>0?��ae��J�����7��Z���h�Y(2b�>ّ2d�`������� rBn�Îhх�����ɞu���F3�Z �nx�k.ji�A�V�=�H#o�^��>�PN � �A����o���q���T�b�ګ���Q�Rm�l�C[Mf�+�M���q/��<��#��������������ƺ��/Q�����&����m�Yt�Bp"GQ_���M��z$�FѶ��sa��7�[i}{��9l�R �s2G6�0�T��F}fd(n�W?0����|g]��=�;߳�s�X(�6��=K�6w�I�,w�m�*!-5ܭ
�M{C0��wkH~���.��4��ա����� �t�-����/p�~/�}������ϸa�6K-5ga͖�W���reE�UB��
����CMB�"c/,vk�n�u�������J��=�.�8���A�h�?�<���-B	�R�?觹`�^p)�&I��e�B�f�
�6�:��=2>���:���(������ 7�e�;�Չ�t�a�>ӗ00�=��n�c_N@�\��.�]%�91|(9)c��I',���OϞ�Ě"=t�jx�J95|�u-ՙ������'�o�����I�M��zE��ke|_#�J
|D4����B��VA�c�\�݁��)��9��U��۹5醽�ۄ�5��j����AC��dv`�G�?0j��ԧ7?� �y7�7�Eg���%�M UPi�k������w����"_�dx��K��?��Tش�x;��6
�(HE�b��4)���c}m&�i}�'VK����n��g��O7�(;�� �O���.�q"��z١����4�D��.!�HG�*J��Z�&m,��Ԝ��rؐ�������x	 ;�Ԇ�Yhu��)�v��M���7_'f�3� |�GR���Y5_d�z��(����G��U�]
��u�,�C��|�\p�^�b�V?L��ؾ[C#�����o�ScS�����������%��"c-��ce9h�G��0���5�3�����7�IvP�?԰�D��_80��M�c}nݩH@
��ê�-��	v�j��Mx�&7��F���d�{�*�h�]Q<kv-ˮ,�����-c��E�d^uDg��Y��Y�|���.��Z���b����9%}g��$��s����[
0������,�u���FL׍U#G{Dqc1ޘ�Fnǜ�L�F��h�JE��R^EU*{�p������Ew�g3�$j�+%e��5�	�L
S�����c>+���K$ߠr~�����Ћ7֌�c��V���3Z���)-�Q{�O�+�Ĵ���.���������!��>E��[Ej?j	���`���z�M.�:��&�bVt����h��h���DBpl��ʇY����n/�1�������A��&7�9�j�4����5bb��m��A�"i:~����<D���.� �5A
*U�����H���)}j.c���I��t�]��Q���x�~T5�a���.�1����s����ͷ��8wo)N!#%"�9bu�n0�c�n�X�5��jm��g���=�SB���b����C��D�U�+1m攆��%E����=k8"g��N��P�o�h$Xc(I:��0�+[�;O��i��i���-E�3� ��}�=l�gf���Tk���NY�^A��A�'� M��|�;�1�g���׮�
�ٴ�VP�!S��$��ߴ,Cm�]��:^G����i�x�Ղ���B�4�	$�l0�5YF&��f�yF���2�\��mw�ٚaB0a���w�(��,�	����n�c&���g�X��t�V	Md����ʉ�-٢�����{��BJ�U���������n��_�X�ϗ��H����w� UO�g�5�v�-x��?�`�hᾗQƇ��x��Ι�X� /Z���y���V��9����[bD�a�0�	z鉁q����.-�UC�+�ѷ�O��g3�c���N�������:�<����a���k`1k5a��� �2v�ҖN��>p�c�,�WPe]c�.�&QX���#3\�!�Y-�n�Y'�ǫ[A��Y,N�ä�i1G��e��>j� ,����@�����u<Aq4����fY@>b��X|Q�ψ���'�Ђ���K���K<�W���q�O�a�4����Vj?��"���%yL�
��Z#��5hq!�d;�آ�x�� +�"%H�5?�?�6R@�[�rq�_�=vb�$&*o�gt��i�eyR��/tQ#�4QA���A�$�&/�Yw�%�=�|)� ���!�v �ӧ�,��6^�#�.eP$�.���a����Oc�o��� ȷWT�&�����zh0��,zԸUYу��{̻C}�AP�-�Q�L�fOL���"��S�έ5B=D���(9on�X�����DF���xY�ɕ/N�c�m^����9�� ��� !� Yr���V��wB���K���Ah�K��w�(���>�V@�TZ$��Q�yJ8Y7�8��5YU)�-�`"�_o;���}�~����kq�����s�\�b��_g-�u&S*T��g�:n��ɘ�Z��k\���t�f�S`/�$1Fqk�+^PB�pֶUi��ӝ�S�m>�����f�[J���O�b&��=֜g�|j���?��İC�T�dl��V�3�������Ս�k�(Ƀ(	�3`�ބ�((܌
01�|��9Q0(�B�u`F��~���&�r�$o|������P�e���c�O�vy:sye�!a��}�����+��Rɲ���C�G�Q����J�cף���[�KZ@�)>d ��	�x`dC+��zBl���%K���5��H�C�r�M�[�J̃�C�i�
���A�L���_�z}��Ҋ�6�5a��r@޶:��m]�۾D��L��]@p���|w���*��ھu��M�ABZ$�
Я\U%.1�% �ɷ$�������`e�&��418�C�K�2�}�06U
.���)/J!G��˘)�֌D�M�_�:�o@�(�4��D�ե����j|� 2�I bv� �*E(&g� r�n��6��?�&��B`�d���*���K�eN�g��L\��|�I/-o=b@�+v��K�k�[]q�P�
��4��𲙊3�+`*�����M%�����O���*w�p�6B
|��rk���t:�˵�^>�
ZvLpOr&qSs�!�8ʳ�~�k�N��Ƞ�h�Oy)t��\�G��Z7�nV�Vv��Mԟ�������N n�W��N��p�����*�!i��!�II3�2@�_��A 	��'�^-m%�\(��n��P����N�Bv䤱��ڰ�Kԟ�r�#�2r��+�D����͞545�oOR��0X�-Ln�wѭ̲A–��=�H�X���Ù�n8��s�Edd;��a[�H�5*'��|jMXc��ﹼ�ױ\WQ&���"��_6�E䒽���U��D�Ԫ�~G�����u�z��T�1�K�Fx.L��ˡ@�M�I0Fݲ5��O2&�¥�KQ�3��� :b�$�nN����#��Z5��֧�p}K�9-00M4 H�9/�"I�V��?Mp��Q4����0tz9��v�j�a?��i��one]�1��9(�~��s(
��nDN�bS؀�;V6�u-XP��;���-���A �.�3�$A�)e꙱�K�4�Вֵ��#�MJ@�s,R)/g��r��Rg疔��1q�K��GZh���<�Y	���/���������\��KQ�s�d����>�35����蚟�[�Qpl;I��N�ڮՌ[j �\��2���M��/|1�6Ȟjʊ���E�I�ŘEɾǌr��B<ZzQ��3���}t"!<H#��"��(��)h�&��p�*K�7��v�֠{�[.ٕ_c��{(݁�T�0���<�3B�݇$p���<A6Q����&��7���_'��F����:�/w ,�c�w�!%��z�kw����q�J�&��t%ڛҩ2 o(N���?�m#F���3تP�BX[A�8~D+m�Xe� qITH��u�!�	QR_%i%��2h�	��24�@�R��� �aͳt$�(B�D��z�(d����{$�j��8΍���.ш }����`PX�B�`��$�`F>�����V9Vz�3�fc3�d���׻�TK��E����J�y(������zU4�gH$��s�Ŕ�#��?餑��<�7r5f$=R4��#�܎�V����r��@�$0�j��5kz�i�|I��l�)D����s�TTJ[-��K��@�dN���`����r���&hrU>L4f!���u��D�w/�s���^�ᶲ�Û�`JrU�8���asc���ow!�6Z�)һl��]�U0u!}p2���	Ju?�$�\?Eoj���\�@7@Z��\��&�fO8���Ԫ6��)1���	ݽ�����a*)�/IH7�EAzU�ڗ4G�Ʀ��e����2W������[<�0[���䞈�lMz"I~��"xE��	F�]L��^�tU̓�K`��Fs�y�'a��-xn9�;���(�(_gY��02��X�(]���Ä���.�W�W�	1*+��"�T��c��i�Y�i���<�٫���n���Vk��ם�pG��Ji�.r���a��|t;�s�x噼l�{w�ͯ���+�f�P�t�R��	+��,��><�%a�L=�9��P�7�G��-˄��U3ɔ����I�������(�iKؾwO=�`��<MϷ�4D�ns�R�H���FG��(�KŁ�s�k�>�h�K��Ҡ�v��:b�m 67�熃1�l��9Jnҝm�ƀn@W�;�j]�\���J9�0��u�N��b��$F2d�VF�u��(5�&���tK�@�/8��?�WL�тVZ$"�G���7��Y�"�&y�u���\�)Kd�F���#c�X�}�c�`zY�_��M�B#��F��	hp�|1t�A{�6C�A���!�7���6��b_o@�J����VjS�^~W��2NO�w�5G��%�f~I��K��`x����6�Q�`�6�ԆbP�����TvK�t%F	�;�鷍��[N3!�w�鵧?�Z�x"��$��Ǝ��ßj�<�Y���|A�$� �c0/LQur�P��"�b�B����.s�c7~X��3E����7]V\/��ڎ�¯��A;���}��Ӊ�J�=$���{И���������^P||��[�H������'�p?��~�v�R�k*y�hx�̒�p�;Ѕ��1���0�a�d��.�a_�B�'���
D���y.���Ș)��Z/�-�ҁ.����$��g*-�B��M�����S=Dg �1�T5w���{s��N9Q�Kѧk�(j��Hm �����&�Μ����\�Ņ�?��}��-@�fP��\�Kv�>�����q�/ݞ�q����AAy=�o���8z�p7��a�"vT}�/2+4�X��c
l�J��C�R��I�S��ⳤ�]�փBC9�cD��6��M�侉�>�#��R�E#�:��M��f�Z��J�"��(��y1��9���C9B�w�	�\9X�7�^�A�l{om�uL�t���ox?�?U�+Ur�� %J�Ot����'���11uHu
����Cb������V��j9�J���PPv�����]T���5����g���\�Nm]7�'���-����s���������%��7]��8cH�ۢ�C�8�ʹ���JQ3��E�h��'�a*��l�B�6�E����{�>E�.&s>�,җ�[��'��:�s}�O�r�_�ɅKء5u�0э�\m"کC�D�	|��7>SlxK��ger�4lX,Q�a�aKԺf�a{ܮ����C9�N^v��x��YU��R�i�ny}j�e�,&�x�2��Z=;`+tv\kǤ��@��-as۰�R��!pZ����6��P�KƉ�|�!4
��:�p)0�_�$ډ��N�#tbfC-�X�V��g#�)��8��(�4��yqt��0A5���7L�Q�M����.�k�%��$ Ɏޟ�����d�qW��	���q<���i�_�S�8�(�0e���)����2o���	ɏ�)��>�%;*���y���xPN|��?�cYʜ}�#�
��m�}V��194�lݱ�U(y�ob.)pT�T~P��?�`�7�W��H�*�o1��=p��P������������������Y�Amñ�F�^zsD򫐘!����3�ȭ��!R۵ހ�7����a^jw �B��rj�d'�2W�q�[��&�ȧܒ]����2��Z�5���p�*C� �p����D'�T��q��^
k��6-e#�@`��������1/�{��E&g�~���܃rJ����o���~ٖf�f.=�4/�*�@V�k��q4%�Ba�i�0�����-��g�t�qf���̮鞢�+Xj�E������.�&<wP��)0Bi�,��:�㢇T#6֖~�_>dp����Hpej<�X&��q;�2���%d���t?�?��h�- ��o.�+t���Y�a �-	z�3[x��|�Z2��.�N���*E�;��`�����+@�=0��7�-ۉ&R��@f}C�M�IES^-��	��-�����P��~]>�q�UOCMG	`��J�Q��fb���@ˉ��%��֧�{.%
��<^YxxΙꅈ�{[�Jy��;�U,���|t���v'+���8�y{�-/Q�}�%[�`�	 Z�^l�
G�4�=��x�5��%���߯�i}m�95e�`�B�����o�xv�(��7�@������,�!uU9S�pP	��}�:��}\6X��'�!r�_�\�~� 98kg���N�L+ƍ���.�؋�4&m����jv��XNoI��������2��g��{ɞV�6�vz7ٿ�I������M�{}-I��!!��n=�@<T�V�������cG����F9�k[�GY'��:�$w�0 �
��<�����b����5�� ��UP�
���d�hi�;l�����7��B w�;��]X�l���0yČf=P�����q����=�V،T�Ə�2���ƼX9��Zȁ>�T�#5����0�+���˰����w2^�u��Ѣ�OM�[�
0)O^�̀��EI�*2 �:W�q�'L���X	&�fNJ���Y'�#%�_]���|ov�4t�j�B����q��1J\�h���_�X^�T�j��N1�{!����^Qϥ�̓1��r��J��,Yt�*�.���֧eu g��0����2nEu�2AObD*HÍݿ�TH�@�(*����'8�N~��/W����F��r�e:�ZpW/:x�R8�(��q��u�E�<��U��\Ӂ�l��b�����'s��)e�<ҝ��*b<��Q�K��>�@�#�H��7YՎM�$N�z����5lq|�����hЬ柎����U�l�j��X�!���p`A����
/@y)�=��N��\6f�W��A��rX/7x�?�P�Q���K���m�{����]��5�>=�XVAC����s��6D>O?~�p�|�`7��D7퓑?d+���m]�.C�8��oy�A�t	5�z.W"8�s�3L�HUW����T���2�f�P�#'�9�u��Z��g��3�y����'�t�M#����g�+4�Z|�#�*��y�j�Y�~��Eug��ͺQ��0�8��A՘J5��+g�-�#���ퟆɩc��ݥ��'*���R�����,RBgB(��E��p�)F ^|��^5�ie�J�?Pǉ�g�B3��;8��d�]Ӂũ��e��42ܨV8y���W�ז�委������e��o�π�/{ѫ�e�9�K�e&A�� ��i��������J��e����OoC���x���ŨI��U7^��Gxu�M�lS
;�Z������*���Cԁ�bI*�s@{3��E��}�3���u�ʣs�V�*�
�[��s?�*��)�b����g�-U�R��줜��z	8������V�B�Yd$H�͗ɧe����9��c7��Ŗ������M[�CR��o<���t�GSF�57;l2 �׫6ľ���\����S*��
"(�C��Ұi�` 2I��! �~z�A��q���͛��T.sk::��Ŗ��:K' ��3I���hPb$ho@_4��>EE�3u�md1��b��]�!��i�a��� ]&�vߍ�G0����,7D�lﮗ�9��&��N$ř�l�5~�l��J��9Q�����N�:��ȷ޾�hP�I�`�[�^�pl�=�� }��R;����	X��uI���C̫�""��݋�� *&�!�F���Qt�lK�(���\��\ə�8c�4�<.�p���i�����g�G3�LY��`#�����iy�C����ysM.�H^�a^@�����@&��Y��1)�c��mr��^�l����qFyפ�v���I��~�-�h��IOC�d{���TWy�L���ȏq����?C'��y������Td_b���a�}8��f`B�t�[�ޮ,ej�i�yt,�ɠ�K]ŝ�mC������l��ܻiX��Rk�M�T�ǲ>I��O����ن=ܩ�4-����~��|�}u)�y�GZ.w�ӕ*����)s
$V��Ý����hh:2� ��%��m����	�\��T�Α{��Ɩ�P�1��4K���{S�$�V�ج	=�g�������I�T�]1�ARE�X�m�����(��b�^[�&�i�-ٯ�9�8��9�@�#:'���=�I/�G$�LJ%�s�^T
6y�S�tk���P �Cf��Vj�N c��B�N�7WPv��k�Dm�Ƌj�d�I� ]AEx�
ym�S�;%�M?�y��߁�͟���6@��|M��v6se9Ȼ��ε¢h�p6'�^�01��G�I�R���ys��j,.�|��/�n��9D���3`�����E&��~ ]���}���"��sXL��0�4�s�S����ܚ�2	L�jP�ebɉc�
�p,�1� .F�6��p�>P���ӭݟ?�"Q��Wݛ�ʥ8`N��L}��������o��|��n���p�-a˺�:��a+�r���|�z�_G��3G���������2��Z����ƬWA���G����<l�aFJ�	4)qD'�=Em>B�P�тh�4Y��<��G�ℶ�Sũx�3�O��_���Q�c��X��o��B]L-�*�؄9C>՟H;Q�LĬw2j �����)-6Ay�ԥzH$9�i���Dl�Dq��#��Q���ݐ����CH���.٦���5�̗�f(ﻐ{y��!���+5���L�)�`_����wu�qc�_��[.[�a^nE���=���t�^S_��F<Zv���r�t�(4d�i��k�F��{:�;�* �h��>-����o�4 >�ේ��I���rF$j�T�+O��tW���2�x� N��h_��l؎��۸�{A�Yd6�9�3���C�p�-K���	� T�z������;��O�#i��@V�����,mJ�,��X�P��(��1;&֔-����W�4k�Ҋc��o+��T��0��X�J?-�%ժ-�V��X�H	��u����(۱�.ί[���No��1,;�t���y�(��2�x�A=�1j� �KofjHɢR��g-��$��1�=��-��*���qY�V��Zo�{�
������I�@�����3*�%b��@6���h��Ц��y�R��l
l��s��h����5���2nX���\�j��R�p�|lT�>��J]����=S�����m6+��C|}��u������gk�0��.��ǾV��Y݅e޴(	^��g�ޔ)��"J�~�]ܟ��[��r��c���'�#&j�W�,�Թ�k��gF�a�{5� a9�C��/�6�A=��T�)5��E��4J:n�@���הd�(L<��F Ǔ�$ �̔v����r�+�X�4�-ٷ�J��C
b�JF�����e�����^�o1��d�6��I�o=I�է,�Ad/�7n3�E��0��.ӄ��7d�9<!��C�����Ntt����4�	%k����'�.u�����g�[ 3����[�A��;Vw��#p�>���	�mߺ���\�����Q��G��f5,ZuYa�?��J��O��)�R���Gi.u���..�.)FM�ǫ�����Cӷ�t�<Ǎ�s��'q� ��5�C���ɮ��l���]q(���p��Ȯ���ݬ;a'L�:K�̧�D�H�-���������i���4����?DV����9�Y�R�D�m�f��}��fG�kÖ�x`d�^PLa{��b�ڡ��!�����uE���;C��R+R%�C3㓓>Ӹ��A�T"��9�P-P9}*��e95U���llj�`O�������n����"d$�[���O�tj�l�J����� A����p.�$M�pG��i��������͐�-I�晬d\ǎ�^� �����{�0���YDd|B|D��d @� +}��ѫ��&�(�~���?{x�SJ�$����g^X��v�Hj�$sq�O�Bj;�~�{���ٺ��UdH3H[������a�]�$��r~IP(?(p�׬JՍ
�؁�����>�ƺ�v�!#��f���U�IY�D��`�Z7%Q�"v����n���1���i��q����Ӻmv�<5z宖�G�s3E��y�]�T_IK.)��,5�E)o���vF'݁d�X���ח�N}?�.8����}O�J����d�8�j�П`�6\[oD�4�ɊE�bF"�`{�ߌ��Vu�X�0���E �|yU,�6�I�M�z9�E�F����m���6nkd2�y"�_;�>&�7AL��z�`�����'"$;�p�#1����+�K+��aP
>��y������dK/�p����g��A$���K�����KI�9��wK��}_1L#3y/�҂8fl�Dh_륿�D��*�-���S>LM,P0<�5��EI���V�Z�=5�e*v�7�3���"���Iz���d	��A9�CL��/�r�L>��ܨ�ӍF��3�Õ�̂�y�b����F$���'��(�C�O�oC��O���s�Ӆ��v
��܊��H��3��
�:^�d�!�#�y.0jYj\E!�٩�d�|5���w�M�=����j/i���e���n��7*�M�ϚG0�eA�y/�>sL�zj���N>E^��B�R���\�O��'4bi�i�"I;��%� �7�e�xI߀�Ϗf�枴)O`��S�@�*���Nie|�X]�U�}L)N���)jh8��t�x���ը�
�-�؉��f�3���f��eH�P S��l�����	����v(��XG�x��F�ҥ�{�DU`�2�� M�L"��`��7.��	S�?97@mэΊ��`�'?_�3�X�ٙ�c�������Նï� ��7IܚOU7jش{��hk�|�r�&�#.2��U4�:�e�7,�#�"�!�ǃ�a�ߛ�5^�!�0�>�15bIu����>?O�`�ͭ��"�;h�@O4N�c2�D�c��dљ1��p��䮀���-���~�N��%��>1��[� ��l�����	�oO�8}�w	��&���U������mDX�z�lZ�)�%'G'Ӭձ��8�L�I�1M�V0\����3�)R�A

m{V�&,�d����3Bi�_�.ѹ�Ak_@�n���O�%hq15"����iޓ,-��HX�W���W���?L0y�FI�,�G���W<��L�w����,Y��O;��=�E���j"F��?-W}���d�I��sl���o���,��]x9T�h��,���I���Q�2���4����z����Eܕ�U�>�@��h��`S��:�7�h�O��]���T�{�
���@��_tp;d2X�δ�pm\U�iP��֪�w��}��K�6���_�����Ɲ��B�IB;������9hhi쩴ʺÁ�n����k���3�U�~z�^o���2�+���2���ڏ
�>BDdI�,�K
�� _檡<��/~ �$,�w+{��|�?j|��32Α��#�[�iW+�С���~}%����Ϧ��y�5���k�q��NA���,��O)��K5Z_�XNs��E��x����SK'WV�{8�G*���j�ؗל�e�+o	<��-XB�]�;h�14��v;��?=���G�d�pN=ZF�`F�>�rBB#O�����$��J�MO1m9� �k)�nC�C\���s��37ɻ��Ò�C�N�I�d#䯷V�\%�#����� �,/Q�!�BıA�8W��/B���#��琫���M7���>���Y�0���6��G��H[���$�����$o#N�'w@y�1M�p��	ۨ$1#8��i���W�6I���b+� �
�����~�].��kl�ϟ�w����͉�jI
(�F�wɰ{��+�G�y!la�<���Y��_���XfrgW�*)�$gPJ�E�	�0��%=k~#�;�;&��X2�]mZ�&�Z�����<x�LI�B�tsM�������N����r/�3�~]��$��f|8�M�W��]���<y�!�U�m��b��e'���B�N9.k��+�pe�W�����	��].$�(*T�j����,���m�&���������<!}/XÉƶ�3ģ��Ȭ��Y��q{�����Y_}��*�*�ȼ�X�v�.�[��??n���r�U�@�Ԝ��|��1M��z��3]2F���&2�о�� ���+>�0(��P��Rvj|�Ѫϱ�s�!S��L�W��Ȑ���<�#Т<P�؆+ a��c�k{[&��U"L���t�d�1U
k�9����|���0Mr�H*�͢�+�vN5�ٞY��,�����,���X-git��h���}�
��q�JD0����EesH�3�I�.l�6'xPƖ�4(�߰�[�a���I�tv�v[u'��<��b�&D���"aC�u���\�Y��:����o����?����o~_ᖋ�A���� 7�ف1	�!����ui�A�:�w��rO%~d���a��b���Z�v���:ԣ���c�J�e�M�Y)[L�C&�Q׏�%�	G��
�[.p��J )!�����h��؂�'�ֹ�?}������µM�2�3�}uh��>�O�g�P����s�v���Ԇ�8>��'�3Oy��,�(�N)�5(Y�FS.!�f�nڝ*�76j�f ��˺�cÔ�����I�Go��s�M��L��y� \Q�B�������j}�ϬS%$*�b�C�#��AxZA��m�B��D�n�\zUF� �e[D���X�g���||d�V�j-9��gL��A���Ө�w�{�8f�%��\�kz�4K���X�B�g*z�.���5��N�BA�7!8ƙOV�&��|9�A%���1*��Cḻd#C_�'�쯧�]�A�-�XD�6�I���^���w��(kZ�ĥ*�:�b� ۴�𢹾��{�� ^�f�&Ξ�L��?yå�5��ё'��PEc�9�ҭu�ʛ鸔�p湹9 �QA�te��<#ؘ�V�'+�@G����G���]��yq�P#�Zh�h���'^��pc�ãai��xi$���m��=�"�d+�RNҕ�zw����^_t�T�A��?��\� �_��i���cW�$G��ǧ��3�v\\�˼"�ay[��]�{�"Ձ����h���T蚧��ϘD%<�f�E�R=��a��a�9��J2��ӏa[�f�P��s�BЋۣ�}�X�#6�|�TH�~�"c.V�M}�������0�o7T��ym��'�p@���=D�2๋P�=�\09'�C�<3�,3�<e4��Y�
�ϛ�}�{�C� ��O�P�w<pw?��A�u���F�-v�e�W���Ml!3��<T�U���������ਪ$: w��B�s)Ĳ˷�v�I�A�T��C�x~'���8�H�?0!b�Qm�JKM�Sp�]��7�H�R��:�#��w��`���,1+��*o�3���ߠ}{e@^r,�{іi��/�PXa�Rb*\"S>�/�S��� v�D
�=2�dnP� ��a*���
��5�[&�����*ߌ���V_�.ڔW�Ƞ��}�^C��We��:�w"O2Ts҉@F�eryW��ӷ���w��GB�F�\i���~Eq��݊�b��K�!O=f�:ŋn�v<�71�s�G=�b;�4��z�In��Z|��5'!���o6S�EJ��tT�9�o4�,�E+�[b�q����8��*ʅ��0=�`�6%t��Z�s]���H��ޏ��ߴ+,n��! ��wƞ�}��W������.@
w/�
�s*.C��� D��|	����c��������6�;"�,�T��!+mH�������\�Zyp�B�x�#׶��".w�8.�����4���!ؼ����-m���ŉf�Ez/�3�����,��'y(=SαZ�L" 쭵t��3l=�@j���i_6s�1&�l������7������Ի*�-�:�Y�)%v��V��I��n��}3&���y1��g3St�
�m���hɪ�n��Ͼ�_/�뻽pZd����vc��k��������I
I���8��Eai�H��-ʱ�Q����q����GRZ�����xY2�f���8�GE�&��"�~!-d��ڡ�'H��+>�r�{�5[̈��*߬��d	n<��VBo��P�g��8x�p���<�N��g����ڸ���2J��w��ȵ���.����t0��4�Rv��=���b�ݙt1��5�ѩBpJ?4��OxW$t�HJD�I������A��k���jX��c�F��0%:�-ԣ��b����9"�Lc��
Ge�S���/��g�8%�$rVu ��?�}O���7�LG�jo�׍��I�|�/���mZ�
3�>�ҹ����3O��z�|X��󧚃��]~qc��ۜ�\>���:����8X�y���`����A(�\����O�yY��:	�c�|�zw]H��]}��\�Y)/iq�x�Q��VC��A�F�Z/��g�9(����Z6r��Ҿ���p�u�^E�0�H;�7,<��A���d:ͮL���* h#C�V�$!	3�&���`0�'\mQa�&17+`D�@I�,nu���ޥ��lj������y] (ݧc#&"Qo'o�g�����9#�l���~ޓ��t�#� -�r*2��\5��+˺��۱:K��:��K�����|���#��[
5���v�����/Heuã��R�Z��T�u�u��¸�{W�$��f#�	��R��O兓��I� ����P�Hq�K��,�%3ݳ�M�T+È�V��g�ȉ}��t?���g�x_*��:�[�*:��mВ\�N��.��]+OV"E�Kⳉ��'��sJ)��V������|AN����fN�r�g[M�~��XH�5��B��2�_�ރc������L������aʟAy���f���p�� ���*3Q��ye9��'?��7�.r�G�T"Q�t"CH�A�]Y�L'܏DH_�C|����X����h�#\�o���q(y�|3~�a^��~`&x��X�M.Z�Qcs`w�:�p������w*����;XG�Fy���~�x���x�{�r�0�lC����:?���1�b06w��߰P��tLW���4�VĔm�GZ����- 5�h�7U�E��T�F��κ��A}TFvz!�p��Y�_���7=֌::��PR�s�Z��k�B���;'��TN�`��w���<�K^/gׄ��iA�[4eL��''��Nz#p��k1yh2Q�(�xԞ�d\z���5�L��
���.l����K��Mu�kv�(W �����z�e�}ᯜG��������! Uu��͘�%9���q�T2Mr�P&|���-YzC�lg+�9�U��Jy�z�ps߫Kb	����c�Uu1	ݓ�5>�7�;�%�zQ�|����̟tpo��L�]�a� a�?g�7���pVȂ���-���O�lȡ=~��S� �y� d?�=�)wF>
�a.��b�����W]�I�T�G)t�E�Ϛ�	�۳�]Q�1���U)f�{��*�3c�;�Ng���ņ�u�<" ��&��勊�([wtt�l�"�������>f�.L+�)�p������Y�.{��	�T��Q2wɆPX9b�D�db%1&�W5�I�L��u���[����7i@K���G��H�<k����_�����#��=�y�;�������_�{Ok��!�k�(��(�Щ�%Ŏe4�*��n����F��K��@��J��1~��0L��Ӽn�D�o�� Vk5_>$��.p���CO��n����'P�P0�
��Ղ,�oFyn�<$�5���ԩ�(�K�r��G|�y�m��t�L��h��b�ԠC�5�"�SUw~��ZiV4~�|����3��`�P*� '�7��]�=���t� �����n�(�Z�POR�c��YӶi8MՐn� 9B����v����Oc=��&,��r��<o�^��8��eCc��$z����Y�� ����>�8-��RLV��s*��������9�1���2Aʙ��kx.�~2!�k���'���/7>DO���2�xe5A�q��H5�$v?�����,F��bE �G9܍�a���dt����~�s�AAf$�@��W&�N"�?�NJ�h�n�!ae"ud��.6Ϧbԅ;���4�������nϧ�dY7VWm�A�#�{1�'�M�v�>^F!6���~���>��;�X:�٫�������Ϲ,�u���"4@�ۏ�LB�i�t0O�㗫<w����l�|`��qYfٲ�1̱9�Wfj������kT�<u���/&��1�*Pc���&x��,ھ=�-����z-����Xˆ������W�.��)h�����빸SZB-������Z��qz�V�Btg���,O,�9�z0P��-ȆUܟ��i����>��9u[��v�{xDT��N�Dx�D�vќ7`4�ڄ["X�}��^�b����D��n�_�fOs<-0͋Mi	�	�C�����ZY��,��	X�s�L�Z�/�K�տȋ��0EKy����`�T��|>� +�#�	����{���0!�y��wc�1���XlF����Hl;���Kѱ;����\C[�ҠY���̤��(�D_�7��NTʭ�D ���^���A�a��m�+��,�L����øE&m���G�{}��,ZY���̜�=���2��
����3ğ��uԷ�C�ޣ��$�x�ͱ�������YG+m�jFb<�L���#���6:�����ܼJlHW���:v[�����5:g�n+ �u���3H����PK��\\������w!w�5M`�x_54a����V&T^H��w��tʚ�!א������>�����{��rZѲd'��6��:	=OJ���]@ 4<@ތ�<�����iS.��G���i�k_gt�(KwKo��y��jrhsV��������8�&A7v4em�y���*`��27���n��K=�
pi�aɎ�#ԏ�kJ,k7�v��O���_���얢wc�R�=�e�7#���e,0ڎ�O��f@Vnr�L��t�������������H�&�T}�D��7'�^��2Ȃc�/�����WlW m 㑗��>�.7�Jh)��z��A"��.n�/[��#��:)��FY7Ԃ|��j6(9��d�<��yG!�B�H��ŕ���w�DYf6��)���@��N���	�Ĵ�&�Zٙ4�� �T��E �Π��7�N�Eo��SG��� sK*���!��7����%�