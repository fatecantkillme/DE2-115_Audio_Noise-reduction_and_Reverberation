��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_����m�e"kxu�Uٲ"#oB2�-g�j��h�p� M T�(�P�+M��&�[���+e�ҿĥ��L�.R�d��HH�~����1^^�]-��s�T;υ_�� g|�H�\��#}J�� ���@���.��P���Mn�;gۧ��@�%�vv��0�*n�� K�ؼ����r
O����*�4Me�,X|�-�]#5����0�ƌ�k�&\k����7�pƤ�H�g�#Y?�����r�*�ٝ�u�g�{.A,Y�,���? ��ae���v��,�`C�����f �Tu��<�,6��F��S�
�b։8M�S���׮�,"��!N�J;9���O�QTP��2�_1.����ug����L�a���ui��aICU�*��љt=��ؔ����Jk�F�0!VJ%�a��kʧ�ޡ�m�s����j�m	H!p�p\�T�s?���$)�!�`%-����'8�g���ڒ�o�_י.�F���{�:<���&�h�䜸�k؎�����b�����*92���2B�2�n��&e}Gj�	��]�ou$��7̛�%�x�9R���us����t���N`���t�����?`�_�ɭi�h�Hɟ�L��C�Ȉ�4�#�#�-�������;0G���>�*jPU6Z�/0Mwvp<ٱ:��W�PV�d$P���9��^7U(!�>j����5��T�Oz]P^���[{���E��%�\�2�Ń�ڕZq�B��\�q���Dٜ�ޣ��p�.ML���(�ϜKo#��轔h��
��B���ѽ�O��4�M�3+��X��$��
4�}�A�@5otM��g��*����{`�ݟ&��Ƥ#p��bϫq�2�QP,���b�7�Q��D.�?E%f�}�j���|�#:U���R��>��n� ρ�
_�ˠVp�K�O'$n�,��	����|�Q�.��L�����`�B/�̏n�x���pO�i;��j.��ܰ�=��a@�����%<8a��Ҭ?Tc�La{�k@`��G[��7ݟKd��
T��>+*۟_'�Uf��>��Æbv�P�xj6�����wl{�ܥC<}�m�=�!_8ӄ�4R��Y��} ����K��H"��D�)IN�ţ$�h��|���<k](BOm|���6?�� ��P��=
�
kF����9;�P����N��;,��� A!��kxvk��!�'���3,��{Hm��P��l-�(��PL&��k�P'c�K�4��O0�a�zg��qC7CP�u�J1l1��4v瑚ꭨ���Z�N�W�*	�Fi��O/�k��J�Dzz�~��pm��nE1hq��tD�6�D��u�1��G�,0y��ȑy���PY�rV)~_�/��� �pq�x�����A������O)���z�=h%��n%k�S�f i�,2z4f'u����fI�����(��<l2�Ѧ$���e|�j���s��0�m�!�ee��\*v��]���h�3���L�՞q�P�m�R�
��j��r�[��f��ԗ)m��^��*����q/����*|���֖�
אQ�ic<�h���͙DgFzx:0�����ظ?��2`�a�?�^E��:�OY�F�ݸ�7�	��kő$�7�Ԫ\�w)�{�ʐO
��.٧O��p�<���(�D/֟lXp�@���i�=��^�<a���� P�ӗ@�q�w����U{���o?�a��tJ)�9Y�s��� �e,&?FN��u	�솊��ݑGW��b|�S����J{��LdF��u�n��؅cZ3�D� ���g2�g.�Z&.�}�K�ᜌÏ7!��wC{�b��?�{�S^|���8�|�>����>�G�H$i^�����FF�����*Ub�VY6c"�$�֬y��f�.9�7�r7q�M �ڐ��%��J`Cm3<5\�Y��n��f?۟�����6���,C��K�=�m�5*�
D�Y��K��fC�c�DEb�������N������O\��5��j�H-����yE�A��^�Xl~'�8s���&�!��H\1!�����g.K|̬a$���׸q=Ы��<�#�1���ˍ�D *M+��W1l,����<!D��@�9�sJ�N�(��Ң�Ϋ� Y�<�J̪�µ�� DshK��]�V�WTa�hO�߁��T3���v�#�/{o߫bQ�[W~��r�GzO��xhƙ�7��`=��