��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<���=a�bm��Q�BwU�xVI�`W/
�Lq�;;a���.�-�	&��X�j �@0?�RP�<��?k79�����h=U��a�9.���~6N��p�
���H���K~����yXP7�����V0�>d]\3U�FX�R��"��ø�O ѳEl�)=�&%�E����l�u;[�Wƨ�.�H�!�Y��!��U��8_(�(x�:�{��DRE]�먓Q>t)�K7�w�u9P�Y���Dgu���r�36�z��5�а`�9�ZbX����\E3q����,�����+8�X�聽��rye�k\�9�SLf�9ҁ�0n|�F�3�{!c��u���³����=f����4Kƥ���OA���L�b��xO&N[�>77�bޙD>t�F�f��Ըy��?S��Y��q"��c��#�����<i��r�_Q�-��U�����v>~�'��NliP_8����9����A�c�d��3�X$|��1k��5y<�� ��P3j���M����$9Z�f3�'q6|qZ��pY=�
��>����<R�qW�Mְ�|��Q���0�.[���(��;�P{�rS<�2��m	�=;)+"� ����ek/s���_~�,t�<�	��\�\^�	�s�?���< �.�H� ���<���>]�F�t��?H��[�+O���P�@R�p@pIoP�	�si����/#!X4�]K��U��.п��ܘ�$�ͮ��E�s�Wz�OT`��z���{�|��%��(��C[�J;V�SBk�I���ojj�r���L��|xᵭAПc:?g^[e�Q���=���	�m��W╽�V��M��hj)*��`�?%t��X�c�-���\����X�;N�?�O����,,�-/jn��6B�e�F���~]�?�K��y�I������hA�ܡӲ�4�V2��n�4}�{N�;<*�亂�v��/T���M���ױ#2�����C�� ��U�<��jQE�aD1$7'�8�WezE�m	�@��B6������X弌aN{��%sx3�`g�/���.�=~�d�8D�H��s?��R�f��y0a��9���\�D!�eA�T���4Afل��u�Ķ�P��}���-wà�Z�������%7�x �&nށw6;˞�Mb�n�Wq4J�3565�OB��n���>u���s�AMDu�t��<5�!�*&%1%9ʙAV�GL�����]��ҿ���ʀ�A���Ivyڃ˩>���EyI>o�S�wtS\؏H"4<#a�� ̮���c����-P�w��b%4]W	!����]K��j6��g�S�"�	�/	��Xފ��oڮe�\��w�Yԓ�4���'�������^�DdK���tO��
��-Fv[k@�bʖ5� �;5���0: =���q�Ta�O�K�
��pM�9ΰ\](NR�c��\"��@���M/|�k�[����N�,;�jL��҇�D�3� �O6�A��H��q�fRoV!V�e��Y�&8���	L"I��Z���O�VA͇C�b�!�zQ,�c�jO=~�pxީ �=r�$z<��&^�������_�b��Y�E�w�����6.wr����P1�ޖ��*ZBURh����ٴ��8�f:b�O���*-�<�KVI��×5�gm�l�l�HQ�R ��A.�Ƨ�LQ@,�_:�t�YO�(�'9���>���t�!�T��h��;�uoɄZ~�զ�ϔw�7�c�>�[WK�̓��=5;vϯen[ŹZ�j��MV�b0g]����yP9��i��3/�w�)�AG����E8y��K�ѷ
�>>én�<�"6?A*{=�!����.b�75��zݰcς���ɝ {�R'��a�6���A1�!Ѻ��1�,�\�e����s��\L���cIZ&�)v
�%����K����o��Jv!.zC$�0��+�k��7�a;ٍ���{�����3�ק=�Eoi���G���B&_�j-iJ���K3�.� ��I �Kw��E&��&��>+&g���l��iC͵QF�2}�i�[��֟ 7f�p�3d��)A��+��md��ω0e�w�zG���Hf�vv{ �, +:�����Z���{���}��<R���C���C���F�?|��ԙ0�<��ގ��3	=!H�
��&6^ں^ճ��g�f�7�rl�8�n�c��'���Jt腱�a���[,���8���@��r�V��h��Ix��cK;��MJ�Ã�����5�Af���#�[jT8�����e��:Wkm�kH8��/(h�;�
�TH�*�W���Y��@�sF�����e�����peg�B���4�-_�,$N�CԐ�A��G�9�P�����������7|ъ�G}�ѽ��ď�i!ɳj�B�����3�KsIbb>Z�����;�̚_�C��!߽O�F�/^�q��ze�P�?�6J��#[���礚/VG;E�&�P��Z��������'X5���DHGnU��^S�І�����)tm���2�W�ބJ�+�uH�Dfd��e�|R��v��p���jj#,Y�h�D�<e��>�+��ѷ��Y1���g��V�T�>_:�m��t���A�S����ȭֻ9�aA	1ݓ,�%��S7�<����"��ot�4%��0�%�e�$-�PH�L����;:�d�
C���k����X����+ ����K��D�{r�e�$^�b��K���k�x��b���H1j#ѕвb�2��S�ϛ�%U�a�[P����Ȏ����½S�;�x�@-���Q�ch�G��c��Q_�^���VG�����q���\�KPo��/�H: �����xȶq�U�)>x�h�iB�[G���A64������f|���%�Բ$���4��y;�U��Y��Ej�ɓ���{�|Id#���J��T&]�N����%g�C�e����e5���@��Sթ�oKEs7�.��H���8���&��4����:9A�g���h5U��¦l���`����U\6�s!�8�|�f�Kh^���n��q'�X��������x%��m-�v�#�%�ѥw��9����/��jP*j
	w��E1�7�d���.-��ٶz���q��]� ��X���51�U�"���:͎�Np�qXZl���f7�Ľ&э�¶X憼��Mm�z�Rf
�����:7�$���u-���Y����q�o4��(`����#@�*��I		j��������>�jip"ʮ���}��G�B��3Pq�-C�v����c�dO`�@��<�=w�e�
	}�k	�p��e��א+�V�]k���BE��3i:H
FexN�}�E֤9�~r+1A:������;�Y�{N3��У=���3�\�j�õ��ع7��V���z*5K,z���KR
NM�ѡ�����$���g~Z��ӝY����PEqD�f=�>;P�Ѝ��bf���?��rz�ӡ4��.ݘ�\Ȱ�7�]]捷���"I�K�k�,A9�	��H��������w_�
����<�o���D����L�qY�6��A%�ԓn�g��)+��QP�epdK�+���s��C3�~TK��7�����1y
P�ڽT�S�����	�^�+A���{��拟1����k���%�Ҧ�O�_˜U�,Uh2�3���h�D�[�qj����-7΅��J}i��{)���B���L���3�:uF`�s\�5'����b��5��tx���	['S�gJֶ�<45�I��y��H�/�ͅ�WOy� ���j����6�jb���9ԈSx�B�nO�Jz��B�V��N��������5o�R�.�X�?ծ����X}��Z���8���bWr��X:	���E���_&,�V�F��D�[Ɏ����Ո�����n���>��c��S��d��o��[�j$V���^֝��K&���E�vW��e�tvD��}��td����9�a��C��?�����?U7� ��i��o�C2;�B*g[����>{\�+:~Q��Hw�G�|l�j?���+(-rhlK4��+��a��j��-TZ��ǩ�:�Z1h����ő�bN�lrr�h�/�]��o�<r�˳M�H�'D�T�
ܮdI��qe`�(���K��iX�D,
��e���u`�<a��/�9��' {Dj,C,i儚�4߶�E���S�����  �;��{M���{�0b�lJ2�&�w{�k�C�1	hV�`���;�pv[��?.�Ce����7��GlS5P*g��p6,�J�� 7����������m��-5��d���z���M�UX����}Ja7({�n�e�S��p^�}v�w��Z����z�f��m�&�{j��k��i4�y!9�U�
{x,���# ��3��5HV@ޘR��`�A�O�9�t��D������Z�-��։����~ �*3e��	�^GI���yo"�V��%�Nq����˿@�X���\{��_���<�j���m��C��Z"+{�h����n_�#)��,�6oasvh:�C�jx� ��!�����-Y�>$���L��2= "��ӚM�O���w�����0l����S�R��(�>S䓦�]�B���\l��s�K�pc�&9���h6,S�� ˂�oD����A��`�/D����VM��>C�]�lzP�I�6�K� �4�9L���._��g�9�ħ06�����z�d�.V�"w��a	�B�c�|�I,5�3�&I�r�)�oy�>7���z�����*Ӂ���Ha�9��<>FI4Τ|nE�	~�����nU^��v�k��*���,�?잚�c���
Z*P�n3Qt0|��x�
@���g�����kffn�T�T<���e��u���1��gc�&�I�@�����ɹe�(��E����v�V��D�9����4�_;�*�H�L�R9���6�_�����ط��4)���m�j�')9�JH��%�yRM�*�H�uL��d�he͉`���������"��	{ݗ������r�k��(���������7 �?7]O�L'+��3趄T���+ Tv�A���M��-�7�b%B�6���U b�{�\�<�m`��A� �}�~*�x#X�)��l���g