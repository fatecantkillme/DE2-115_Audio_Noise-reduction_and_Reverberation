��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�8k�)9�k���J�f ۘEN�R��>�Ug:�&�1��i��kʣ�!�I^�,�_y���l��f���I���d!sՉ��A�z�RQ�-(���^�ih[g�����̓G��Om=�h���F#�{�VQ�͵&�D��з�$s2�y��B�Ѻ;Z�U�F��}�L��K9�BSI���Y9�7�{���B��X�C	R͑-(w��h�sA��>t�;�`���N�4�j��]�f��f��c����p����I\�N-;������G?9�f��7����;�WI��P���X���A�)\�0�ӱ�*�=�;� �-��=����d,1�3>���^�\Vn��+���"c�o�ȸtp���^_��c:	�B'���ψJ�&ˁ��=3�ч��au�]%T�Uml)~_p !�*boX��G��
��u��^]0E��{�ɉW�H�f�����T�J����&1���'�'uF
$:��r3-��K�j�@���a �m&��UG�^� 0��
#]D8�ϯp+H.o�&+X��Zc����n���`��`aǻg���<B�n@HB�\.5�	@�0����&g�|鳃S5x���&8��:m��Xk��l�xG{��H�����͡��~~�mq:+��
������)�:�F��0�ZW���?�b��_<�4�&��zHV�cz(��C��f� V�?Ɩ��r�'����Ie�_�ƮA�;#eQ����t���#��L�����
����oC+w��=�&*"���M(�4�yS�g��{LS-q�_��3��cp�0�1;����c+/OV����AO��P��t9�!�%ZR[Z�9>�mt��~�_�p��[e�/ttg	Fj�A������V�Ӄ�ɏ�������\=�2���Ʃ"��W4����X����9|��{`��|��+�b)e7O���0�︗D�
O�'�ٍ��H�{�$Բ��m�c��� ��[;��Ik�5�iCj��-�Q�;?Dȉ>h��!L�'75��k�UxqW���3a�7�2�b���aNCի��V�X�������.�A��5��g6���8�gzZ�E�'B^"c�"`�n6l�q{�������(��+@C�&-;;&�<��;G�&�����}�@�m����=�F�k����l ]���f4���t��bZ�>� �K:�����ȳ�D�G��W�Y7g�����R#�����uR�D�6�.�5M��_��0V�M�Z�@|����8��ͯ�W/�	49��r7o�S�S@��,��m&���3&��e��I9��ъ�Xz��0�5��)��$�����U�N�]����Zś���k������4T����f�8�rܻ��ז1��ψ�f$Dt�l}��E4nF-�'~v*5r�"�.�h]Mm�2 ���Z�v��i��Zfćẉ�z��'�i�͏��'�����MB4�9�ů�6|N	g�24�^S����jR��dW���'����C���4b��e���K��CD���Gs�r_kxO�����&����u�{B�Z��Iy�H�'���s�5h~7�hu�e���|6Ŝ�W�a��ń~�"W�L�F=�Э���.f_������_����?�2��^2��;Xh@kV�.>��d��B����9��rRGPwU��>��-��qap/��N?X&���_���N�#����dU��du��7:Ӫ{�v�9<E"֨.�X����*��g�ɵⶴL��v�pa.LSb`�j�o�k�7��7������dn!1~�k0G>\;��LӬ��$�1�Ѱ�
�vct�1��]�Ѭm�������g�ƹ��Ͽ��L>?���#9�n��&��P2�ܘ%V��&V��;B����˛5��E�eI2vG1�m�J��W���qvI�V��Ѣ��eS�4H��@�C��W�~Y�PЅDU��:�ٶ����Q @<���$�@BI��R��Tb�_A�����&n,�>Q@�<��ά�W/��j�|�,��G4CtHw��raC|3��� �/���F��Ȼg�����Mv�٩/�3̲.����wI���]E@WM!����i��[@�ˁ��Z����YE������3,X�ω9d�A��urpk�7r_���k���M
����+z�E"��ӆ7n*nU6+�����:���YS�����E�/Y���<^_��F�/���A�-x�e�� SWV��=�Ӕ״ = +=�(�	��92��5~��'����bE�0%�����5���8N=�zńZ,1ס�T04���eT�IY�)���D�R���_��B�^,��{�v$��˫��G�� _I���Q(�у�M�Q�Q�#L�߶�f]��a�:�6<ly�0��7�څ+|�~�Yd�fʃ��x��1���cS����n�x
q����#�jȌ�8�?�S0?фA���gG)�K�~���-��
I�����Mm� ���T��<OZ
�z���d�=Ҍ���T]Bȋ8��Ou����.4<Ⱦ���U7H�--�h-���\?P�	tk+�^�8��9��B;�4x�<}�C��q�#�l_�������-�u�t�o� ����AT0;c���{57#�Y����35??;�J�\�nW�h���a ;�
<�����n_3�o�^���P��v��M��Id��5y�<�A�r�T �B|�����a���Y�;U�V�u1�����
Y�0)�NO��/ˈ�!Z��wR.�_�-�%RM��n/��["!��%������'E�,�:ABa��ʔ�L0M��&b��KN1?��+��P��cӴ f��w�$����ې�i�E$GJ�b%5��>��Zzk����3@�'h��q�r9@�e�j��_e��j۬%�3[�ɳ�B������:� �>e<�H����~C�o�f-IH�ѱ�b��N��a��JM@��S�Ɋ��� �p��g�]���6
��9ǱUYW��SO�1aP]�����v�)A+��OJ�3���#��n�;:�tm�z��fqY���R�*�gۻU����]6���)?�4G7
_���������E����db
�dc�Q1-?���U�Q���b�0�{L=iь.o�<$�AU`��f��$��]ϕd��5
m4��&�;4�9�.�z�6nZ&������}�}-Kv���Jx8e���,w���6���t�zB���p�*nh̎�M�Z�b✈�S�Ɉh8��0�	+���;/��R�p�}e`7�.�[�rJ����v�c�h�ݳ7�~@3���/����4�Z�,��9�%��
P��W��b˟�$Β)a��]�}bE�G�� ��:+�i�[�"[ ǡ����=S&���mbݺ��a]��w�q�ls���ՁҾ�^?�0e��X��r�nnI��x������}(��!f���nB��ݱ ��2Z��3�����������@̛����Zs��S/�
�䌹���.ȇ���þ�1��X/6��1�d����
���,�A)6���v/���lr	���������f	�L,����~�9p�f��-8ch*�4^���K��:����bd��;.�%W�5���+��F�����8A���"ȥ�)�����$���t�9�8�s��T�c�=�֚�+K�I�|1�M��k�mc����`����T�����c���<�2j���!����NN��.r���}؍��۾��wՒJt��/Na�"R�cx����|�0I�V"!�?��p���t�z���W{�=���j앺B�2`0U�,e�,2��#R�>u��|�l2 6�.=��9�_���]l���BͼΈ�W�;��&������te�z2h3�,��!����[o�H;�<�pX<X8?�`�����8�W��m��de2᮸Ġz�R��`�׿�9͏�	V����(�ZO������Q"%X�*�95l�貅�a@��X)�{��|6j8�:;�R����־k��`�Ks�`nZ�/�>K 	��=�p��`�ȢV�^���kv vV�uC-"�V>M,�h���,�4[�����~��ό	���\�9 �LL��"�i�&�[w��&!�y��bp/3^-C>�K'|���1D_�$ )���? ���]IYo����V�����Lp��D�F���{r��zr����2��zM�_�cáEQ��7���RFq73�47 ����+;]�4� �����)e��쯑���&?k$ň.s�il*y�+�
�"�/��ɹ�e��L{�Ј'B���+M���;� ��&C	,�)�����wsk���?�Ez���	��Q�0g����F�Si����B{�M�ǯ��=Ђf����"}�"RL�9���H��E�!OD�*r�{��ӄ�yq�%L�]R�H\0-ֈDG�,E������BN��kC�B��+�b�����D����T1�t�+��"�V����3�Ml��2٤��C��:e��b��N�9#���е���ci��l�C�S�����)��7�uk~�ڱ�#z4J�������b��45P^m;�vP��Ǌ)=Y����
N�,.�{M` �r�8.t�.�M����̹c!\�hLi>�O���H�*2R�/��	({"�.�,F�GI����UX�66��n=E~! ş�-O���dsw�ӳo��S-m:�+eA����(��c^��R~h"��&s��&��zI0|-:zu��]L�d�f���s� �K,��E�-Ҁ���9�U_r�����K�z��R��Ө��QY\�@���IA�̌ b�i�6~�i�
g�q�ʢ�Q�-��=B��|�1�D>��#)�n-�����#���i��C9���(B�甇�"7p��*Q���`t�x��tՐ�m��U�8�1}G������ �)a0ΰ��D~�Mbw��y/�h'�N��v�b�<h�A�)���C�,�����x_C�U������y��_���^(��Z�al�ֹxg�z�/krxrS�v�B,��5����`�JKq9,�b�f�Q���'�[�Nh���i �9�LЊ�ݨ�lhȨ�$�F!?�c�P���Ӥj}��K��̢�m}k/��km�fTA�͍a��&ݷ/��r�dƍ�y������		�|��͒iY�Ә�7���1h�%Wt�����:M�Be�<���/6QQf�n��I��
�/�
�%��R=i.��XH� �}*�)5d��I(/�>����NF;1� ��ۍ����7�L<���|�rɕ�6E�ȯ��p�^����?{�v��<��7�l�3$k�h���A��\��tL@���4���xܖ�%��o�������Aw$6 3���]_^F]��:�`u�ƳA�Iz~m|[�Y��l��d/��z/�|��ap�8�7t;����h�ռ�|�yf�Kڪ|]�|'��2;�d�̴�[��Y�.K����.1}��m4�g�q�W���z�B��q^��ެ����0WT�����~��2�$1�h^G��5�*�	-O��_���|�����_y���\{���)q��epL�~�x1t�<��Ci=��;ŉW��������=��H����h:"���W�㦪���qHch�h1,B%0����u��@�2G&W��;ms#HAӒ�A��',���Ԡk��7�ArZnz�Pa9f��J�d�@�2 �<uf/Č�A�QR��HeN�1���[-vJ�"�����Z �n�_ʓ�! �4J�fy.-{�Z�.ZA��u��k�O\�^�E7��=r
���}�5�m��\K�2*B�wl��z�Z)6�,�+�W&�b}<��Wa�H�r��|�@����F�͍����dF4Fr%<Ha�!�}�c�r�˅~�8��ih(�������#�V�����k��%�Vr��,��,��d���M���Y� ��Y-mk\RPa�@�����R����a+:�˹)�A01��#ocv���J���&L��AX�J�g�)ǣ��1���5G�!�(���It'u�g����*U�
˚�<mo��>��P&�k���Y�DTGp	��)�l��mPo�ۅ�R�.~T��ɧH��wF#��\)o�i��D���?�V��o�Qyi��fN�0����7���q'�X�R¼�$���܆�ys.j"$"�N��ǔ��Dl����N&�:ULp9Lv0:�WDг�T�6�(�-c����/��2V��h,%���B�����.�(��SG��Q�{g,��T�NPP�*�l��
���GU�H�P��N�%�C��vuB��v�K���?&��.ԍM6���q��fp�)�F�x�.���FÎ�:�����ԟ� iHz��ku��b[��4��L� �1K� �����6:���u�=����!��x��l��8��R�c�#E�kY�E�~W�ji�X����m���B���[*���p3�h�5Ѥ�"�
y���x�"	oYo�gJQ֋�u�]��7ڦm�8�:�^sӱ�����2�r��V����?��%�6u�\�)<��7�����W�J(�o"ߋ[u����y��?�f;�-X� �9�w/<$��	Gƕ);�E�v�-����!����f{�Ú0`��4�`�7������>��o,|W{���nM�[E�M��s�|�z�����]4N-�-����{7���>bH5vo�1����Ufd�b���W��98�#�����C;	<Y9cQl �X�Ln?�����=ۨ����߮�Z?�UB�~��ٷ��ٟW*�C�ӓ�W����Uu��0<GT^�z�3S�a��ډc"'��;`���i�S�Y�Kϻm�KݽI�GA��@􆾣���8�v`Q�TP���h̶�a�XK0'�a�,�O,��d�ܨ�r��ដ����:�73ޟ,���et^ [n��l+��-�gU.:���q�WՀǮc
e@�8~��%h��+��`{�b
U��o�8L~�~"�*��Fmx��K�I+�<vJ3����x��T h	��ɒvu.�~���F��1>�A �r���mRk�����s�FH�b��'��;�=�C.�i�N��]��^���XzO@L�i�ݫ�Q�]�U�2�u��-m�>g��>�
Fc�RS�C���f�e�ɯw�CJ��0����3=E���e���UI[0���'�!��O�սIcɉ�/"3n�gT����/=�p7����ԹK��W@�G\AAαX\�0f���d��v�&���
����Rܓ�`��/���[T�+�tI>�� �.��κN�"���Ȍ�"����ph�[x�̘#�t7�����?��a����^����"h�xt��w���G߽e�d%�r���}������V�Q�ᓺ�`�k�����XLc���	��7�%L!^�~��aR,�;��c܇5��qV=�?��	���ޣ��1��)O*��!�QѭSA�Z��$�I����67_�w�S�5�6��)��\=����ա��E����E�P�aF�x i�{�sĻܲo	��F�h����a��J��?��ba��}F�p3wI)�r "H�YHZ1nF(��"
�P2N��;T)Ju�Px�������-r����j/X-� ��<@(��@����I���v3.b�)�I�+�h �1ʂМC��YY��{�۶;1�[�D�E�P�٢��MЏA��g�f�M1a��ɤ��oӓ�@g�$�{+�r	���b�Cf6u�	��&$����W�J}�rh���H�aS"忼0�:�]�&j�eyz�뛈�K�>>s�x�p��V��l�Y-����%�؉������j�fg=�sv��LNr4X������:o���
��_�1j+%�������� ʲ�_��cl'}9s�bK[�Z�p:6\y'� }�N|\hD�ԑ�q#
�f�]�ISxA�%`�2�VYƴ�-��3��)n&4xu�鞍�9���-*��s�ni��v�N4W�t�`�P٩|;]Ќ�8[Qu ��������U��~�i)A�W�$|C�xJ�и�K�P����|g�c2u��Zp��u�ܼ�ހ�º�<};Y�>�
eN�c�ӓ��C#g�|�W��j����s���F�C��"ep�E��1� �ؒ�Rܭ����D�C�����6ףh�����J�tĸ�"��/��#g��Yܷ��d��5P��k/
Mgy1��?$�A�1��ͽu���%!���*�	��U|$��\n�^K�|��4�/�N4�gQLBw7��sHÈ�kd���FY���zg�Q��۷��D�=�{�ʓ��@�Z}�������퓨�<��%s��/%j��֮�76h����J�1���p5�4\������ZjO��Q$��|	sg����"�oY5I��+;�݀f��I;�5�o����rxM�-�a��)�'�Ɣ<jU�%�D�(�7�������$&y�`�C����'_��vb����4��;��4'Ζ��x}a�vk����0��o[�����͸t���k�_�l��%Vu{�����ML^ryDl�}��8��
	hË	$��&c��2��o��%<��PQ�p�[���
ޫcE�ۤڦlJl���7��"��&���.[��6�Qj�&���r��Rz���
12�V��	�J���_��A��c�+���Ne��^7l�>�&���U�^�T��C-��MA���LIK��D�/k�i�<:7s�_��n+�}Xq�^�Jk~��5�{�{���������^�m�m2=�y!9�j�?Y�tev��7�Amv��.�����\��U@�hV��t͡#�in��f�`�k$V�kחT �vl�r����H*�|���bӥ�8�~�$|_	�&�1��ņI�����{�4{_T���˽;�s�Yo�#0ˮf��-�L)��%������G;������y/O�s+�������7@�:\j��z�����{��F�myR����X�
-�ʌ��z�-@)��?���ir��8����0 ��(5.:�Q�g���
�aK���/��8���ӣ��r.��{j�	����U%��ADQ��s�m����v��;)"$A�h�H��M�-�?d�h���	��Z�*�mT��D�,3J&k+����7�z=C�}���z���j��9O�T�<���)$WEUUߤ!lt�#%��4�5�
�,A�'���Q��C,��(߄�b���CɆ�jȐ����mKԟ��Ŧy�mɡ�6��>A}ב�>�ݰ�8�t��7�>;�%G�-]��NPP�@<8�V�.?@&�j�]OS.DR���iy'�б��(ˡ�-��w��Ԥ8Z>j��t�Sd�Ek��I� �����j��ry�}G�S�����,]kYyvK�����E�f�6��Em��sh�M����pP�R�w|e�D��m�dU�o���OŮ;�B�Q<�tl���9{T��Ū��*We�.3yI���V �(�O^_Gn�q�'�+0﹉�����ߑ�c����@�*8�ʋͮ3�'�1�Ϊf6&���TcN���b�&������ ��S����=C�=��Ւ���ǖ�<'C�(J�8�j�n��]�!��^���*�F�ג��[�^�U2���p��nG���=ۛ>�k���@�@��^�F���pBN�Jֶ�QX���Pi� �u�
��bJT0Ͱ_�9�N����c������>�P����V�������ղ�:Y
�l�;���6�
SV��t�� �S[l����i{p�ө� $��(�d+�������ld��y�*a��rM�4����P�����l�4�1TcӛN1<�B�y��G�~3ƣF�(\g���{��m�ǃ��E.�r�yl�<Z��~	1C߫rZ�k?�PS�a��"���-�������!��Ja�A�iK���+r�Q��~��u#U�uYQ}k{�7?��.�Qٷ�v�wO�g�}�6����%�ܮ�T�@�(硃ً�E��DS���{0�SHi��a����ì�
��!��7�u+g�t�/N��E,��z2䖖-'����R̝�`����S�;+�4�YF�56�CmБ�|/���oT��!����ӕq4j��̋�$��=�a�����d�8�{٩��^�7e������1>��U�'l�8kn
)�7cr��|)�tg�����Sk�h�	�JN�j2����S�9O�6��d����U#)��~� )m@��!fgښiv���Y�{��ۈ��[�܉��̪���p��JGAo���t^^�ݓ	�I�7�ʒ��^Xm'�N\I����l���:�����)`���t�ސ^P�"cJp�h$/��rlD��} ��k���;��8��qm^�"Ъ\9���#��KA��<°�VC�̚���;�Qf�4%S��to�)5}�p0� ѭ@\�xߒ��ި,k'�K����6�ES.�3�o����ez���g���O�L��e��W.�� �`� �qD��pB�}�풳��]<H�X ��-�G�#_��z?��;����Uɂ~�g�;��9e4ژ���nw~׋a�td�Y&o� ��1�-��1C&_B��W���3u4�OuE@'���ז�M��P�8jC��8�˚ �0u�cɜ{�v�BRʳ���|��:s�M�8z���m��wN�%����81�̎W\�Q'6�Ʌ,�ݹ ?��8.M��4�ꥤL��3Q(�UdE4�"N�S��㙦XΆ-���F�	���ë�O�6G�58q�Cϙd���e��Ưn?�n��wk&�PY.�x�o?�p�"Q���B�P�PؑQ|�.�PA�B�l
f���B�}v���jur��NwBo�S����7ЙD�s�s���r1�yNMk����,�@p,�:���A�{������X�y���u������z����b��y���|n��?����6^"+�i�yNWH�Zn�Dd��8\(��F"��@o����o�W���:��Y�s��*�$~::�5H!�)�ey"���������V|��^2�O|V�|^ٶ�6q�8�
����?�[��t�}I7p�n@x��n��e�7t���jSz�/s��s�V/U>c㳖>@�D%�� �4k '��q�����/DK"��*����+q.�D�QuN �=7MϞt�#�h��1\@:����P>MdHO����ۆ����4`�Nd�3�,�8d-����0ï�P��˂�"H�N�Z��;d�[><}�N���W�pE�7#��E$c������wxnZ�p�w1j�l�����w ��Z)L0b�j��7�*�qh�HG����<�./o�^�.�`���Od�э��rR^:��MC�XI0G7�oQ.��Zx`e�,�my{��f��A��a��S�d�}(�б��
�hM'O���1:,�0u4�Pr fa���Hk���N��щ*���&P7�4ώT�����g���F�=e�0�Q6��Vy��ǆ�K"�e��w�SR�T�k��K kH�u�o�5�$c}�[&g'gQ �"���7�<�Lw�7U+�Aܼ�L���M�0�W��ToI1��e>5Ads��a�~;�&g[��S�������%�3헉<�|ku�͑�ӯ�VȠ�����_��󚼄�1䣛�c��#<�G����0�)���D�/e���l	>E{�;�IP��d���P9�n���(ۻ`e�?��& _^'�
~�#-�z�s��[�g�o�VJ�I��ػE�;�glZxi�<=(r�鷔$n��Q֣D ����4����[����D� 0��y��?��[|Qƪ6��S��F�P��N�����m�N�`G��s�z��"���λ)�� s��C����<��6PƑz���M�f'w���Fk�{Wi��M����w�O��,����E�ɋ�*�,c+��ɢ#��an�O�^���� �yº�#�� Y����%�ħ�iۋ�����A��yC�y�eD&M�R%�<L.��*Z�m9!�-���RE��9"e+�aI 0C�����*�\h�\i�k��taRӮ�W��v-�]b�Y��jx�
�p%��k��=�\5}��l�h~��f>Z]h�'
�jn�&��	�Ī���W	薝+϶��� �QB=76�� �z��ؿ=�~��<KVQ�`X�5�J*�~>�Tͷ���OlB\:���i/��S��/�W��%�&(���y����l��2��6-X`���_�m�ёAh1{����!���X�	��)S�y�!���D�y�cM�9��TT��i�q�q��J�(V�'k�3������Hf�����;�V����\��i�-���(�&p����.A�sY��8\'K���ح~C�\���(���V���;� ��2	7φ�p�WԁX�_+��!�����*��ntY���������5�p��R|$6=���q��B�&dJ�&u�
LY�!";k3*�u\>]CNky��LhP�n�1E<1ct�z�f��F���}mM4Q� �L�TܖN�lȈی�V��s�>k�R���:a��T5H؀Q��5/P�aȑ,�
�-P�G�)DXT�����5{`^P9�=�%U�x`�FL��؁�)��s&��uⷹ��P�~{N�_`��Qj��Fm^5*,]�	@k_��s��R[#�Vm�,�(,�]��t� ��&�#�M0�?vZ:ڨN�z��+����ͨ����J\��u;�'�l��@K�5;V�,���bH S�`���U��� e)WV�!��rC��1D�ZÓ�!5���FY%-�� �˄��<�2��f��W2���r9�R>��<�JZ˝')�:YM������i��s�#����G��Xb��l��r'��o��v�wϧ2Dj�2�*b�k�Z��p��Iq��n��)�*�<�1�L�Z�w����12!��<��܂�;^:z�jnI�{"�N��Ek���?����\3Oz���u1�H��pU�Gc"d�F�����Xj�߯�wy�M/?�y�s��N+x��ߩ<���Ok���,��f��XX>����-�f��5��ݔ��2nq"hlZ��~~U�;���+�4T�2��@0������+�o�̺�m7hG������7��nƤ�L} ���I�]��s`A�k��^U펎�n[������?���
��E@$-�~�)��ַ�����u���,���'�6�=�u`d?q�`�J(��`iޝ���
�S�n���m�X���ܓ�j?���U��k>@����̪�3��Į����x�0Y�j�nc;����OH����i���E��';5�j��W���Dh�U6�5�҄�?z�O�}NaW�3r��|Ҹx	&�S�jQ.n*�W����[�c�7�� 였�!�V�`���H
�W,�l�3<��s�0\��!��I�}V��h���QH�J7�w��֩�Nh,�w3(�V@����I��#�t��F����I.�i Fz�Bm�laL���� �ϱY�y��3g�sT� �(	��-YK��?����
h[S�ܡ<|8�3Y����k�Ds�F�����᠞��5B�u�g�ͭ�:y�k�}�ІM�HcĴӿ���4q�.�W'��P�@N���ѹ�8�0�mA5m�i��V~�����[7-�5��.�~��u���KS��u+���M ?v檝{y�X�U��i���C��o��6r���������)p�I��3�D:#2BϺ&�K�]�xT S��\�����	.���M�}�ņEؠ a��G���f��'�K;��������I�[��ʐ��c9��D.Z�Y��{����n���� S���c���"���I����a��ө����d�j�kG�g�M5�4SK���I�t�W ��˪+�K�4��Y�-#7i���49徘/�(��4t�h~f δ/������ɉ-���K.~��q_�L�Bm[�����l��a3+�Mݖ�?�U�蛟}+�0cAm+SF	�3(�A�Y�s8���g��Un<ޒ��Փ!9���$�~ΨCs3�0�͋�����������~�,�}�ޗ�v[���;�ss�#�D-d���Q�մ�i'���=|��O�<{Y�s1���6�4u�[�]�j�����L����#�"�Uo�����e���r�X�rY����g���FW���miڅKa9]���=�����m��"��I��OC�
����ˤ�0��Z�,���7�퇧0[%�qt��>*2'�ToI��L��[���br���E��C�9�~��[��{%'�a��{m9Q���[1L;;�<x�+3#�n��F*��P-���\.���	�S�I;��c.�&��6�����)�]�x<6|b��ܧ�|��!�៚��S�yb����{4�N�ç�b��3=[ڬ�������Y��$
�կ��?�m�������A�����Z��$HzMh�U ��.�ߎx�
�Ba;m�DZ�<��yet%Ɨ{5:q^#ݙ�<=��a��x��?G�s���/1o:����o�'0[��~�I"���$�'qdg&��]�s�]�u�|�50_p���T\�O_ꙶ��܆�q���+�V�ï����+O����X�y��R4��sp�����G�H6��a &�ٱ�@�r_�m��դ����G�0ٙ+9��>3�G�)�;{X4��x~R\�ٕ���q�p�t�ȋ����߮��O�T�t�y��Z��E"_���Qb��Nt��y[�8P���9�{��D�)�w��;=�ѣ�Zkh�$uCo��&ܿH���$����L��tUyh��2z��T��H���K_�����R�h\��&��b�`���.Pf�ڈ�_�v-�o$�����j�+<�w��$CL��m�#h"XT����
�[5r�!∑C�!n�}�%�/��V��@�7Z;�)�i6��K�
J�.�Ojxb�T �/�\.�����2&=E�OZY����`�����3ھ�V[U�;�+g+Ӂ���p�^��B$��1B�n/����l��$�}L��z˺"��0�|p3�W�l��fY����wp�r�4����Qh���+�p0U̸WS�V�S��f��o{bRg�}%���(�k%!����N�wk��h�Y�4"ŅF�X��n$VaS({���(�mm�X+0;zJ9��O��~yʺ V���I0^P��g��X����h��J���rS�/SH��40��`)���P�(sg���cV�O!�/�U_�U�;�!��8V0��w�P���W�������U{S��(�:���ow`�l�<f�k#��MO:Բ��ЂqH����9�X�Ȏ��!4I�B���
~�bN�DҐnt�Q� Rϴa��4�ɴ�f7�ʗ�("�{.c���B��`��4V����PK2	��s���0��~���O#��J���gN&N\�~a���8�G$�}�f�k�շ!��ێ+�2��;`DfR��ky��I�m@>�n��]�$�={`�3�$,;���K^) 2�{(��L���� �5�N�'bj�����.�f�����Gn�\�k/�}6U�x��XJI�C�Yw?����������'ڊK�#(�3�64�_�0Z�J\q���9*(+4 ���A7�Q��!H��	�%y�Y���p���a?l�Uq�4�5�ZT|��m 8�f5z�s�Y��&.p�$���M��nq�,�D����'G��L�I�:m�ƍ�wF������NW�A6b�� ��E�k�z�u�/�;66;*��Q�'���-��Li��dkt�֥C��h�R5�rhS��9U�3u1��z�]*|ď!��suG��l=0�{��6A&m�n�.�Y,n�F�fCk Atϗ��!P𒷀��an�<��J�1%�~B�0�-~�t8��U�I�a#�����ɞ�[t��[nE$��4
$���I�����q���%<?x��,����4���NV粬zg/�d�n!����i�5V��y`%���r��� |']�7��C!��6����9R�#0�zj��p�sq�aB�]��O�n���x��>M3�bhc�!*=sc��S{�鯷=�,�Tt� �P^�� �����ʒ�y���'�=Ɵ|�O ��Q8aȢ`�K���jK�N߆�U��^��r��k��#8�R�hr�D"WR��[�q�L���H$
�m?ݧ�� a��@��;��S�ɳ\�a礜�3#X�x����i/�0@aUYÃWx+W�S���@T��O��8)����w� �w*��k��|k?�󻑊T,�A������8�X�i$�V�[w���f�&鯿x�ək�
�k������ue)`h�ZN�u�qd��@�2�.��Jvn�rׄ������
O��� �P��4Y��{�7�R�c��^��"L��Y�\&K��i�c�N�;JL���f�{�":�(���)toz�b-��_�yN����=��텥�m��Xw�3T�mz� u�e5}2&F��-��4j흓��q�`�#	��46��
��[Y�������;b��-p`a�,m\7�w��~H��i�Ѱ��<4�O��Ĝ4��w9��;tN8�p�I�۱8�5����I����@[ {���8K=�x��̮Wd�n���ed�5�%��~�G�R��C�-�� !��u��m���^�Q�êm�d����C��m�h�b������������E8p"Ɉ)�C�t�m '+��r&`U?��{����G/��=|�wIF�$L� �ey��Z� 8W o�Z�Of��l�e��y�Y��>�Efc"oî��+t�<���}8��߈��&p-tՌ��$��1�-���s��B���8wf��ߞ"~Nrs^K����d�J�[���ꇨVL��j�#&����A*�<h ����HwU,�~Mhbh��Vsi�C�ǚYL�J�G_�#�E|����/�{2�C�CY	cq�gn8NЊ���,�'G�%�x։W]��lj������n'1Ai Ԩ6	IF��ln#�ߢS��xz�0�}�ul�����d�����r!~x��J�)\H+4�Nt@��x��ϊXm����!��R��띌s,�Pܧ�VEXr����� ���؄�_P(� ɐ�KB��A�څ�0��:QR�t�~�"1�c��Ss@b����2��"��+���@�1 �`-c�{ �
��ߥ�Y��.��M^�~������Wr|�Z��!���e}�
�S[�$q�T�� dI���D��	��X);�4�f�)Mh/{l��F�Ef��*r$��wT1H%�93�ʦc֘p��H�+��� ��� �dd����Bm�53�l���4`!���k3����gD� ��u�۱�O�rȭ
��oTV%e�Clr�$Q)'�xzB�P��I�q��?j/����]�:7��cz5'����=���$*��dU�W��E����&T�(-
lu<�q�Ȩ(+�����}Z��ݹyV?C��iڕ*Vgݍ�t�F�K"�KO~���H�"�`-���u[�dX�|,Z/��YX8S�Lq�����]��Ҋ��@�J ��W�9���i6�����X�t�׻����n�#I5�)D�����������5��L|���S��#�� _�%h(�"���[1�����!�+"l�۸��2�Ҩ8b?�g�{� CGĸ؟��4� �{
�ԡR�^�+�Θ$�R|Y������m��1��]���7��W�c:Q1��\K,}�Щ���9��w8�c��(��%Q��ss9�
i�1�� ��WP/����2e �6y`�zGy3��6��^��f�U���&	 �
#=,��L����,�Ʒ�B�O5g���@;� d'�ك������I�ك�t_/P���	k�A
��޾�ܩ����3oh��^ڤ����j�眦n��φ� �f��p��Z5���.����e^��)YC��ef黀�wf�!u�QN[y����\���I
�-����a�[��<P�}/n���0qmGQ�����"������I~I�AH?q[��Q�N�k�����^��IᷩMs�E�1��$m�UQ����dv��)�ŏ��ı��Ȯ�6�T%5fK���&TJ��s��C�];��t��>�
�=��'m�^>��i�B��2�
�-��6x���������C�������M[q	;�Jд?��H�Ⱦ5z����a����*�ݾ��"�!�m���F�Y��u���R�j��0�1:��t4{c�c���ƅ�)�;�M3x����X����q��
�5��wU����D��
g(s,ݎ���(��i���Z�m��%�N1/�E�U�E�P����)�=Z�q���)�W���51͉��������<c��<Ζ��T��g���Y�B1��/�W�G���5��&�T�>1p"��fG4]n��ڵcro�t����:�s�(��B *���MuR��A��6�Ҝ�"^�a1u��Du�ٹ�3�F�sȼ�`{v8Z�#	� 9��٦�`�XC%�O��ݝy懠�d�1a+8u�I#�us�����$�8U�hv|*�LYxX���^�
\L��~��'I��P��E�fX۲H���G�39enWp['��OװN�ŅJ��X����{��Kh������a��X�	h^�m�J��^=M�����:MyV���:l���;P�k�F+��������x�-�P�[��gp�+�4�d�BQ����2�M3�K|c�G�	��h G�L�P`�8d-�����V �
��!�u8�x䊂ӂ�t���[�����tFOoe����s���v�1eP�V-���1�4�xI.�`�7��^VԟE #�F�ߦ|Ff�'����R�L�N}Ӝ�0�7g@�fw�y��r�ݙ��L�GF��@Pr*9v9)�_����o�Ҁ������f�Ǘ��/0 �yًޔ�?������7�
�R����O��J>���rts2�����<��w��dA��W��U:$��e���g?�e�%x�Fչ��ѿ��߽��foA����R�/��@qy���
P�r�/��i��'�	��d�n۴�Ѳ��.��ɍI^])��+q�%�בb~���0�s�7�&gB��2����Ҿ���Xm'3�m���!7��O�0g�(����.Z�_�:X�%IyJ1��/%�:TM�y�B�U��`�R>u�U1˴jT[�@�]��J~bE�d�^��(�Qb�;T�)M����ZM�����` �CC����t(�.�$5���waO{������2^��Yp�ƌg<�q4�ߙ��pQn�/�6[�J�#̉fL���J�rZc48�|w{<��(ʰ	�N�1�>h8O#Ғ���<@��	�e�j�>���Zj��!�I�E���L��9�`��m�0x�d.g�;��<wus�+$�k�= �2���X��?�Kb����P�M�ʹhpg\��q����hW�9
��� _��U���y�� �Ġ��@Fv2�\O-N��^-;E��x��۳�y�7�+'/�ˌO�JQ�
܊Y��(h�)�J���i����(ȱK�u�wd?��4���2��p���v�� a��%?���nE�<D��)vA�ಾd�*�� .Gv�����#_�6���<�7=:�|���P@7�^w& x�.���
��e��8��b1�M��Έd^3����-���;� %0�O>��ԤZ���@�!�u�R���64_
����7^��mÄsM�H����`zg���s��o��Y�5*���@�(Y�EJD˾XU�@Jn��K�t2 *�� �|�������=o}���Dm�ҏ~��ƹRi4���\��hOe4��ѱt�yT�ߔ��P�g��Kb?�p
�lQ�E#��8�28��V�Y�ptY73�sX0��z++��%a�||���Vq�ڬi�EQǆ��ͱE
�N4�4'��=�B.l4���ؐZe|�f,�F�GhT|V��t� q�D<KAW��d��-��+�3���Q�m"�c�&�t.C�g�"�Cj��T֤�e��Y#w�
6.
��E�,+��� ⤭AZBև5� ���1M�[N�ut��@����`�̓��.��!7-��f���py���{� �Z�7�THn�-Y� Q�BxT�c$uI�i��UJ�%��_�N�+f5��nݪ�k����ծ�%Ч��Ș��Z��=�IB�w3�C��Ͽf}�؋��E��"`V�n�Tr��r�y��b�p�5��q~_�#�~g�̠�Ӵ�Q�8I��(���?U"�T}��`0��ԍ��
;ʿM������Z-����FK������Ι�Ƈ��:~�%%ە�:E�}����8Y� ��S��{�M�+Q�H�l)����Z���E����k׆$��nW�7Q���JE��6έΨ�K{�!��^�GAx��v�1+k�˻�����#�_炛��9������~=�K���6x�bF�ݴqSP[�К��V;X�
؅U�R"�1�2$�r��w3'����hst����ఎ���c��y,_�.���ii]���LU�ᇦ?8��fp�M;:�Q��Q�-��!L�;���S��5�P��I��Q1w�Rښa��@�r�P�<�J�v�2`�1ھ�%!��QD������4�O���}�LpZ�����&��xK%����^��rg�3q�;���uÒ� �o{����±g4�a%����ݢٵZ�%3ԙ���zn���}8��0�*@���Y+�qM	���n!�:Zm�Q ��M���nZ:`. �q��9��3�5�*�}G,�5� x� W��29�c��j�B��[ʢ�?��M!V��)��3�9J��u�KvY�{�p @Z	t�B
��rY�o�q�����Ю!�e)��Z ?�+��߁�"7��v���ɾS�iCX�f[b:�y%N�	�h�^�.��|a�<�#/C����������L���	F�!�
;@�k9N+�Iq�/���|s�L�f�מ�~-M��ڕ�WEͺ3�YHw#�j�m�σ4N���W��A�w/���W����R��M�Đ����Z�_�sU(�x I�m��	�|�.��"3�o"y��C3�?0i@ծ�mF|6U��w��&�CNO�&Ƥ8#�1/_N��VQVO�X�C�PW�F�J؆./W��Z|�ޣʓc�x0s��Nx�h?^�G4�X�OJ���s�IڭVP�ZN�"
3n��-y~��I�����h>�`9Ϭ	��kEy�r(:�}U��WGԳ��3�3���I�E���F�|"\�2�
R�'�,���w(���9��EXL�6����y�=N�f頪e#��v�B���ݒ|�v�KB�Mf����U<��O�u(�yj\��Fm���W����]t�=��B�]� Ǡ�],� %�,*�I^\R�1=����]�x]���>f7�SЌoq�\�̆"bH�&z��W3�m\��k��'3b�n[�!VI�MC�š8g&�?�34ӄT�5�=��Z} �L�]���$�*��Uʼ��Q� ɑo$�!="�c.���i �$a�E�8���o.�mնd���].��V���5Z�C7A *�KH�����1�r
��0P	:���Z��-��9����x��	~��e^mA�`�T���A�J��~��m�z���ޙ&z=Zļ:�j�p���˴�3�B�on��&�jtPt;���U�Y�(�r#�lp6�s��Y��)Q��E����χ��P��^:�� yk5cz��ip��e��Ϗo��l�[���?�)�S�W=����:�����m����즠U�#Ϣc)�n��VWh�B&��2p:`��}E�[0, ���_(dY`�w�"兏Z����ͼ�Ң��-��Q�:�S�*�Է���t.
����f�D䣽�.�q#| ���e�~t��OU$m� d<��6jj*�������!Dь�.�E���`ɍ#�@��d��?�z��2w(�j
+�!�f��q��J��֑�Uk
Yr����	_�P�8�|�.���9����B#��J��p� 8��OSF��{Y頏̿�.;J����.��WDo�"ŭ�d2x���A|��?S�L�>؛N�� ן�LGc�W�U������`������@23��i�Ɔ,��X��4���:����o�5�N�KD���U�St>������ ��E��Ay6�)�� \�,���;�Jv�Q;���ۮtҾn�y���v��­+�j�_�0�NWv�^Gk��
e�p��74�����.��To[&o��:��Bl9G�ŧK���s�!U����q�*bS�R���y����3ˮ���Q?Ƭ\:*�d4q��F���ɪ��ͅ�[R��������}��Yk6q����Bу�áz��Cb'�g�y�$]��$��D}����,�a"��f�M�( �6�z��8����Y5��ρ9�8lP�j���΢߷�R,��l(� ���&�&��a��Z�	]z�1������(���������u�!,�g�Ws zv��̖P������@�S���y��GH��R�S�c(�� �A��ۚP�f!-&��I%i!H���=m�AWF�}������d�a��b�<�M��ي�3��r�ȼ��1t�?�,s1.3�̎�jms�?����HD�
��UxKS���k�SOo݃��z�;����T��k)K�RM�^�s��>�6�	
��ܶ���82��h��قzk��1�c�`(&�ɫ_ư��<R�X�X"q1?L{��i�Ҏ�mGHA���>H�ث�I�Z�d��zC��Z{��ڗ��}�ju�W��X�kT���M(�����:g���V-��o��rwGX������=p@d>_�W,`�M���DE"o<W>�9)k�y�@_cz���P��[Mf��"	R�  ���c�t�:�U�s9&����l6��-VT���B�%
�:P�9	����˔�e��OP��Q`0:yYN�h=���� ��9H�G 1��lw��,��FF���|��w�����i�&Pi�{���X H���_�|�{(V���6_Y}فQ�f���Y��% �}�f;u��ÀՊ�;8=�	��|�5&�	M�ϭ����{�DE����N~�}t�w�UGjI�p1 �����C�̱��o'_���*���6
��������Ƭ<�4h�!�!j��( Jxv׍_߽߮ezbIԱs��fo�'絡j˻�}:LE<#�N����Ѡm�Hy�Ք7�1�-��A�H��_@��yUʌ�S����m�~s��lg���c��1��q戟�1HU�w��|c��l���\<�����3H	o��@ڒ���i�4�I��ʭ��&�"[s������].p��ģȎ�1R��������U��8׃ D�W�,<��9��	;[	D�5B����P�;a$�7˯����U�w����R"�*:��DE��Y����,+�h���6�-�� ����Dyл������{��B��������A���C_��6�h�\��m�7?k�|ݱm����� ��"�W�uV�"����>�Pw��Vc����*����'%���	�&[T�-Q�r���_�Q�[��Q���j"-�����.�&��WY��GM1x ,���e�s� 
~�*��T��%�|̊!c<rV��los�	&��=d���<l�Q��T�_	??����R���������)"��mF��+	7N_�����Ä��q�����}��8:�//̆VaG,���<W��aо��|\B��[�[��|�b[���a)w����A?;����@�Pq?\(έP�T�#4�L2Z9ڹA���;k��� L�&Q� �K�:���H�ܿv��d�z��l�� :��Vi(�v\Y�������f���pYIx�I|i��1�<�mc�����?>�}��ν��BM�����9��2W����j㢽�R"�C�I(W����6�[M��ؘ��h_�-ǝm�"k�s�2���"�
���]���Y?�%�`w���	DX��}>�"�a5E�r��B
��*ɒg��Ю��l����.y�(��NT�>�/D���.��!�@j�p��&.���Z��.�~��J O��
�o҉�`�|^Uɍ�D���m/]����1�Rט2��Wr;��hn`Y�׎4a`d%���_�&M��<� F3�8dF��r��-G@:�ch��^��:T9�
�-S�As+�IV sG
�oG��m5�v�rd�_W����x���X3S�mAxV��7=r%��赫��P���"S��Pc�rc��ڳڲ�^��Է�b�\�iC��]���}%9Vtf��s6���a3v��n� ���|�(K�ԋz�~�i�S �̅�#CW|?r�r�U�.�Q��5������D��~"��c7WuS�u]#��tOj4n\��VC�(�&�g�.[Ԣ�zٲ��!Ç''{j<��˾xX��[@]��`�x��y�����������7�^��C�v�(�FFΖ5�W'�6(=��<��E.j���08.*ƶ�g�G�)G�ݤ�]pv�k��5	x�%�R���QY춉P��p�SJ��c������^��I�#z�X��^j�l[�S��?VîȀ<�U�/V]!!��&eq�ש��;H�n�%��>���m*1�~�[Q3,.�0�.�U�v�{�1�¥0o%4���F�6��؞�2V��t���d.��M{�L��.:ꁰ;�k-���˝���CcF_��p���Ú��O��0�4�a�2:��4ֻ��������ᠼY?��~��E�d	�T�|����FS0	R�I��Y�A��b.�E�ʅ��
�����j璘>Aa���ٮ�W�%�r̖�R��Xs<�޺oK�r�SX"v�+�Af�moJ�`/����>�:f��ȉq%��8�6xۤ��+,㻶,|?�A�~n��(}�	#��WtS޽��'�n,�|����/�/!u��}=�^G�&�,!re�Nb�J^BxG��EI�qv�����f��!LL>R�M/V�*?��a�N��>y��=����h� �vK-'�������9�n皸�x�W�3��&�\�eXK��D͏c�襵���9��ŷ	_Nн?�/E\���4��,婌�u�\>4Y��yG��D�"��Ꮗ�f�ݭ@��ڼvM��I.�G�&�n�:F��1/�Ϯtc�ᆄ�~d�!�`UY(l!�xe��t��{�L�s)���k&�������̮�c�:�'k�k���4�O�Y�[S�����OWJF�-��D�oS;�е�䮯/VF�z����˕9n"3;�ц60\b^���X� #�kYA;ho�Ŧ�.7���!��F�=1a��G,��@l+�&����#fH���'�2�л�|]�2�^Ы��\Pm�:!>�4�뽊ğd|��=q�����n�~W�5��!n�/7�7	#--�?�VV���ٶ$�v�c;��KJc�b�E+n7�BD�s�����s�3��D��/gJ���o�c�â�>�&������]fxUn\c}�a8�x����K?�*xCna,
�����PX��.��4I��A���b*n��I���LB^�4�x�p��$�~h��~�B������c�񐻬�߇^������80~#�|�Ζ��wi֢��m+�QIm��P���ׁSoRdc^3�҃j@�.�@ӂ�.��*��g��� ���:��Ny�s4׋<��:et��|w�,j0���f0���(m{ ��@aD�����B��.����	���'��;��p��\B�Nh�e�L�p�����}@ {ohEe��� �ږ�yFNI�=�d/���`��9B�{E��y��/s������M�Xt�e%~_�g�kn�B�M4�־�γ���\�2:V(�Qe��=����q=@�f��1y���]h���˛��#����o���:$��S1�R} o��>/)�B��DJ�K|{�v�z�0H���q�Y��ܣ�j���51�N��Łî9i��&�8kS���_�d[+}~}.�7k9��R]=��36cЈ�,"b��I�Ҷ��M�I#���u}:醵�>�U��Tх��N��	~s�Q\i?5�v�>#
�y�hy�p%rKB�/���_��Ѭ�h���q�ٸ\����'�&��pB�ý�s},��H�E��l�\O#�c�%z��|�M��f;�w�A2l��F.����D|B���t�u�'z\��=W٘͠�K����D���7T�>�A�`�����&��w��� �*�|/D��ƈ���ח~	�I�T}�_��(��Odڠɶ��뷠'$���&Dz8<mB7�2v���rX(���������Y'���Xv  �D._�Kvb�X��_!0��8f,�k	�1
�Op4=r�Uv��F� ���n!�j��4����$�%M������m��Ňo� {�}��T��GV�����E��݇CZ	2Ls!l�)-~�����J�M�G5&�&��n����(���^��b2��/a��`�� ��c�r׊u"�}k[:U �F�r����mzI78e�+���gГ;̃�������[��J��B뾣�j�y�┋�ϊL��
��� ��;ҹ"~��E+i�ۗ�R��V�rq�}��ϸy+r2RSv���L��7K��꒭	�ڥ�r8����V����n�%��^~
照��%�%�!e�pg��?5`��3�~�S��ʽta�D@en. �@FY,���k�|[�n��N�H2�֣&�����qT�j߹�ޡ\�=�
M��|�Ѷ4�Jg��X+BP�qؿA'�5�}��R����"�1F����߶�Qf�`���_�m-��ٻ�kФ-���IdU���j.��Z��ἴ�E���h<�@K��'����e��]�`�Y���� ���"�̺��+kV�)9�Ε�Ex�����2�-�!��m~�0wZ��%9�m���࿅{�lɡz�b1�
]4��	�BM?���q� ���&�u�;E�����@�P����Ė�~�#�'!�1�R6i�r��?zX�7��/����tT"H�AţÑf)�g��OUE�>�6]7]�{fvf,Ī���E]���)f�7P��&���G\���ߵu��NC"�u?�s�h=vwn	���Mm�`֤�xĄ��m���1d!����Wc�(��$A�Ɩ��|�i���/H
���l�R^�V��}��ç�h���yu�}B�' �_��x����6�� ����e�	�f`�5[�;�`4U$GB�C݊k�T��/A{U���j���P|���Y���\�'���vۛi�}s�+�mǅ�K�ASm���Z�uT�>�D��w�ug�\i�N�h�'2���ԄӁ@}���_C%,du��hh�^^��Mm@�_��n\'�;�&<�?���������[/7�:[ӗz���n��s����\��r��n���V!}쭿�ktn�K@�׎`���d&��{~�z*Ħ������,��,	o�����ʿ�?��N��e�A��Xj�q����?5�yH��n�KAc����&.9�ʩ5��p��
\�v.ɛL~^#J؅�,C�#�����@�(<y��rf]j:���$0��V+��bSz�@��v&�{��ttu���H��	�c���Bu��k\X������#o����3����!y��K���[ޏ�Pq`�`|�[���@�Av<:�>D��f��i.�h�K-�
L&.��<����t����V���X�����_e�v���?F���?x��lr^ >'�m\��H�F��A����ݞt��;'Q!����ɗ��-敻Ó3���=z�[�1�uR�޿��	��Ǥ F�-�����6��W��:4NH~�&���n�"�M�Ud�&�����R]�W�{+%�P&7o�Sw�n9Kgf����Z��%J��W}.�}H���d�*��W	�����0l����J-%zw	i�
Pܔp�O`v�	
_>dd��9m;*>K�n)�+ w�*�J���v�Ǉ����@��|��Dɧ!���*��|�և2
ߟ�j�P;lmѯ�s��t�Etۛ ByמZ��4�}u���17B!F�Z��~n�)"�ɾt�
�H�W�7�{2w�V��=�q7�u���@^��r-�%��l���6��̨E5(��D��аW6�E��|P�@��)��:�++�6�z�T��２\]���>���{��/{.)�T�$�Bc��ɍ~I��Ѐ(��a@���#@����۔	����GP�N~a�˩��O��e�\���G���~�"~O�� ����r-s������X>�QѮ���Ӝ�4��j��8��}l�r��k��b�h�r����t�Duu0����&����]|6�Q7�U����AJ@�6��TU�����Dp.��Ĭ��z���/����;֫x8���[�)� ���E�;X�����f1|�ӽ|{�(0�%z5�dE��=7�~�=b(��E�^~S�D0<+;H�����gοwaN����r�qȝ"w��g7#��{��(<��%��Xu4�'Ɨ��Q|�\�����Lwj�Xj(�q��t���x����t�׻j��a$#{�=��-�<d��N���^���J�rΟ�E!���	#>	���F�$Ė�`���_Ov���a������th�`��!Ԯ©ˬ��;���@��'ad�)�����cJ֖��;�'��e��>Qwj�Y��� �jL�R9����1��o#�*4��?AZ�삸��f�[~���Y���_���6XDG��ښ~T�_9*-��������H^���^ ������S�BȲ�m�u8���V/�=���A�Q)��OzQ���"����j��`�`����~��	�|�۬�4D��;TJ	��X�)�*�Z����R�E`�O0����E�/��-?G�(���ta��nj�}��&��O�6XٙБ��ww1B8�=��d��l(����5����Ɇ����(���`y�fK��7�s��4�|[��ﭷ�����.k5�ĬΪ!���K�o)X%2T�{�$Q�\0y6'ebJ�}�2E���_����:̰�^cX�$�ZC6��2g����Xo�v��W=��^�#�@�wX�T. ������q�r�HU�%�8�b��x޻�A�6���?i�<m�6f���HJ�|��8�V��X==���D�nC>X�~-�Lb��b��j��ڹ��=�ם���'W��<~"A���L(V^Q1NM6��W^�mpJ�\���g��R	�<�.��Y�g���'�jȎO!6��C����4��XQ�Ý��E���P�Ji)��"J�4pr��*Y6�dɫC��9b�����[(�����3�H�gX�C�Zo6��� �J�k�m�|la�ڃ���b~jr�����(�y�5>FR�=Cyw���g/S�;���;ѱdґ1Cf5�&y?�b2���ft~%s[v)�ɇ�ƙh�T�*���;'�ڎtYZ��Lr(�����V�C����9>y�U���[4f���S�0��_lj_mw��aF)����?!���5����Jg�r�w�������m�!��B���F.V��P�|_���P�H��?Q�C�7�JVZs_��Ex�_�S��`�lJ8�`-�̰�8�G����������>��"�Y?�)Ǐ�,�1^B�2s1�_���l|�W�o~��V��{	�
��E�TQx�����Z\Yǥ��{�*
��2��Q�� ��&4Q�?���v)'I�3AS^���o��+<ڑm�BۉQ�'%/ʖ�f�Heesd�k��OD���7zW��(CAT2�擋����l�#S��F:;�PP.��ŀ��?�.�7�������$�1G-�|ς��=&�nY�^��4�������z��ݹ�m��z����JK����߬ƨI��#J`��)��X��!�s�]�~U��<���L���~%-oY�e�s��I���TN�.d��	.Kz�� wM���U�-S0ΐi^@7oE;����T*����9;N%��{��>?���v�cW��B=O(�1�iKY��L$h�w�� "����!�)�%Ϟ���/
OV��bmT?�hP;EBz��ہs�LT�ue�2JN8.�-�h�:�~I�����j�@��Ftc�"�|�f	
x��Ў�{E,�{]g6�Q�~��J45�]�{��p�j�R9HW��e��6 �U�u�����E�P O���,����%C[<�Qp��W��{�)̔C_����b��lW'yD'��wI��Z��V�1�}��ʳ��6�b������;Hp�[HZ��Q/��k'�X߻L��4&���XP����?�|�1)���7�:��<��ΈgK����q+H�rբ���8e�����
BB�.��v��ž��hχ VLmL	("��!��9�4�֝�]�Tt���0�W���Ʌ�=���1�V�1�4�޴�����(Bh�))�ѿ�?,|�d��ћ����N �́]���s�~�2��v�yU�ԏ�.�8��^��n5�s��n�cӋ��kJ��qg�:{ח"���������"|�wk�? ��VXn��aP�D������M�=}�S��J�Xޙ:�to*��̐�h�c��zQ 9]�)�;D�dJr~:p��f�X��f���o��g�h���A�[�4Q�9 �:��m�A��!�+fr�StB����)+SQH�h ��������bi��9q�A8�>�5o�$Nɕ|�]?�n�Q�?�۸�L"��2J�#�8��M���0��qig�|��ݤ�}hZՙ}���h�Y�<�Qz���a;�>��^��D�6`6m��); R���W��.�O��U����!0�6��UV�l��i�9.����bm�?�H�ewST��_�#�e>uL	�ʹ`�f�p��}�����8X���!�w���T���X5ݹ��=�m((�bߣ���T�49inĒa�n;���v�3�6�V��b�k��N�~����<�����z�ڌ�C� ���#��s�b|��VI%�.��`�/ �cvQ]��LwH'!Nb,߆2���;XW�ا�#Eي��n��hw���������A"� ��	-Qu����k��[xKKqm,a�'�WaǙ�;�,��0ɼ|E��~ ��I�ؐ\�(�������8ѵ��P��~�sCgt��3:l<�§�|*؆�Ō�|�S��y����ɭ��O�[��� ��ÓQ�/�Ȍ�-X�WO�S+q�f��Dǟk��0|�B�҄�_;OO��ۉa�dM�Eeie)x�UcӓM�M�y��ĥ�)�JAG��"N&�/2-��&w�*����� ˫�Q2D�-5f��`�����]ߍ�'X��Y�����(N.�rc	^k
���	��n�����|����؀��ӘU����0�c�K����+6�Q�ZJ?�mW�y|�~�!���Ԃ��bX������i
����@��3��i�lO������O�ܑ�G�)��9���8]}���� 46�D���������T��g�r�� �I�2N,���t�7hg���vy��R��[ZL�׋U�$AI�l<z%d�$/]o���2 l5ݪi�ծ�^����������g�HaiHxa5\0���?u�Wڞ�ᦇ(E��I����y�/���7yn�t��۶�v�M��4��lZ*��ܶe=���zḓy��u��37�ҤQQ՘gT0�%�2BK�R#[G�
��t�չ�go��8�����˭�c=iR�~���h��p_�o��@�s��a?,j-�2PA�n��M{��o-)f�	M0�Q�{.? $�	\���w)�hky�0�C�{�j��L�YK�k!o�k�S�d���κ�s���?������d]�q8�?G��{<ˍS�'u��Z�}Ղ�[��&".Sl�~�F"��`Ή���B�7Z��d
5�M5f�Y�$m�j[����޷���Wx(��Cf��æ�uj���Z��4z.��o�aL����E��t���mp���-�����̒�<�j���/�96)lp��\�9��� Y��6r�KZ	dkf�Q��җ	��6.��`H��]6Eܕ+�Pz����0T��s�����4H?�qBNo[����D������,v웯�Q7��d���w�a{�8�����I·�0u�ߌ���ڔ���(j�k��r'�7�M��AL	F	m����/�t�_�ƻ"j�PN�a���Y쯻�Bh(�Q�/�׈vrګ����%��9|d�TZ��Մ�ɝD�g���k=���i��C��R���j�=���������g[�P�,���L�i^��,��sZ.��WB�b�An�����,?R%����Zc�f���?I�����_Q�*��a"�1�,)�OC����3_ �jdy� g��nm�m��0�X���C0Hcx.��b�g�rЗ���&1׿f��L��)Ұ�҃���f�e�8 ���m��j�۽m,7�AN��6G���ӱV	>x���\Z\�O���Vr2�j����r�!o�\,�y ��������v�G�A6�"�d]N�%M�]�[;�8J���I���@��/�1o��@a�s���\�����p� ��IwY�>������v�(�+��2����H��b9H#�-���5>��P���NA~��3�GP=�;ϥ6��Z�Ҹ�j���I��4w&0텲��<o\X�>��,�MX�QT���Scp�&Ƥ�|bӔ'�qNB�0�	]��2l�X��6�a�Asb������q/�a+/�B����T53YC�U(�Mp{r��FÈ�R?����-Z@��?��a~AJـ&��'�9�/��]�Eo|?����G��ՍW�}*H�0Ƅ*�Mp���񛐒۠�H!faeD��=�I�^c��wm[����n��6���㔄,���v�� �P^�J�W�%�����_�4 ����80*��+����b�	�ߤr	I���nw�=]�Qכ�S�KR���,��S��TH�%	!�>Z�o����
΢�ʐJ���Y�Fz`�@䧼��>Zh����Ǖ�'��f.J��=��_z|Z���Qo;%�`�:�}G�H!B;!UH��Cr���/R|\�S}��ß�d@�"�X�nb�Ҭ��#fQJ�]
��G��m�m�F�%��db��L\RK���oq���఩��ܞ��g�(�%E�3���^ֻ����}3�/�0Z@�M���W؏юE{������jQ�d;.T-B�L�г�[aI�q)�&�}�᫾m��5�#)g���:^=#lV�6����=�Na�H0��f��y��"�xZ>4��`���?1CY^E�IU2�A��,9v��Ma���t[rM~<��2�q�1Yh�*y���'�&Ɋ�4u�M���{�#�Ͽj ;)����9I\��ꩻ	VAN�|r��v_��7O�>� �ux�`��_�����@̠�i Q����������X𙮽m�(p���h�.�D����:¿��`s��d���A��	*~|��]��RZ��e�}���휔!���%q¦�v�o��:�I�v(������}�rX���`�&��i�i�FPv��xv���)�'�x��H�K�i
;}]�{G�����}V�!2�_�r .�^� ɡ��9�8��o�qeG7jw��
SV��M*K��l��-� :�a��Mʹ���k�����RV�a�ߞ�&FT��X����O�!��>FO�]a�,V�6r�zY���E��l��L)��+U#�0��j��ʂ���!A�m14��j��,�[���)�I�׏ݓ<�[�A���<}u0s�y���R�1���!;݄�Q��$�n�P�6�����ۡ���`�,;��/sߤ��!e�@=�u\Dlmݭ�O���<�P�E6͵��n�PC��������}F��y�?���*o���.���`�?��� �w2"<7��DnW＆$ �9ј��_>�"��+��ps�	���~Ҩi���#�����ډ� �EaEG�G��]�P)�L�d�H�	�E�����Q˿���AeRYE��?
(]bδ(�X	/��7Ey[��V%4���mB&�9a���ŒOw�95b�f�{h���5��_Z���s���/�s;\�j�3�Ht�[9�պ��C�;srK_�p.9c�A���h�i���̄�g�+���l�gm:�Ǧ��������z�1eC�ND�40ZK~P˓�a}����չ[�w��}��=$\���=ǡ��1��z��*ܰ�qb���R��'6���:����[�i�]�"P���$��w{K�2x�3�b=��R����_��T	���Ԝ�����z�����=QY�5#�G��k�=uT�	= �zh�)��u}���j �D ��f���^E�~��u�P<�ȕ
�Ș4�g������ݴ���X��,c@u��zTĺM�cL�$�/�)�&(�?&���$&^�#04d{�I�Y��j�gy������b1�8$����c����Ҁ.T������;{u#6���?L������K�A@���ֆ�����D"�Io�u��*��R�vMc4�ɚu"
@x��/�*�P�HJ}�\�6��C�U�s�iI�Y��Z�YfX�*2jZ�!�4M�2��ɞ�g�x5vK�ș_��'��E̹�3�|�ݾn��{Qߐ�p��ᆧ!�^G����v���l$���h�B1����I�y�90��'��_�"�}w�o�Id�bBM(�S�xP��|;����an3�����UQ�/{[n�(�@@Wqf	L���}eY-8�]hZ�'�M��T�|���a��%��5�ehI���~�2�lA��ڽ�$.n;b����n��س��ޚ,�T��a��Z�8,8��w��4����Q�ZI�j�c,罷�uo��Ԥ��@�����5]&�'>��,��H��򷘂�͍UC�2\rx�%uo��v��Ĭ�om&O_��p�X�Av����l���7*,=Û��B�z��mSx����ܻ~�fG� �T~3qfB#�����>88��"R�:���0�S &DE��{�A�}	�wG�Wp�|Qo�z	����b$9��B�JAS^!��
�@��s�%@�.y}b��-V[�l̀&���š#��[��a0���OC��7P��� �]�=�P�G��d��F�r{�W�9!G��l�@RD}���/aKX�[-^�r��c{�Qj�1�z���Q�T�]��É���_$7��on�I���d�55 ��%�4��SxC�r˳j2[���t�^N����}J��4�)Yt����~�=m^m���eNkR�p��Zo�Q+�gm7�sk:6��{O[yc IS�v*Q�����*r7B�`8\�z�!-��ޙ%^��Ӛم?�[7p��nw}���u��#��-3��k�GI����GX�إ��%ߦ��aw�/��w�C�Ԅ������ӷn�
��ޯ��l<�].T�aI�
�������Lf����}�	9kj�:��{�!]����
_���U@��`G'���d�}HׁP����oR
2�u�=^�� f�!�r<��BO��d	�4�u���%��'��I��C���q��Ю��<��,�Q��؜S*���>&�D���j]���R&y4�f@H�M4�I���5�<,���-�!ȕ����B�QK��^��w���H ����a�{�}�M}�cۀ�w,�dx��Z:��o ���
��vJ���_�� �+A���"�T��I��L��ë!���j�(Ti��g�^�D�kN(}��I6�<̵8l� U	|�_��	�|�$ck֛ځ@t?��1��@�o ��.)�����*��+X �z��.�u�R�W^�Tyn�,�y%c�N՚��ߦ���tN�rRS&1�[�7<����^c�$���:G; v�5���y��[F<t�H�[�L8ѭ;��v�����DJ�c�7�q05��)�ܼ�^b���rI������%b���OR�@B#ﴷ��Mّ��N���!�e�B�mِ�|��:b8�2�."hY�n{�Ճַ�q!\�1�\��#i8�&l��M Wc&�+68M��x)7{���m*=��D|�a	dC}Y��X,v&�+�Ε�~�Q�����1�t���%|��G<�g.K|<z0���S�����+���PL�-rTl��.� ��4�I�a�����{��S��A��t�*ߢ$�dki��C`���ݩ��m V���\��3�H�$��c@{<����gq�����)��~q�U�7_䳾i�͔�O�eDX[~����x44a�[B.O}� �X��O��t5٧���ѡ#�hw=�M�4V�������!�Cg'�w���Ec�/�zA�x��h/CƼ��W1e�1n�A]���Xs=��О�j��1R�!m=��*,�<�t��1�9�N��!����X��I���;�ݳZ�zp$+^L�#ƊDz�Y�e����]͌C�|�:L�O�@=�3V�&o�X�h�䵃V��qfW���f(pns�L�E���`���ehU�F�[�3�"�F��H�o��u��	b�&�����06謅\n8�D�-���}��?U�w4?p��IL��)�wq7�n �	�f��M��0��x��*Q��k%�x��G��;��wXL�7!�n]�S��߈�0G,l��>n�O�:h�j���Zs��bz�'�Y��z����<����� L!�h��װ��w�?/z�8�0
�^���\0a� ��&c?�_��GA�;�8���XƂ��G�w�ςD�cr�3�V�&St\�Bo�7�k��'p;�䓬u/�i��ng��pX7/�V/D����hs`5�`�K�#�Q�1����/M{������鰴�u����P���2Zɨ{�k�T�LC49ZHw���#qi� ��o�L@�o}m��ci
����3/�aZ�&,u��(�Y�gJ��g��(IfG�Uw�d�K=�r�>j�H��]���l��t@�lQtzqݶ��Cy��a��dA;��������+X����1�ȏ�� 3ݭ�e��!K�%HـB� Gp����~��f�ew��"-;�\=6�g�Vm-��R��=�OK�3W=λe���0�ӑEw�wJ4����X�[�3}W���?-[��B�]K�o*EJ$���Gk�iYS��]8����P/~+%�a��pʈ{�ޝ�D�"c�Xj A.��ǧQow�Z �^��������!�$��!8��t`A�[�����>�x�\:����kASo6��/��uo�Sٕ�C�,�c�_5�6��M�y�?je��&���;������"�wI&!e-hy�jJ0U4� 4<%y2լm�'rF.�j]	�t��E�v�/�������3H�S�(E*O�ɂ�쳏gzͥ��"�ע_P!b	����"��/6��&�"��{Y���0�Oi��cz�s�v@D�n�И�����X�aF�Y��o�bud��Ă%�5�kž$��4��Dˋ��ҟ��IƼl����ރ̹"��X��!��Cy�+�1������tϼH���&OFK���1�W�Y���!�"��bf�'�C�Y�i/�Q��ʏxV^}��,��H���)�^\�.UąQ�9�(bf"�v��RJiJ��C��E��&o�@��c�=Q{����Β�8Ĕ��c�r�"�Vz)�R�[��쐱��#���^�=�}��^�xt  z��l���2W�K^���51Y-C]1�� k?���i=�I^(<@m�ba�d}�hRKU0hgK�T�o,�c�%jպ��r�AP�&V��;�ϐ~"f����X\H��f�5%$��sY�4ѱ'�d��}��,	��f\r��KjoK֛2'�:��Y�+�b㍿yuf����,3"��n������i�A4��ZD� L.`=�:��s����V���g��x-�kɩo�V�r��,eK�����gc����P�#O�#aJ���ӫ'?��+OA>� ��5	���c�q�����·.��4]�2����2�HrH��lta�3���Y��lp��9����� h��C	W!S,����lөh�ۻv���n%+bM��*�У_��C2��_�LR��V��9{�p7 �f�����q�_�9*��%5_�K����r�U��
�����!hJ�9�v�=�{Z$0{e���+��B�ϣH��=��*�ge��`����(�BF�E8%���P�i���FƝ���M����Z��;��J+@؟^�5׹�X�U�.7z�t�v����~�	���8�k�A�(z?��k��2`V(
��n��]�?��2=�/��[��Z7���OGm��Ԝ�i�r�e��̼�,h�<J����6�l�;j�%f՜V=н�!��������j�m|��;;�,���-Y���)��Y�i�;��(q$��`Qo[����$�|q����X~?�H�:u����b��p:�euh�k1|�?���/�ɿ!A�J��!�h-Zx������4�V��G���V>b	TJ��C�	{#���3����X��`��t��۠�b� �H�eJ�׽�H��zX_߱�`��}�uh�Y�j?_z�`$`&�-�9>G���*W�S� ӕ��w��J����@�xo^��C�=v� ���m�=T��0�TǕ�at�Ki~Z�ŋ���^��M���w����`]��VL����]��ҙ\�i��������b�����4?�?���
b=Ig��iAY��d��6�
-��ε�� ܟO�>׳�t>��~,�ڥF���z�an�~�.mw�*2�M��5=9�h��_[mx�<��`�Ri%}ľ��|�����=�^�"�TF�Q�T�`Vc�i�g���r�:r�E���+�;�%���i[ԬiEK׌�Y�`_��2��fz(M�t��,u�KNt	_��D
�\��9K��FSM㍂y˻����A��~!������������G#	���:5˝ ���(7'K�4��)�t+ń�9���i`���-�����@ێ�^w�s�u���\�f�o罆�@_�T�2������~�'��f�z�u��@�����S
��{���M��n��xV�?z�}�`Y+����y��k�墼�_v���/�c~:s����{�%��� �=V�©�F�7��;@�6�Im�S��÷Q(_�pL�?}N��$C�#h��Z�G���}>��B���ӌK� ���zsL�/�;u�[p�`{����A=�U�\�2b4�d��{~�f��� ����m�'��PS�>o\�#��:�ݬdv$��!qW�����*�5H�����.}�f��
j �C22؁���;,Տk���.��21�>Hc[���uf0k6'�5��_l��a��<7M6��Ն��p�X�E"��� ���l�h|��<C�PV����P�V��r�o
Xɪ*��l�F	�+�D��&�=Y�:�Rb�\%{�����Г?т�@Y�)	�~�G-3���&�Y��  ׅ>[�;��w@��®8�t�M�Uf��1���	�th#�T3�3ݦ<Kq�J�$��K������_�E�v�x�=���m����8�=�C(&)i�C��z�p�"�#��zK��J._4�[ml�����moyh�Z�?h�3�:�i{�����wC���N���]�S�sM��zN���J�:�
t�q7�#�u�<���}5��k�������A�U��g�������͹�s���ұ����C-N^��6��J^��<}���T�(꒖-y"���������+XX�*q�;]�Z5��Pa)�'Й��+r�t�`iL�tܬa6Wz0z�1W�"x��H������ӎ�9�����&�Ԁ���@j��.BB4��L�i�#g/
])U%f�����L!N9l��{-��9pM*Sb5Ì���:�=R�!����P�.v��
��ݩ�0Q]�sȚ�EtuE�b뛣��В���h�3HŵTy�ܭx�;a�g�{�D���Z8���2w��Ŭ��b�����MT������b�K4��*,{*�(���o.���̺���4��\��xt�[pYa e���n���y;� �N��e'���h��&�_���ΦJ"�Ln�p�V�{֕�
��oxgZ<���V`Pt�ݿ�H�sC��n�4�G����v��M�Ҏ;�-O����8B �닃ڕB�y�g`�۽�q���������pŬbu�Ė�$�9	Օ�(��qZ�?�65ڊg���HD1X/:Mt�O���Y^�\�%RIU��tS�=&�W��|fV{J���.]�.�v�MC�P���#��%�����D�RK��O�^�tTR9
:���U��R��E�e���ޕ4�Y)��<��p˵���,�wE�G���}�&W�%l�L9�������Ǧ���c��$�f�`DahO�a��p� K�4��Q�����?ԡC��J5/�g�8�9����Е��e]e�lUJ�Gĝ��vP
�`��2����K׆]q}�.�V�����z'�+_��ZR2R��+#��Rj�CR��\,hl��q[i�d�}�s�9ǝ�n��T��X�ff�yhgr4���	_2��~k���4ΕM��pW�����Y�����He%�D����i	X��6������y���cH���fM_"¼��,��hQ3��Jls��M�T�ӦRs:̬Wq}_��b+q����BzR���:<��a�JK��!=���!��n�I���$!~U@� �F�nP��\^����S\���TI��B
��`�A��	���N����5,��0׶4�:z��_���U9�GӲۼc��W즜�YeT |j�ź�x���
	p���X�~�N��֮
��ݙ5��p ���bJ+�Yz��}w�A�X�������Ji�RVE-��e>��=���8��v��:��BL�)C�
y���1I��w���m�A�U��T�1+��t]��"��E�J����,�ٍld���'�c��<�nc�G͆[�{/��]�{l�'͖]yt������P}�>1���3��|s�*�Sp��|��0�5����$UN���U�oH��S�>�N52�����f����_�R�$��=�s?է$����}n��� ���Z�ҶO,���w��!R'����'~���:�:�����9���˧��^a�>�m6����\�T��Bf�u�cU�������&E�G�B�6���f?��7��6����� NS���@�ZUY�����'�Ԧ�EMS�+���'by�Ѽ��!��gޟ{"�alF��y��o�V�r�3 �n ���~!
a���ʵ2�!�*��Û����n�e���!w;�F-g1k��B���8�\�E:1�;&��]�Kj���Ӏ��rrՄ��*/l�A-f֪u1B^�օ�AM_߀��bB��!�<ypX6���%d���m"Lg�����|p�/~�Y��u�@N�4d]�с���@-H3'`}�҅��3�RO,�^��a�z۾0xuǙW�̌[����:����ۂ�묯ml��H5ވ�w`p�V�W<�hf�){X>v��[��8<Z��Թ7���{���c�g����^I_>y���c�d	P�sd��	i�mSb���}�U��f������G3���@��,;�bB��9£�	0I�D����T�$ԇ!�
���)z7hB��ZM��o���x�߈_/sX����#u�P��!`�u��V�\��B�Z��S<"���bV :�:R���=��E@���c_���&|Y�˳�U�,�N�GѤ�U�O���n|��'z����[7�0L6!",@�m�_��
���~�'���? �&����I�mM�l9���׺�3b�E�zd��.�tA�ȅ��?GX��o~B���c���ϱ�d�ᖑ����g��èLn��lp��I�5�����o!�<��e��y�<q~�(�;O�Ј��)��|N��pb�[e,͊Yn�1� AR��'���@	h��bVK�b�#����b��@�JĬ��2J�b�v��{(M�D�a7�;�Yd��v��u!�v/0�;O(�)��q�ݩ�i��&ǆN���xsJo����|�f�K�9E�*g8q4LX�o��j4D����x#.�^	�0�`�B"R����(��nL��.+9U�	�P� U�Z���>茖����iT[>yD����
k-��D�e�Y@�9� ��d����S��6��j�Xk-{ҫM�yl��m����]�������VT'\?}�;�Tr�3~���*ǵ���4�
�&C��&��5������߯��o��O:��c0�	35�;�P�� %�g=|��[�fwE�1�ߐ�ɵ8z<�%tsF���<r@�f5Yl{zA�h\h�M#�䓳lבt�NZ�M�܈��UU͠��$��5�~���2�0��Y��ޗ�o���	�8��ڢ`�@�
x���ɾa�SÇn����^J���0�0k�c��8��l�n ���0��u�b�a{?�2S�^��.�)��ޱ�5_�2Q�Ӓ�w]�&�2��#D&�f^n4���YAԕw��<s�+�Q�u�ә Z��-	$�w��E�W�Ay�"�G�y��IP�f�;�v7L�gD�1�j�>����i�r�Ӏ�5O쀱!$���t���7�zr&U�4.͆��HiR�-����V�X��<(q�$s��禕�Z��+a�J��a��?r \�\7xC��0|X���'�
�;�o�p �n|M+:a1v!�t�<4l�~|,Qi�w�(�9�#J� UOK��HD���%)\�Pt��f�]�� ���Y�#M�{�S�$���l�+.��@^X�/0)�3"�(�DD����i���n�A��&2�P�|誏@����w��
 �C�b��y=�=�V��F&A�:2cuh����¯�	/=d�q��&��_�,�	�}WHX���08���7�L�ѩ���N�EǷQ-�BH��; ��������Ҡ~��
m<�8�v�(e���&��{�L�]�ݱ
�EQ|K�ok]�׼�R�f_�*9#Z��߲UGy�8�}�!i�㘫"D���΍7��ݨ(\��K��T���E~�mD�(��?�����W���o9<,ɴ��o�m�G�͙q{1�� �g�}����u5���9Hq��]�n���w������2:��C@�Δ����6�pd�8?z�7�\3���v���<kX�#a"�N�v+w�;u�����f=��B}J�qs`�6:M��q�s9��9�~���R��g�ۯ�n��x�e��E\�cゕ�ٍَ�͑t�p&��� 8�����IP��b����ؕXp	��$��\�����	B��D2�[��Un:��r7d/�ẁ��]��J�}��Ǐ�Wm�r��<�-dk#��U���
5�)���s�g��t8ʣ�s!sy��� �'��,�[�(���6�����ߕ\���_֐�XJ1����o�T�(Q|䙰z�DZ���f1���<����^!#�Q[���
�Sr*�I8�f=��l;���xS�v5��w�.R7f8���B۴z]�yR#Җ�(uW��1P��a��]	,�����d�������_���d���ú��n�)��,R�7�M�P:[��Z�N�|�'�pB�ra?Jo�8�"/?������u��
�[vCd��E����3����.Q#)�JH8n���;S��-�b\�[$R4b(� 5�fI;��^m.�>��a�y�2)P��X�1����Fs{�}�FM�*Bc�}OP��9*�bV�q��0n�?6��29pһ.�鯃��q���8g��f����AT֌L���ƞ��_����i��O��N�N_CٌD|c�j�s�Ԉ�W������L�����7W�^�w�;�E ��7��$0r�-���UJ�{�㓟<'�S�n*�1z�a��l��(�A���@gV��� ��#o�(ԐH��5���}'����n;�E��W��[�*���1=�O�;|̪���;9A�]O��R���I�V����T:�X�u���Y���'i��\'�k'։k���1gUƲ��Jev��4]�k!
����z&��?��՛h�M|e�Փ=�~�����-�ë��&ߩ������ldN�.��YV'g�c	��(�v.�N�UF�P�Ux|oZ���f�u&F �����'�t�8�>��������Į��Vh�o�nq�'��]���>c`�r�su�õ�,��P�
9����\�V�J��&`ྯCA���&]��������9�Y�.L��֑�0�߃��@�G�A�ޑ���@(��w?���XR5OL��w1�v� D��;2�X����G�W�����n�K�[�l9�ʖbר ��<K�4x{.twz����.���ӒqY�΃���Y�j�M�g�?ϡ�Z�d��#�zc#^s����Zw��u���}0s�:>��}-$R:�~����Q�֓@�Q�p���e4K���'X��54���Ex���Ai��������ٙ\�ױs��Y/#��]�fAw�$�P��;8��z�k��"� ~��Pb�m����D�	ݷ��#$D~	�P�H���S�,�I���OXJi�)��2�)���#{��␀�}H�������U��^*��Q�V!��ҏ�Z��"�'1�E_;bx�k�-8�2l���{Cu+.���o=QWY�ȸ(ʾ"��i�y7.t�!a1jMC�U���0��4��7�?%�N;���	m�1R�������O��D�<<��;l�˯��وfޫx��n9v��,��Ύ)(!Hg|TԴܴ�7�޿�9D��jj!�]�"��ǒQ�םb�%m���<�A ������yz&P�	T��
4 ��VG8�)��ޛ��|�Th�akS
�#F6bGb��Pkj'r�+�*c?DDkƍ�d��	�mhs+D-���[]k�)+tI�y]�&l��ǚ]�M��cjE���lyP����#��I������-ø���\�xp���(�fI�"�Y�A˗�d���Ų� �����y�[���(ɪ����Gzs����>��m�ï����L�w�&��. �Z���ha�T��yJa����TԢ涇tt	��fe�u`��SSE�KEكZ�$�F�:"�%�ET�K��[�߅-�|���:f��1\"�I��D2�K/��8֞K����[�Ĺ����lN�Gt�l%_�z�ªi�n�-�lu+�?E!HO%b���B�\�CŒ\O(���]2�1}#��Ý�Rg,�����+)R�m*BĄ��,!�ǃ�~��'#!�Hꤽ�]�5��e�>��`�%gR��G}#r
F
ɝj0|A��e�4V�Л+(��,�#��L��b�� �ߒ�+r��e��t�3~l��@pYIѢ�� ��N&��C���}˱�ߦýIcE`(��;���.�x�`'�Y��*��~WU��
�4�1[%�z� s�J��E|�wf%�1����||f�ɖq@D���������N�zq�~�a	�Ξ��S�?��n�$3+K����)���~�` ��@��cNL@K=|�31�SA
�J�o�GJ.�ֻ}��Q��'�7n��M�~��n8<+�:T� ��/%d�� ��E��Q	:Y_�������W��ڃP�����}�'����t�:֕Ѝ��p��;J�1�3�$~!*���LR�=��
�+R�v����j����sn�!���t�U#:��Bj.�C!�E��7��0�L�װd�{hT��'"�W-�ut�RGܹ�Q�vY�"5�MR�~|��T<���h� �w�}��C���+Q�������#�=�:ֈ�Y�d����Ot�rY
�nw ��[ɧ�����&HB�&�"�tA��/7~n������.W���2k�9��3]�Ŭ�1�2�Da}���������kn�ڛ?ۿ�ҀXuc��������ְ���6�r�|�}iύt{p�u�th�q�0q�8};������48�/F>��6N��ͧf�5�m�[O}�5�CR�<���dw8(4V4c�,%�4�#�P|�O�J�6^�K�P~��j��w�#2촊�Ȑ�C����/l}����ATd�����W�U�Y�w����縐O��~8}0�ar��	����K�.$��`�V��Xc��t��*5&YysU=l�:�����q(5��ꆺz/daч�шͧi�ɧ�Z�v�=�ؑh��JrB�[l���et7�L����>]��>�~8<�S��T�����3��\��I&"=�h���V�����b�#G��1�a�P~�2�Q 
v�Q���2h��ٓ��:�K�#�Y
���=2�G� ��9.6�����q��7"�p�����e���.�'�C��BJ�y�)3�3�"�h��$oj���#)��`"e�2	�L_h����|y.���3�j<;"- �>Ǥ�f�C�LX��1�H5�B�z�?�i����<�g���K���L��U��y�f<�[z�ܞ��2ݹ�ۀ
m�,|$�jFQ�f8�J:����-��,ٗ��Q�k+4�� �[��r�����b�I3��d;y����/�פm�ӧ�d�����*zVX�`v�tm
��EX�1�ѕ`h�E�رl��r�O���Ȏ@*��B��z$�����ⷦ&'��.�aD���$v�6��Y�'��1s�B���:"��e�f�@_���f3��d�g���`2��W+�2����>GO��Ĥ�ro&A듁�!֙��5Go�Ā]��U�����T������~&B�����E�{�,��0�4��[#r���8{�W����0�������� h���w�����`綣��مS%�\��M���Q�c[챘�d��a,�]B%�%�
�R��X��)�V)�b&:u\���Ga�pd:��i�{������!'*bq0/����Xa�� ���@�O9�a�|^/��i/�]Vb-7�W$*dF��	�ߘbW���s���ki�D�t�2J�>���$[�M����}e=�&1	΍K�(b�l�oG��K�������{Py�r�z�BW' u"���W��..]�V.//]���S��i@d��_U�$k��������!�-$?#�@��}� �䗂B_�ŠQ<�6��l��fD�Gn�1���-����|Y.jH�'��+x� �PH8�z�7Ɣ���X������$��P�T.ӡ*tv7an�8�v��`_� ������b�9nR�WC[ UC!��Y���S`��	T��YE�t�8���oX3�_ �Ch��͉�F]�X5�x��/<������`��V�f��`%���wWf\t�i�u�o+o�r_�M��C}�*�������T�5�E #�2uh���6�w&Bw'
��j��:*f 3���Gu���\|��D+��7�\�?��e�����}�W��B��NN�EMNQ4����S(g1�w���.�B����e5[��b��U�Y��E�;�R�