��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<�w��Bk���U��8_�jJ_�#C��'4`C@�k�����V1��U,�Kn,@6 ���|G�v3�O��sy��T�B���MD���xM��؜D����ȸż��?����S��M�?#O9K#{�������ZfsE*�y%��.�i�	���w���~��>��\��c�#H>O�Za(���Ao�?$nx�~�Yf���Ec�`0A�����/���4K��`� �����W��_��g�?�/�U�p�P5wh����l���ZTgyX����k�W�4�,�q� :���k�ǛBd.+��m��	�i�}Ú0>�g-���&�3��Nj&Oy�G��֯;e�ƍ.� *�+�l��h���Φu����|%3IK�-���b����&�|��}��L���V���$v�w��|�n�y?��Om�� M��t���j&m�.��M>�~�ڗUnQ8k�x����i1��N�5zS�w��T���mp�S�d�_}w�G�Ge(-��N���uM�[>0Ԋ��k��̭�A�g�� akm:f�XU\s�6�{X����~k�wU_T� �,�v�ko�߱���ͺ����?nP�+������H�����]�b��ٕ�f�fV۩����'��/�uqC��I�����c�=/]��{�߸ԕ j�))���%��GG�P_�2���(��`�Q����]�4Cq��j����vv�+��?D����>�ݿp�����Hv��hP��U���ͼa;��gX�f�\̕֎W�P�]e��(�Dg��ɒ��
8�|��pbQV�5�%1ߒ�o��}��Ş��D���i���`�����c�&�Ye>�IgyW^����a&a7�����t�g�\�i�'F�J��Nq�����{���
�T<�({G�`l��x��2B��� c�8嵂>��LKd\ $�4�gKp����z�  �*��4���>�5��1~!������"L!/��?�F�:��Z+3ܥf9��H�#�_+/�.m�������pYlx"�m�m�J�pY�3���>�9��U<��ԅ�5b��:7�]�"��C
Ӄ]�����T��wb�M� k �S^ilF^#���Z%�<�������� �S�����KA��)���./s���ۆ^!��-��&�ɗ�=�J0Yk��yb[�"�|%���Xp<��"HH���3!���k�Ĵ�o�UR��x܏+G�`��(��<�X�Z���^�hV���|5�%�ʱf���/Wiһ%���/���|�w�XÎo\��NK
������D��}M�C��UoEԴ�I��,����jO�������j�`1]+�5���6C0�29,xQ�y'W���c��¶`H�%�\t�2^���X[pݓ�eE�MY!��X�!�LǊ���R�?�3��mhW���*�e6��6�\�z	��2����H�v�����Ua�%����A�̆Aʠ���`^�*�t�R|P(kaas��ʮK��z�6���N��62{�l�JDZ�_2y�-�O�~ڿ�k-���n�BG>�{�d��G�<���*�M�f<Єԗv��瀪���N`&���̵u������"�7��[C��VH�d�ȣ�8]�V�!�<>�� &:��\[�@o�é�jܠl�/^��:�t��Gf�%�d(�Y�+]���s�'�Q�$@i �V�ɿ���x��c�ō5�8���.L��?Ho�Nσ�Y�P$9î�6;Ts��FJ�-�%@{�]���:�"�^@��?#���ѯ�ʈ�:����k� ���'}}�q#�3|��eR�\��9�C{w�}�"P6�m,����+�Ν �f�m��(S[�����I.��w�$��zʓ�,�t;��ܹhJ�q���U�=
��l;@7If��)ħmVH�K|�r�s!��H����/����w&���IAY�a�w
B�:4XG4Q����`Ë1|q+�TEy�>��R|*�%Ɣ�^<�IikzasN(�҈��I��޻F���8��^�}�f�r��s{e�(�d��2�
�*�����cN��>��G㘷%�B+�����~��$R2��M��W���^�.��⧦7Ф$���XA���Z�k�[���;_���.= ��n��� 1��6����C<���;�%嘽�g@o�*#��V��&
)���D�@�"H+SlZ��ś��7[Ԙ�mk��K�J�%��Q�&�9Wke�� u�̑��\�#E�s�&\bʁ�g���ZSY��2�i�ƈ�T-ُ�\:z���T�l7��A-�ؤ8��з���Tz�4�=Q1��.^}��+�������(�Z9�A�0�ۘh�Ү_���k���g�Ӡ8t�8HB��%���%��O��v-�{�T�'
bX���c���UCKdZ�f���|����_k�ˏ?Ie����&�+��Ӡ�<$�}����9�"�.P����m9�ƽ9�yɩ[!e�[��I3�mևy w��z)���x"81�����p�g8�Ԝ��XoR��4�I��7K$:Dy�����J��J�|�<C�5a� AR���]�*�e��v$m1hAS��O~�D��Բ�K�H�
�|�}8ߤ<��E�8�X�Vri㒝��3d,9m��'����o��/f[�-�o�f3��K��-IT�k:6�l�{����dɢ�T��E5���0�1d�����3<.�n\��uo�}o�,�	��*A,�yF���pɒlG>�$4����B��Q����(�;�%ҵk�?� V�n6��|�
N�{wvA�tϊ��Z�	�%iE�~	]N� �<ð�p���n�С�]��X�D��mu-ʺ7����S�=�S
V����Jf������a��\T/���r�XL�����B��$�<�4"�ѮO�Xo�t.��We?�����j��k�A�U���1'�H)uj�~y�'�>f�Y�fOԶ	��8&}��jk;�zS��f�C��󎐽X��3��'Ӫ����a;�>��դz���4��P1�}�D��5Ռ-}�0�[uo�J�������3�p%M�-I�`�����W"<�J��'53l�~�r^�,{��I�Z�Z��{2��� ��VFȤ�y��Ao��T"%J��z�#+8>�e:Ҩ2X]�➌b θ�m�B�:`_
�w�h$K~P�]���D�%0�Ta(�X�S����J�h�:�H	��#N]>g�G�q���a�2~��ڵ}	O�����V,)��#�"���c�K{��W�v��_���߾(�/���V�06�(���Z+������V��@?�1�'�����uX��Y�����$ŜBx�9��)�e��3X�W{�y,a�+�Uik'���*��O�'~��t���w:ה����0�\㘆��!��%#�ƮO��W�L�N?ڰ_����˶�,}�jFס�2�����h��:��{�ڞ������=�ϲ�t:;�w�5����ۧ��"j�9��+����1[�
fNșƭx������=�k��vH�ٗ���,�,��ޚ�?�&� �:�?uL��������G��_ߝ1_�1��}{�>od���?�S줘��d��������(�0#�M�wb^j�4o�l���Kj�L�P��8��l�䥧T�{Ű���Fo��ȿ�P�
�� C~�-���]ȧG,,I��0���wb�*eI�^@tY�k�˴�N�ڶ|�[�E1�Ri�6��Q�J�+<y�j��0T����5�uO1���}�T��Ip�0���K%.P��u��*�������J!��D�ߣ_��;U�9��fn�B㠩1��/����" �1��*�i;���x6'�?�"�[C�d�6�^N�����9��һ��ar�^¡��A�2�������`J��5�r����HB�4��t�F�)��� ������ЕG���6�6N�\����듣��l�K���WG�cR`C����v��c�^�6$@)�2~�
�	c2`@��A��_�]��]\X֭�$e����B5��5�dú���L��b�x� �d��"�p��:�;:�N�~���]���Y���~`�8��P��̮�j����NO��/� i�M�`X<6�I�i*򨥣g���-��h+<̼��{��Uޑ��|?傣�	�XL�x-8�&y����q�h}X!�FT��cEK�r���K�_��c��c�PZ��纇���	�f�Z��l~��H��qN��gkPZ5���wP���F[���B��=�n�)�/�qKh���X�X=�͡^{|~ǒ�:�3��]���H6/�T�k2�(���Ʋ��CL�3��%�t�K"�����MHwTL�I�I���U+��؉��q�܎��O�[�
n:������Es_[_'�:�H�# ���m���n�� ��qf��U������8��id���nf}ݏ\|c/�c�Q 0��V &��:o�UO��N�U<��~*���N��9Z]���?�'���A	9g�a܋<�hb�Ͱ�c�2Z�Y�	�K����ڸ�M�\��|���{�S�U���ռS���I�Hin��[���jw2��g��{����o�w�}�8?��8����ϯ_f�&l�M|4,u+)@7j�
�Ut�*� c\5ee��_��"*���S>���B�@�_2p��o�������n�el\�(r�vi4���׈K�}S:���I��T6X����V:G�_>��&�i��Oq(�{��6p���Q�njbCY')�x�Gͦ��b�f�o)�J�Q�F�f��c,"(%��t;���S�b����V����B^Q��8�6�@q��7M��g�U�^��y )����՞f
�O�t>��Hl�
v�p�!��w�/�$��}�*�w�8U��O8�|'��/܍$�lZ��%��ٔQ����t��K̺V�	��#?�WŕVW�Z��e�@�WITW�cC9��]���2�|�������d/����[���[��j\D:�����Gw���ni�:�ן����CD��^���r�" ��T]~:����m��{�I癣)��8i����kk���ޝ��61C�������8o�,�r+�N��Vμ�J��Z ��*�K����C܉\�D21�{c��y��YP�,�N�i�r=��^Y:	���-�.bn�j���~�����e�� ɶ������%�c3���a���z���=m��+p8���~��-g턤��#�G��N���N����Ђ�=6'�y��xfTcl]ä�λa��L&g~��vlޯ��\Hh�����4c��������\������$E����NC�W=q�2 &�7| �u��wT�=@�--�@D��.�U8�A~�@k1�V����Rt!�|�Va�x�7㓉���?i�yG�#��AxMN�˾�-O�����	��X�g�'K�Ԩ[��9* EsDX�4��!"�\�Lt���a�.>�WH�r��UO��k�宐?'TY��`����*x���̍�B�}�?Ykk�۱At��H�������y;u����+ I���tнG��{tL�~�G�l��P�d-�O��d@�7a�읷��m��_1�4�D�نCaOˎ'����(Zڔ-@!���;�����BBzG����ߩP52�|	=���P�*9��=��@���Q��7���dO���*��h�̡���O���=�5�8�rL&����3��%���z��'Z�+��A��R�lq��`cy��"/� D��)��;"��6{#O2F�Tf`�2�q���Tn���Pt�~�Vȡ���K��f%�w�2N6�:7��~	�#f�u��WX��=3d����*d��p3�TW>H.UF85�ȁ���+;K��B�b ��TmU�������Oj��2)"H�վa��i�_'��d�.�������D����`G5UVN�>9�YC�y��HJ��m�6J5xo��0��=�*�y����y!�/�zƷ��Bp9.PEI	JD4pƧ�ӗ��֔b$lM�r�U�R��`�����8��Q
�����y�G|�j\j˃��	��?�?� i
Vqd�"9�m���<m�4�a�p̦��m��b��4e�*e��o��:��gA�O4���va���AOF��b� ��#t���1b��]����Ƣ3�O�����ϛ���P��B��4�O���/�+�=���LK�%���k���(����e<V�|JTPi�i��� �U�Y�8�� A�1!h�O�ր��E��t
��h���@CY͖�B�'��6�i�!���D��˿�O��*˚�a�;�Ǔ�1M'd�w_�1�!���J�V�[�F����$%�oʚ"�M'�ީ��Dc�.�Ǟ���0�4� ����=0�|@
5LÔ���m�d�6�������yl׽p�ݿ
Ȍ�7���6����c��-��c�5���H�-���fǏ�)hG1**u���	RTDZ��qbS�3�܉�E�{+���J�y�h�xO:�x*^e������%�_ PM��A����jAF�}��oi܏r��+�Y%M`q<�4�_��APmQ=����#P4�OJ�!}�UJ��yx90���Ɋ�h�cb��j�/.m`��l��T��N�� ��a�Nޛ]�*�w�1���yL ��N�K^h���o*_9��_=ק�5u6׫�,�å�[�ޜɞ�&7ѰU��.Z��sJqQ�R��	����:����&>h�F�yn[�^fAiD"7�h��[�B�x	��u󳂂�zO��Y�6LQqcEB"%��<r2����d��u�؉??��n+�Fz9��?�rR%�m���퀽��"��u��.������+k�p���j�Fs�"e����^r�h]1 =� ������j��U;M�X��i��L�-g��У-�sL/7vڧLBے_l�J k���4Z���F'ߪ?���?��r?���z��)x�Ax�fK	j恺n���2������2Wy�5Y ҉1�]g[��
|������C5��
3���aL%�d�_d��jQ|A�����������ʌ�v��\)�>Rvr�tڍXo��߀i�XB��)g)�ВȐ��Xd'W֌V*v91��9R�AJ	���K�{F޿�/��l}���ђ�J��\�Ջ�*f+����Hlz�a���/^��c���N�V�+�ޓ�Q�M���@�'�=����� ��"D��O���2�c�� �\�O�i��f��{n2߈�cD1
K�Z�R}�B�Lg��|���M��4(���ٻ�l�C��@
���pP5��4��b_�pZ�0��-p� F���i%hA��J;1��ܼD)�#jP���_7����3��K�c��!���|�/@��F��|��6@ױF��	��j	qJρ~��i�(�Jc��a�H�;u�O�e/�d��Q-�Y�~��I��Q�Z<�V4�m>c1�}f����+866!���2��-��%�e�����M�iLqi�y�C8S�'�>��J���A,�!`ˮ ��*�򲐱j���?�0�GǏ���1��F.���g���z�P��N��Ot��* ��_C��Q/A���D�=���>��_K�4W:��:���{j���D
��0%���'���n\�o�P���r��P��B�o&� �T�|�
�;����8����ti 4�fe�~}yTQ`i���p��p�T�5�pQ���d�k%��:%�,�����o��o�1�¥�q3�6s5��d��lb�_ ��tԊ�sƑ
k6�(�����vT�z�71`ȅ����:3�]�m��N���q�M�u@��wX<K=-��|�C!ϓ[�z���T�*���7�F'fzػ�Ø���U��FWK��OK���P0���9��>�pOz��!�����H��ӊ�l�5�5H �=/i�ڛw2OѤA-�,ټt� Y�q��ڏ�(�T�KE��������x����%rjj�R���S�?d]�X������@m��2%i0�w����\�@� �r���*BZ2RbwT��4�-~�G�/{�b��C(R(�5.�A%l�?��G�L^�xj��H��'�v�!3�������&�q��L��<ڲx�.'1���u����<V��(���5�mn�)��$ 8��2�.l]�1�#�*����!�~��8מ�*���h�opZց`�p��c�]*6��$
W�[����=~$��aʹ�~q89��Z�u�l'�
D�W|�(4k����Լ����3ut�wV��M�j1͸>�Roؾu��JW�
M���L΋W2�������3����QB�#���D�A�nk|�r�^0Ԃ�ھ�t��d/t�=��@���2�C\ ��u~��nx�.�^D��lb�bWM��͇�{Ծ��M�x�(��٣\]�hJ�S�m�m����f�*Ƌ��Z5��AH��q^k�����p�:�	,�_�Occ������Q�&fwo�[dף�G�iB�G�L�i�Kh���ħ����VN-�Y�\�t{NEn�я�+��uJ&o��ٌ��).W�@<]�Q%0��&��1P�a�	�D2z���!��
gהeq�Y�z���z&
5������D�C=0�7X��5��g@ǻ�ܺM��mGkR��P����N��;
�U(J���=��4�m�K~�A8V�ns�W��*����Hx�v��S嶯זKE��?hr<�#6rX-�k=��,,,��m~އ>~����Ne)��"�&=�X��m{w[m�9�"!W9'��Pi�d�EnP��
�q4��5�cl�v�a��,��1��ut˚8�Ic29�A����H�*8��;�s m�).�@�@[-�[|