��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�8k�)9�k���J�f ۘEN�R��>�Ug:�&�1�X�,l�v�E�%bm��̅C�bo�g,�A$��3��J��X �V���V�mR.�Σ(X+��0֢�9�p{$��ʚ��|��7���E>���ƑF���c�0��x�L\f����&n�\�ϴ3���T�K��yI��	kh^>#=�˺Z�}��4�L@�&x�g�J��]�1�n����hН���1��^ yl�Mg:	J4K��_6�u�īe��x���[�nfEUR@덡�g$=)��Y�d
�-$� ���'�VN�n��T
.��a�N%0�~�o l�cM�6�a�X0}�����!�1�o[��n��_X�dAV��7m�]TN�$����b�%��ɕ��G�q��e��߉��8��A$zE4J�6@0 *G�m ��"8���
-�����.�sDs2��i�vNߺ���7�,�������\\�e3
$�d8�<⊉㍊l�ų$����*���옔&qQ�����"5L ��ݣ=A�u��9B8�;mW���𯿅�1FR�
G�*>
�Q5 e/ё����q��*Hd�U���(q�_�
BҊhf ǎ�r��<�G���C�|�3��^D�px�{��>#����k� e�/��/X�t ��qr�"��Z�W[��pJ�������^{C�dj4�k�I�����_'��0�V��\��7"�\����ͫ'ў��>�kX1��X�}kMV���%�=e�'�k���~�Nx�~�������M^����A-���Z�gaI��q�R��G���C�~�$�O�p��!���G4Ģ$�˼|��B�Q�y>U��D�l�e��lÂ�����~A��S̳��W(�]�����k�P�E(fO-G٬���g��S���gnj0ȳMB�8�#]��U]����'��>W��������ի�o�����]�Tu���EJ��{xP��eF ]�^�8��.)�7aM����^�)lj�q'0�:�H�4��/B@�w��p^��u��������ʪ����%�}��H������ӪIU�$�����kn64��1S�[��A�W��)`�!Ի!��YXz`]<}�}e���R¤��{㐾�ղ�>����xD���֮�7���_���u��6�3��_Cy�w�X���UE��e*=�ɳ��6	
�*�/�y���hϮ4r�]�]M�mGɖ��pZK�����������*�7��ڟ�θa�?#�!���k2�^��Ob�{�C���GDD�`�?��zbw�&�k �>_�E	T���O�X5k�d������}|ږ=f�ЌDW���7��p�R�T��5njhO7?�]�k�*��Q�ζ~�k q��X�XqTX��y�
���U�`�ч��U��Ҁ�p����oT�n ��׻�뱱ټ96��VB��'���U�_��ɣf�t �D��V�Å����\9d�aqHY!Q���a'4V�6xv������} �w�\�Vn���\;�G�&A��|��Z`Ĥ0y�F�]ȑ� '�\`j�6S��.�z
�	��Mu$!o�Y}���&o�m��6gy����{�@!
�A�
]_�m*9���a�"�Jbƞ��	�B�Eƞ3[���q&��!%�ӣx]\�@�[�ؖ� �i�a9�"���-�_6��ةӧK����o���y=��p䲭�8�� �K�&X��!,��1_E(��pP�{?���O_:�IχA}_�rCf�1UE�����EVE�E{yj��	�G�7$�e��B0����Ow?7e\<�^s��3U�I�Z��j�8 %f���1 �V���*G5���k���9�\f{ңՑ"�l�Հ(���q�'�%�S�ۤ9�أ�[U��$=�&Q1�K���#\��uo?T�o����@� F�����.�����"�t';��@u 0؁��x�Y+��\DRy`�N;*ѳcAk����sp変�քߣ���$�{�HR�����5�*̪�46sQ@�\W�=b�}i�֑i2����Kհ�ذ���P�s�����'>�o������o5��Йq��,�`!��9��q���¨C��ھ3y�{��o*��_����ڢ�> �X,Qyi�����-���6�i��߱�B���I��I�UQ������w�d�=���Hz�lO]�E��4ȝrg�É	h����ʇ�~����-�d��R�Sű��6T.�<�[@��,;"m}�R%	���pnB���nW��7��y�����G�в��A�(�?��}�Х��l��7�Fu�Q.���li�?xSI�b�2iN����^�o'⁡��Lǡ|+oK�A6�a�� �Ң�@��#�'�3j�\E
'��D����Ő⓶ʂP�]�QX�_�큓�����n?�Y���3�	p�*~��(����!��*]�����찛�fn�'���@���X\�6�;���w"U��^�VU�ѝr��ǁҵ��P
h�Wyq�N������ך�� T>�����Iʝ"�5%"�����_�[�p9d�>���+~�t�R��=@�"�\�'Hf�ǐ�zQD�X��/�-�ȍs	���h�^�E�AA�?ӫ&Rg�P��do9��r#"?�r�w�dn ._��k<�>�$�<Y:���t֟�}�2H6�3�z}/�(s):�X��9΂��-Y��[�|cpѻF���\;����U��b�)D<BV�)T3�e P���� :����޳�m�&������Y��m�Ƅ�F�0�-@製�TF���d�[.�DP`�(�_Z��C+��N�l�ES>�����RF�.�}g�Z���9B%����Ե�1��zm�'jn&<}n�Ƈ}��{�)��=酚%�<Ņ�5o>[غ��UA;���ʍǟ+xV}/R��OI���`��Դ���,Г��;k��X�b���@Al�/�L'�q��d��G�E�#j�[�@��P���䮏V�CcDrрg�'\��n�7�ao�d��Xkq㒐��B�f��b}'��ئ7��@�{���H4�|��g]�<������\�7J��!��l�B�R�`�~�Q�-�Bc�3��w#T5���1¼G�E��H�I�����\*6=!������+�Hb@[Wq�e�lBO���Y�4ɲ<+�m5q��d�j�XN5V-��J�AU��J�>�	ZM9=�����9���̰�ꠜ`��7����_�X�\�u9|��]	.ؼ}jSXw� vؑx��"�{�����n�ވU�]�.�P#�"&���^×�e��W����q8q�����i#����j���NS���#�
��q�'��ȷ�����p{bo<׶ӛG)����xpn�F0�����D	�H#C���W��p�>��54O4� v�����q�-p���#�m���\�B��_g<����������e���vr����C>�x�O���<Xi:�r�f�ۛ�c�P��$����n:%h�S5n_W;�)����i�5�=��pP���Cs��h��~��6�ٮVD��%c��:Oq��A�ؙ�ޕթ�D�6y
��ȵu�F�ޤK��oߞ��L׋����P�D�;�AP�q3��}��c��s6DJ�LB�Z���ң��M��sʹ&�d��!��;�U<�N��M�5sPa7��a�wGn�{��U�<�G52�� ��(���1*�SJrQ_t��sƒS�O�{������k�l���.��W}�SB�%A���wE�/XS��X��T3lDѱ�x$7�zPV�X��QQb�8V�XTT�dT�N#Z;_�g}���ڲ�X��M0���?R��^�L�/���������^<�_��U�W�>�ۤS�m�3���.f��kC��%Fec�^�8��Sd.Dz]�j+�ʝ&��)�
�����řP��i/��z���Z��,s�%���=]�n��'�^^�?r�s�+��/y[�L�[O�\СɌ|O�w�Ya��&�R���YIVOi�ե
�$Q��Ƙ��M��l��QH2�^��FZ��3��\��$5�����HP�+��%��Q��Ж9q���Bf	1�}eeG����)�.$TR��6n��d�{��$�%@fNy�u��F������C�*��l���CA�o� ��t���W�i���a�3`�`dD�o
��0�P��$��Y)?��9�M�? �O��Tע��|���Jɗ����U�qK;L�	�	%��Y5�Kqy�w	}C���*�ya����̃&�P��5Ŷ~���I����� �h�XI�+�O6�'Aп���a�����Q��r����N��c����} ~�nW-Y5	�j�W:�wTwi�<U+��`e��I�n��a�\�G�,��9� A �����H) �T>kp�Pu�6�4PX����>=�(�+�C�Vё?]�����#¢}���Y�Q�w�������N?�Y0�:���
n�/��**κNG]�j�yCqAA��v��ϰ,�4�e���ƫ�o}b�G�șD���U����f��މp�]Ay{Y���/�[��݅���?	^v�[�u������e��j(K���FF'02��wR ���̊_��.!�,��>���=�R6+�p��4����[{�C�Tpf�B�߄�8,y�8�e�W7�8k\��O
5q�^�3p�L�-��#`���arK3r��%N���	|�cy
��_��Q��#K�(�E��N������m�=h�M|�s�n4����<H���
�3��ÊD�V�*��j��s(���,�*e�S�k�C����Ai�C��.�1[uC"�،�
�H�w�h��
64�Q��c~_4T�R�:�t.ci�[�U��¹��SP���������o���[���ik�D2��V�~;bg��BY@j�ƨڷ����@�K9`0V�'����D�w]���T(��!s���Mk�q��:n[��n���K(�z`�ډ#<ȐݲhQb!@�>:�ĩ�kGtӣ��z'���e �>�͑�Jn�T/�u��*n���f�<���������3@�����KI��E��>"�	�q|{@���<��uC@��������V��ܠ����D�/Y��&Ž��~[����a�%�h�?2��0u�@����S� �j���f��bm�=Ӷ��3�;�4�ߌ�ex�EjW�@ܢ�x C� h��P�U��rU'�7���z�B�Κ�s�L�@��=���3C��wJA�-�*�*t_����5׭�$A�j������ŧ�F^[sN�G�S�iLɱn��{D�k�鿹��1Ґ70��/(����k �@�gx��.z�G3x����)�|��]�e�7����ȃQ�h�����r[��I�xL��$N�'9��� �K���929Y:ƞᯍ��w��T�R'v�\6�л�XĀ�`��>:y��*�	M�<��ŕ�����L]�T%��xM%������1z~�D�ǎ<6|��|4[��^�0�_'wN	̏���T�s�D�Q�P�x�[s
E�2�D�$��n�'��K�O��mE�Sؗ坎�}R��`��,�<3��@аs��,�}~B�ǰ1Z���j�	��(ǵ<;Z�Qd�Ck����Wnvr7,;�*ʅ($�8C=�[���=�Ү�N�'������o��ʷ�]��A�w��W����0N$(U���K�<N_.[w�a�z�����_zR9�C�j[��J}�]��ʿx�.;�|�xvu1O5nB,��t��cS�A��v���H�f���jf��B���wo�"�d��Z����`�BB��6�Ox+G��o�c>�)b{��M8sz�5̝���Q�2��w\�@ڕAj��8z�A�R�C*�Cl��F$�8��'�Ϟ�fXK�(Q>1����͆���D1Sa���>�����.�7�U>S�	 �t�No�~���gPwT.{Qy�jX�^m�]׵��5?.{��E�[v�Q�2i�Q�	<��s$��̡����o��E�Yk\�r@��3� �"􉆙�"n��a��������f~��w�_��Y�5]vͰq<����p��U��PD2�-�E�;o>�v?�|Ŏ��j߻A�_��y��Ԉ���}�ŧ� bC�a~)'���+׮���v���BPX˳��UYl�4��&����_IVZ�k�$�[q{�7�������q�F�ב��Ĩ���I5�`�'k~��@����7�C��f2y�x�¡� �O�f�S|�����N��Q�����k��iZ��u�UN�?ئ-��?}����R�mk��:3-�V���z�2��: �D	���=�zX�TO���L�q��"�r�P~KM yD��G�g$��ʎ&�4j��>>	���
u3=s�@G�G9����1�F� ��;V`F��Z8W�?�{�]�gQ-0��٫<��v�����ﰒ� ��(�۔ir���6 �6�Ϊ|m���������i�(�;����-�"!%LDGx��H��1�����X+�[�ܫ�����YV6�s���R����{�
��N����C����qD1JJ��.�lcfWw�fֺX��Щ�f5�mt�4[�{��]z�eo���Җ2�n�*�g�B��<)[C(��9���P����<*m��A�~黛E4�N�����ϥ8�L���2	6� �0%�/f,�uV,i�C����M�����9��S̄���V��v�)�Q�z��9:��fpf^�~5?�>���v�^!H�"�}��k�<����aq*㑿�Cx-?pW���2P��`Y.����7t&�Z򥇕����7v瘤�U��{�5-%V���Z�KE��ĕe{5�K������s����kEn�G	�������3Id�rG������u`�^�(����wz'�I����ɝ��m�Ϸ�	�Gu�6�3B���^�!�e�e��w��	�e�X�n���$7�?v�r��؉����M�#O���s�(�2�����P��o\�;�Ħx*C�}��G��Ɵ�ç�O}SQ���P���� +�a$�?v���4��=�v,�-T��p֨5ݮ�ru"���79b�F����rx<ēZm%�2�U��CN��n F%���:Op�+n����`=�Sd�5�n�"�9{���aiB�</>z��B�+�(%��'6+���RŬ��q!�[}����{k{z^�"�3t�Ѳ<J���b�,W���/^�~�f�Oи�UmN�qh74�)��s&u��K���43e����MP�9zO����Z�K'kE�j		E��
RLn�j�f8�3�p��qq�T��Ae�0o��\���D�_���w���	ଇ�,�Y:�,f5��W2o#M�<�6�w6l��5/�V��"�"oV�~�`Z��E��HM�Q�yܞE6p5.�
�,jK �A��x�]Uu�	*%E~���S@��Ro=��Tn0�~�!�d*n/�76�g�I�4��"��	uv~<�7B1:���sτUPN	����p\ˢ�z6gf��ȿ����CLz��qCwLX��g�O�ɊQ�ěb)vRLA������ �Δ�O����^�����ͩCAct�ϛױI�zn|�Sj)��4���z"�Y�Op;����pT�ȪLLh��*��3���|�8
o��{IUI��1�������*�Nr�J��4��Q.���,ڮ�+�Qw��~!����##l��^��u�����ȱ)K�S���?�bns~��	������oKO��w�7S� �t3���B&��3j�v���_ ��f�:�ɱu�+;���lʾĽ�X���3��VG�jS#��l��n�����@$�Qݝ�Ϸ��'�s�}t'�'��k���N�4���:�!�j�Z,�n	rq��M2�tp^WtF� 2J� �UN����)�pƐURvT��2r�RtD&��Y�����v˃Z8~K��FlC-��lku����`��e7�v�9�P�P�ry2�N?-����W|��p H��R��ǧa�4h2 ~���W{m��4�b�>|�X	�鿷ض��2��L�V�g����L���a\�?~.Z�A��U4��)��M(��dhT�f��Ȗ���X�}��;�A`������2��w�5�
�2�ŀ0J]J��	9��I		���y�����	�SĈ���uf�(���D��g
�Hٽ�K�Ss^ݬ�6c��_�|K�K��B��k�Ȗl�g-.��
�lh}��9������4���9!��Y��M#&�j�i��WEq��@��
���B�`}�3��
�0�������A\A�}��A�󯐍�Y�d^N���>T�g����8ϣ�=��HN2A�\����~D������}:<����˹=��dr���x{u�r�g��O(��?�&TT�3 X�iYvE쩓%&A��"zM)�d(��j��P�j��E)ޔ�ҏ�ј�5ц)�I�>t#B1ϷyL�� ;"����~�:��6���\%�`DԂ�Z1�� �N�^��8�Qt��R���3w��7z�z��>�c�>�GP :/������B��S'tXK=��S����!�"h��"�	<3��Ф�y�]sҥfx�CZ�^ԫ�J���LT ju�{��Ԋ_=.�7�9Ɖ�+��/鞷#_t�T�O��U��������7���w�Xo]�o���l<l8p2Zz���8RX�H{C)s��OȮ���U1� ��Ӆ b{�j{��/̡i"X��L#s��F�jg��2�h�oS*/q���*D�؂f^���*'���Z=�Ŏ�	����>��L����+���%,�a ��c.��;E�@|�ʙ�F�Ə��p�Y;N�e �ɏ
�1ʗ�&��j�)����񁇶7���1>43�m[솫'Ԡ���:z��������<AA��QU�u\�.	�<�o�Mu��e�+�������|OI:�x~oF��������I�	zCא�����WK�p\<�՚�6�a֝
o�>h���6B �\�
K{T�@j;������&�}���X�Ew[���@�<c�q�>L��l���������7�:�\�$���xjlE���ꊱ�ో:�2L@G�Uf9Փ�5ː2�R��2^k.0bq��f�����=1�Tz�ASQ4���V?Ui�xe �$
<����k����
�4`��r�&�@� a�H�5�>��>s&�嫬�rP�l�y2ku�SKU"�B�3�m���ǃ١!�hIİ����P��Bf`צ��/ȬJp�oNO��~���c�<9ЎUd����M�5"�,�m�p3Ǌ��O?���L7�B��[.��'h:sH-����Ɵ���d�Tq6 �'��L	Hv�]�~H�t%�ɞ{�8^.p���ʡ��$�٤��_ϛ��f���s�dշ�mfST.�m�7�#V[��XBۙ�����f��k�hd�-%H���l˴A$S�H�V(	bc۱ E�c�� ����!�˗tO�8�Vsu�O�d���X�'����%�dD�2�_7+������PG�Lf{S�6L"Y����C#wf�\LN�w�������{�)���9�B(Eg��I��IU�+H充��#p7��Iv�:�8��~��+Ҫ�}V�JPº�5���7gz ��E����G#�=���cÙ%�����(��?C��-��G`&�-����I�L%���͋��K�����U�*���9ͶOW���4|�ƍx@�k��8$J�*w,n�
v_E0E�1T�K5��eOܸvɱ����v��8���v+��o��'��_0��j�G�D��ܸ���rK�'d�� �N-�ʷ٥�L�G"LqKt���X���٧B"��C�r��S*�4){�z�����}�=��0�G� ��M�;���3���<��&�x��r�[k~6���y%9Be���'%�H�^}�O��m\�$DL�-�Ts���Ȳ
-�k+��Qc�	ఏ�e��?�Г|�ϕ�f
�	'�ω��7I�^hj��-ҫ��o��W���!\z�t"˩�0Ij��^f*A��v(z���+�\W_-%��6z+'E�U��6�m��g�;/&�W�/�~���N:>`����k/9����Xi���?�!�9&�6��	`t�COO���eq4��|��S���˸؂���,���G���{u>f�~X��^�e��������A�2�Z��
����{̷m��\f��g֔>`�s�V���r�\8?�`7W����;˶��b�K~1?��؊n��!ȃp�'�e{��y��J��6�Ռ�D�4�i7��I�O��AV��Ƭ����{iu�u�W�C�nd���|�4c��#���;��k�I��B�)������$�pW��~��ݎ��üv�ޔ&�¼�p3��$��H ♫��1=�D��r������&5`D�v�z�vݗ2��R$�f�gJU�����:%���+�����,/4M�ޢ?�n����#��� A�v?߀3�D[*u�Hb N�1���P��[�g�	�߳�;N�%�W�@`"�K��B�=�� �+8�OT�\��J�����X��tz�֊� ��b�=,t����	>�M��Շ�UV�Hԃz���J�Wo����&�>��G!$͜J�Yg����Db\�?0o��7�	���G����̧�0����0Ѵ��M-k�Ǧ��8��{�j\Y᲌��+��]к�b3�.����Z��e�[��S��0��-xk8��I��B��՞� ��'YI��ۯ�����_}�wN�n� /�����O�Q,��ɽ���Y���т�|��Ȫ`�=��a���{�G��(bS=�x�3������"��:^JܕMgܭo���-�4�x��)�t5"@���·��<^�r���S��_�4���7�w1ZHé�F�A����}%���lw��N��o��=ҟ��Q0U*_���e��}��_hpJPb̝�p���~�f}C�������Um�o�ۘ�J�R��t��5�K�1�[+o�z%O�ݞ6�{ƥ���	@z��oB(�IIu�aH�2YtC3�e���vs��u!�B*�BU��L󅍀������=��UD(���1�U��h����H ��K��܁��Y����Җ�lp���x�ӝ��;��~�{��U���8U1ʢL�6�B���ۉ��ʓ�h*��{�9b¡p��9�ޡ ;�#$��y��3�
�uwa�P2����B[�����\�7�U�ߡ�v�<�7�6(>�:�[ˇ�j��qcF�ɴeМ�R3iZ�G��t)�ٝ��D���>�ޏ�Vy=UK[��Rԟ��s���*��]o�}&:�wY}��s*#i��uB�l��&y��؏(�X��i�A�ҭ��sl_n��������ltB��wd_d������Wr�����ĤI �����2�:ซH*x۰�Z[IJ��|S��������#KN������7",��[^J�#�F-���b?$$��gh���=�Ĺ�,[Q��_�awQ�I����TD��唭�6��"�j���fϕ���A�Eٯ�Rϙ?���<���
|�Ĵ
Q�9Ko�3o�ZV�K5�5��Ƙ'�S�O���E�oL�""��a>R7���Wj� ^n�a0�U������M%�\|��ge?�c�VsJ�Һ� ���~2�ĩAI������1^�ߒ��~i�����^�@�#�p�\��!��:�=�g�!��3@MyING�c�j�+�$r�ܟ�[r�zE�_�鶯�K �|n,���jU��
�����=�_��m�|B��rR|?����h�*�GQ��^]���7��@���f*���l+3�TY�#d��q�'N߹�	O�~HCO�_�j~Q�ŋ�.|񚞤O��V硿�p�"��vfEq�?��y��3��c.	������UKK\��J��s�<n�9�&Fbrme�fi�b��
� ����U�r��O�*Ҍ11'W�uϓ[#c>��⥀)���s�4P����vħ�߃K�MO���/��:�@��D�)*e�>�,30�yP��6]]-z��jw�|d�/���P�4�F��J+g�
5P�Ҙ�o�����h.�����sG��M�Mv�(�q���8
���J� ጎ)ӔM�G
7=h(9KWLgHj[6�7�^����$� �����hV/?	 ��xmu�:qY�� ]Pż�Hw)���~��W��7Sj��7������ Ä�2%�� QR=}��N�pOS:�DF�)�oC�X�-ۡ�͹�BpR�O*,�J �d][��#F � ���ƥ���\�I�kjij<U��Y��CX��*1��&��;=D��*5�+����C>
X@0q����)Tlp|z�B�W�`�b�O���rZ���Un�a�c����-��>�"�Fe�;h26��y\��w6n��CEoG2�Q4��3�[=i���$�,Tb\qOP~ʲ�l
���8�x��.~!���lWq_/Y�@�{�}���~T.��t�كIflc}�0m�	V��-N�<~^�~������A!V-���[�:�&s\r0�@�49�TuK���V�
����@���������Sƽ7�y�16�<@�w�P��s��8s������Ԟ6�t:t1\OT�Z�f�Gר�-W�t&MLH�z����_W �ÿ�$�m����:)ly���k�����b��c���)f&Ǟ-��y5E�p�q+69Al\�c�����^�>�)Oa��=��*��6V���Jd���Y��*TS��ZonK��?�@[J$��WoͼP�p��ۇ���s�'�X+&8,��$	�5���w�� ňl *z!�*S���G�:�5�b!�)*�������]��{qL�P=���V��	f��k{뀂ь�[�L���/�m(調�d:��4+�Hސ��O�J&�}B���K�{���
G���6�\�� �����!�?�ó��T�SB�$cүGU*@Tf��~��@�x3⠿�|��4k��${'��t��0�tF8P��X�G�����Q#�)l�g_PJ���{��3��$�1����@�c�p���o-B��M����(+���'�(j���a�� S�DEu���"	]�U=�#ڌ;��|v�L�����?�T���K��mX��R
!u�>�"�g��P9����5���"�M`3������i-����UנۋIq����!Zl$��<a��Q���F��6|�	��}�B���Z���xy�qF�u�Why���@�R֝B:�i�Ҽw�H`�v:t/���E@MƩj��m��s��w����y�_֒����S'�:�� #@�?��ͯM���v��F����l1��
�u]՟W��mj��w�b��ra�ak�:M �A{f����B��5ʡtŪ��s��h/��eJ��)����!��H���1
c��
�|y��tx���&�eǠ������o2�y̱L��Rfͷ�D�!�l�_8�_�^0Ci�:�)�ѧն����qA^@�nw�т�vJI���AF��G��#�\t8�v��]jkO	��d>%�<��2(�QN!A!�X���կCt�M������!���i����a��`���g$`��N��)��K=�O�ky��
fO�-Ro{M_Z�wN���`��'����� X'�%%�8��A�M�������B�	Pބ8
����p޹v��(��nYX�vtA�&w#;~n��h�S��>OCH�DVj��<v�pP�t/��C�'��`��._M�ޣ����H'��s���Pi�׉���.o���N���
���Pi�eFt��trr����Or�%�B������@�LsՍY�vs2?Lezh�eؼ�������DA>��x{�~"�1K�36q]�*G˷��`�p����qe�Y�|�D�yZ	U�:fvޚ��}��S���I��+�2}�!��,�yN�oe.?�/�[oC�y!�������YP0T=��<n���4k������)�|o4�5W@�*�C�6j8�-6Oْ5V0�`z�������T��lpǱ��\�6y���=�o�6��O*���?å�Q���� g�ڤ�m��Q"z� ���w�B��w��>P>r ��E�(�\XUi����k����;�~�Au}F�vN��1�]㔕��V���ހ12�,7|�
\�w���<+��aڹ"~�e.N~�lW�)���։x�	�(x#�_�����-�,��dq4�/���B�6�\�s祩Uی���'ib�W9	��:e���`�<��I�n_��!֪�8�����P��Q�����>՜c
=�mP��KN��f߃���I���;�C:�{@�s���{Lo9��!SQ駎�����L��n%�ev�^ƟUbe�<�Ǟ�sZ)9_�+�-��'��+21z
��օ���4�D�s��tux)/[����ݐS�}\`�ɵ��35�DWW��-�#�L-��7��\˛�$����W2��"��Nc4d)�,�����5������:�����ߒ9����G�E� �v�����ǝ�0�8�&537u_�Jn�Z�>�s8�jF�ud�G��<����]/�
6�f,@�����i+k֣L!/(䂚�%�=��c��Ŏ�u���U,��Pc?(͈���('���^�}��oN�G^�Ü�q��]�]_����Z�x_�z1k����cWQ�J\UV��0A}�J�?М	h�������Ry�p��|~�I9�c��q�#uzOtO�#�Y~}���\錁dk��TF�-�0��/��f�k���$GM�H�'_NpƄ��#��M��OVx��9a�>���lQd�cC�ZH�$�*՝B/I��5;�ѱ�Y'�}��J��Q�|˱P6yP�B���zr�0{�P BEH"[0t�~8��;Oz�F���N��d1f吷EO`]*����U����s9|�XVv�)i��#�}p�9-k�q��N��ݙ�"g�w@g�ʏ��-&)������Q�S>=h����j�$�4}$Ck��`�3�O�
�VM�����>)U]��"0�y�Ӄ-T��B*U�=����B�~+�9Vug�����սC��H<Y�<�%2�/&*'��lKx��C�\"��� %\D��6>Ws��z�7�*G���3����R�LEYZ��#z���|�S�ڋ#E!V_~�Y/���h&���K��Z�xA������߮+�j�y�Ϫ�T~�g1�b��]���;��KԿ)�D�z��(b�4@zw9��n��G�B:T.��E�}X�oB���#S�'M�h� _JCk��q��8_����S�D;Uz�&{Ƨ��F����E�0e����q�~��NU�׸���p U���+��ж�7��y�7NHi;I�I���m_�P�$!����Ѽ�������n'���w�Zd�_�ψ�����6��x��R��O�ּ�	�ԅ`��U4��qFUP������h84�Y[ѽ��F؝��Ş	\��213�r�B���ZAX
L��)�)F�B���[ �Nq�i���z��U{�[ 0��gǽ�l\�h�:A|-X��" �����)=��}R�H���Y'��2�DmL��=F���"��ÄIs�{3?�9�u��!�AB�
�BM~L�tN��=�]��q�H]�kO�H�����L¢U	K>N���<�b���\��B�T>@�ezS���##���zNA
>U�K5zod���L��W�v�@Nj'1��� q@��p�Ѷ�e���9���vp#��ռ�Kl ҔQ=�nO�m����
��"%����c.g�0J��nf)����1��r}���f�c�gd,B^�
u����߁v��ʃ�km�8k�,9�C_�ƂHe��3��	g.<�H0�c�ǉr���?�Ǿ �x�ѯ��$���9�5��Y���7�����7����|/������G����{����<!�y1%dny��F�N\2	O\����U�'�gh����j���+\ xiZ�8>mRs���S�x�&�Q���T��^��*9���7�M��t�?5����[��y(fZ�w�n���xwUr���'c��;�e�/�V�S�(S����Xԫz>�W�C�GEK�}v�0'T��E��0@������Y��_�őM�5�D�#X��Y�i&o�h��F�=�X�N���qG �"4P0�tD�@<C[�wD�=�B��(9���E��q�l..�=
Pd�m	�T��۴Q������z���xi�����0�ڶ�_?�W}Kٍ}Mw�D��y	">ׁ��K�5��֖l��*=�b�Nx�!�]�bd��.�@���y��"�T`X%Joz�����1���V����v%��Έ����� &ty��[��2/�-�@���/5�U��͑�ǵ&�8��n����d�y�`��w]���6#�}�N�!����W���Iz�q��u�?��%�:�Q���K���7�r��'0�7�(v�U�a��2��0�������bn%���b���G�j������>�1/J���gZ_R,��g�@&.��l�-�����-ץf���Ј]>��m��}�ur���s���*��)�fZm ����B���2����-:�TrW�[�Jl�z|�^����i��6~RE`Q���B�ϟF��"�w���0"�*'���ĊP�Y#]���ipjc��(������`vҌ`�F;���<�r�r��yv�F��A���ڭ���̈�v��*�����0�6TS�5��Jѣ4~K�a�8'V7h2��m�Ӟ��˨�Ȯ���}��/��=D+�V����K{���穛s�!�w�$R����I!��=	�yUKR#u@�����=6��z�E����w4�|_$�vkm闘cW31a��{�&�?�֛��Ic:�Il:�~����m��-���
��r�YS�b�����s�q��$`V��>��I��4`�T�NZ#�,r��a�Ŋ��ذ�?����v��H�Chl��HVzv�� Uf1��PJ���ˀ��J��>-�R4s����C�m��P�CRL�j]�
�'��>,V��aF�uء��W���7��<:uꝚk������[�:B*-�qp8�<��`����0٥�wp��/�mvwvx1®����B�W��$܊	�d�I?��(�sG��V���;M+��|Up;��K5	�N��b�bT��d��/Fx��*~���|/,�cQ�Hf�aR�H�h6�t�ƺ�3�t��M�}5����R���Һ�1��?�Z��������,�J|6��m�8�n`�� *�\�D�;������׳!� ���%��z��(�q*��*3�de�gBܡ���Y��_�/R�o��E�B����=u��K��''_���Ӹ^<����	�g�9���#��i���?Փk�{fS�h_���e����rfZ�%�[�5��J�y��Ob~񍋮r���h��u���;��\���*f�|_!퀻��-Nۃkiz�X�RKE,�([fKf��! "��q�8Ɔ��������1|y9�Ƚ�&�4ik{񊷁�l-�e�p�����7a���Tשϖ���3߲l�>��_uFEg��L�@����8�)�V\�x���6�Š��w�p��g��c���1��i�5�Ȑ�x>t'
�1����m�wy�o�y ��8r���qi9ȫt�x�N\���,]�1�y���y�3��޷�P�C[�����I҂���k!���	��'Į�:
vr`D���4+oT_',���E�\�%|���e����%�d8~��*���"��
L>�n$�C
$��|��dŦ\Z����,��t4�17&he1�&n�Z�&�x�@���չΉc�T�rZ�3�걄v�=�~����D/R�7��p �:���C�:,'d��V܇LY��}�� 
M�|­���(�ve4�^[`��%��#K�C�� 9+��5���2�Ŵ?�[G�hIϟP�:M��]ҹ��;zqpQGd�@Î�'K�Fzp�9xe ����[��\���E=���U?״�kL�"�W@�T/�,e��	z�s�@����^�Nr��00Qu �<�6��S�O�Ms �V\Ds(��Ӹ�����O���IY�-��ܰ �3 r�چ�^����N�E���N��Eo �m���#��Z�'���0���'�0�}u�Q�M���hJ��z�'#���=B<��|��cZ���~vמ�.����u#��}.YX�2�b8�BS�^���9)�T�&UCZ\v^�2aӒO� ���δ1"�[�E��*p��J&A���S�=��˳&l����0�9��cxא���ʜ�^Ay5'�I��gɈyD��-� ��x�6fq�?�][?�-t��4OBOiq�R����(��و�p|$O��+'���[CEF��c��˓�vƉ�9�!�9\_���as�|"�&)�&�ʯ�qlCO�!bڻa��1S���&1�����f'��	���R��Y�3��33���v6=~��W�b�;Sא[�56�N+��	����P�'yW�?�%bTnf�0N<����!�Z�Kͧ�]`)y� ����S��q����$y�[�"�d>��f�\l�拆?�H�rP�1%�kFi!��A��2!H�&�Ǝ�n&���9�92� -aY��X�T�Gy�L�������?�C5G���,͑�D�����J��x(g�3��L�<�{ ��i >Xu%�h9�Q�zǢ�i�.�Vi�0u�7��x�*آތt�&<�z>���]c�is��$�`L�/�돻Q،��4̦.�f#�LYd��������V"��Ov��%��b���β��8��P�zQ�^�E���X�g~X������=�­�]���?��[,��LS�1��ϟ�M��q7i���I>�e�=l)��$�,��&�Rw���Ot�Oӊq�N� %��	�֭����8�*����W�N�l���� bv;� %��ڰ�1r���M��K.Sп>!}�dPl���k嘷,���g�g�sh*�X�ʨ-ߛs-� �ۢ��:�p��#gc��� 	S&����]a�������PƸ�'�-9��G���X�yg3t��g�&0��