��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|>�qT��>��*�0P��]�*��W��l].UDY[q����<��;0��ꂂ?��Q~ͩ?E�Ûݾڝ������"2k���[�մ 2�c�Ü��N?܌�7�;�~y��}�Fv�J��)m���v�t��s"4~#��e�w��O��,���o,?�1���>����׎uM�Yx��/l�yБk�!�^k$q�u"4��w�@�jь��qUD��n�gs���2��?���d�㩢Ig�}#�Z�
�̬�\&&�0EP�`a!��J�7���M�`�8,��Г^F����$�����z
�w1PY;�$�>�K'FOa)��զ�[�X��/�?0G-.�rd���w]�_�֗��
�p�dl5Qk9�zN	6�\iz��/��!Q(Hx���w+ņ�V������@21���d�ͪ"jg��n�q�LR0}?��d��}65|�g�$��y�� .<�ט����y��:�_ht�� $�lu�.H�F����Mz=h e^�צ_<����^/�k!U�,��_{אָ���ީ@��~d��Y�UW y�H�k�,�<#k��G͞?�%Շ�5��^�V/���W1����`u�j[��Ao��+�'�*�Q<J��������B����W�'��ƣ;DRҲ_��^�-�#�'�E����R���Z~�od�4��>���]p��E��@]���tݍq�"�?��A�������3��|A��� ���WpYk-]o�V�G���b��dLn�v,�Y:�-� ��ĸX��ي2�Vr?/�S/U%]8U�6~Ir`�7�N�9�iIj����s���aYЅB�����U��E�HΚJ�0�K�,��/��U��qBs�_vw�.}+�>�	��<v�u�ؿ���]Ye���u�T<�;ѧE����w��Wf$�Ij(���d��a�.�Q>Q�,v����Y�>h)���,�Ɖ�_t��	�&�r�K}<�nj�>���� �Zt9;����D�!�n�5s��ww��ˣ#�,�b��@�@y��n`�-�{K�����-�(Yz�vN���-a�q,�R��k{�+����0� �h�m�)�=�zL��1�Z���S� RM��>Xp~��/e�{����TXU��76g��B/%�6�Z*Q
5�-e��<��b�b�^�9Uvh��w�l ,O�B�}%�Ͱv�)�+����%���4��E��ǯL�pw���ɲM����C���?�JЁ�E7���OH���CnA*=��z$a�Z�{Ba��,��?%�h�qf����x@ޕ�IY��{?�Te�+��ߵ��Pg=�x�E/����D|��ڹ������B&A����as�ɘ�62|*�B�%bż�`xU}K+#��GΩI�uI�����X$�U�ἕ�!�g�
G�:_��Δ̄���Eih���`��U�1txM�P��8��cb�S��[�.��JȐ� ����N����x��q}����F��R��ɢ&�\��%,}���j��qZ��p��K�`0��A[e�}���J>����^��������e��HO\�D��uګ�Y����.�����`����prbц���ҩ�����������͋D��p���H���b�����x�D;%�,����^�92�q�uC�g_��<hޯ���)�{�F�]����)����t�}����!��LS�}��ڇ����]%����ހ�U�G�+����
��#��W�:!��4x��_�qVA��-�3$�a0�2���!v��c �Q�W	�%� ���վ��2�u�����jJI"{3�U��i���2j5Fٹjk*?�E�ϊ��>/۝o�9,��`����G7wu�~��q�p���M4������}�'�K*n����à��/���.�ݣ[`�d ��lPE�B�'C��ٰR�$���n�E�nΒ�ח8v��#�V�9T�˚S�J�^6�;,���f|=��%r4�).c��k��a��P&a���/l�'����|�l��c�	
R�-����C��r��w(3��X�� <'i�����T9<ool�h� ���E"8E
hI#��k�%K����]��8�5#t�7)
�����Փ��@R��4o[��|��w	�ʘ��!�j���2Io�35Q�)�<ZΚ f��w
���!<��H
ȤSM���J� ���ߧ�ȭ
`2S��&~���~�a����S�m�u�/m�T��.��8�0�W��?'_��T���өΎ�!m��dds���j�H�� y���\�oݒs�"���ŞV�)|c��{��P{�bB�)�:����q�C�����_��ԓC�u�PL,�h�,�^����?0����k��vH3�?� �q���6�����0�D�vI����R�Sc��M�)#��d���bOX��Y�I��T�!Ή��El��kMlJ��}
*>�	���񅟅��f!q)6�T�ݨ��:�K��A���ܠ/�ة<�-��ե��a���yWh��?��Jm�>�Ý�rB�	ܨTH;��z�+���U�P�6���B�*T��혪!�V����Z�;�҃$OZ-?*Y���3���=(J�����d�-f� 
<b�D2�q�����^�tT�K��tbxr�z=@�Om�*����A�Ju��T<ߛ*!��$������D�~R�̓G[d��PΒ�0wBw)���-��~jH�M���8��g>U�~�JHJ%а����1�+�T<|U����z�����0T�=�͏�IqM����Z��rp�_�8�3Y�"�f<Y2f�PΕ�?U�_�к�}����Dd3�v&
�T���7)��l��ץ��WE'ܜMp��E��� u����τ��J�����ķ���v$9Z�=��O��1�&0����|��x�*�=	n��kf�̾�]zu�c�i��\��p��L>�ye<�_+_�qU"zۂ٨��W��8 �k����k`�2���l����C�!ޜ��.��i�@`�����"�A1��@��D����dI�BW���M/~�%��)�QĹb��%}�����|2ϾV���U-IƎw+Sv� �l�˨i1]y��<�\ѲK��)�  �Z��b�p�)�,�t��k��d@��欟pԛ�ݘ4|(�Ye�^;g�	�vN䳱�� E���"~�-�@�����oy�����j�KI�c�����3�vY���5�}���($��fx�4�He����*.468�H���0��~�>�-r~)��K���%���f�u�-���B�wW��?�p|�q���ȟ<N��0�<�ӗd����*E�� �H�c'7������q���U_��!+�$�VP,��} �fW���T��?��ͬC��H��Zw�0���ܪ�����N-��F ؉�)��=�\�����5U���W��/�H+wDSܕ	�~l�+���^I�ͦ��jkġk��,&jF2a����	4�g�ej���yV���,F�a>$ï���ݏ���J���%$E_�L,.���W(k$ >�f�(��7��:�9�!�	�c&aPqZcB4p*��?��DH��RG6>��o/�?����������Jfu_F�I��Qu�m��g_�kk,�̨xܿ��P�4�1��EIJŏ��H�Lc�: S�%a6M�M��@�5c<�	�����*@�����9J����ר=P��%��
a�Y	�Y�4�X�*k�����ժ_&�E�5�6��O��iRI@U��	�aIE�y}3ʾT�@���0�В�w����#n����?�Kg�u��.^�p�:E���'�L�?�E�Pœ�ۍ��ji����`�,M�6�z�6{=Lj�gy��V