��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��/��Q�w���a5P��B�~�/�'̙���S{���^�qѝz��'�hřD~dVr�F�!5�=��[�\�bYzy��d�(5���*������j M����J����Cw&�u����Dg��>_�,��o��3�9=]�sn��5���A<�-��Y�,���AU�G���̻N�	�Ϩ�g�ϵ�w�Ω�k���R�9HO�o�u�(v�W�T�yVL �q^�Q�0/�����)1�cڵ�E
�W�D�t/�Ș���~x��R�X7�]0|��?ͭ�m׭��e��%\rN���H�i��8A(_�P��0];�ű
�0�"��(bJ��OV�[�0h��ɛ�}<pB���oUqe��]k
�\3��Hb��\bsIĝ(�GV% ��Y)�"���t@����o�5��#
�!&q+���QI���%�!��4�y-G�XIb�*9��O �	�x�eMB����|���ß8��܅H��>nR�>N���3����-	j�c�3W���[&:9���n����V:W{V�2v �su5�����b]��%�Wk�P���_�l[�*h@X��➀K�+0��}H�S�d��PN�|��ݻ���':�qdj�CZm��.):��(̰ǻe��a��*��[`&�m+� ���p�p���5�#_8�Gv��J�S'��mq-��|�Ĳ.��r�m��RA���1�M8���q�� ��ʨ�P�_�I�\��8r-/)Ͽ��6p���h�G����b-�g��,0+��<v���Ž~ J�a���"S��	ֱ��h��2��\4�4����`)���ܿ�Br��_���� ݒ2q�dN8�uZ�����N�>�C����Q�D����C�8 E��ᒍ��-�!l�d 5���XXWb,�78����-NQ_;_?�����/�s�����7)���Ph���H�f�Vw�}����{D��SsBogX�I��a��WU�)�,w��G��D�Rj�� $ʵ����;˸���&����]���$/B��5[a@���������8`"<W6]��5x�V�-�݌�Ei2�&`o�k�k�;�X��u�*X�kz��N�ڐ��@ō)�x)M&h�+L�_P���GO��!@���$�K�q��
�a��sA��խT��O���orP�
<L������P3>[䇈���Îc�Q:���_�� ,2\l�kcw�/IQ�mw�+�V��B�L	��ĎO�q�
�ґ6�iW�V�a�������x�F�P��:^�؎uL)7�\+�t�Q	�+�tC��,C;��8��u �ۼ��L��Q����]>�>|x���a%��2���7u'��Ss�,��cD�����䙕)g�������������yT�D����[���Ĥ�m�OD��e��é�4cٟ�Z7��b�Kݢ�(�1D�f"�Y��VZ�tg=��R��II)����79��.5��*u̖���g��4��N����O�Kux�<����l�kp�v�r�����F7B��;fw�=�?"��f��H��.|�4uJ{:7�O8◇�㑿��lz��|S�� :���{=C��[�!��ڲ�mNܶ�SӅ-`6@��R�m7��8�?�, k�I@K���y%L���}�B���c� �w�I�����_<_���T�E��*�m�J�`/R�x�6yW��;L4Nw�L��/X1�i�o��J��ŎF1�0%��L] �Ql������)ywZE��!TX��VåR�d/�%����^��vp;��Dhǚ�X\�Ɯ�L�����A"��H�E����9�5O��p�q�|@E�v�Z؂�DQ4���'*V�F�"(��d�IB9�����Ǚ	���;AQ��F�h��8w��&�UO5��=�*	Dm��
�նe��h��\4\,�Y����rǸ��mQJA��ڱ#�!̇\$���$�8[e��6=�`���*�w��b��W%׎��UMɖ��*�P��t�|��v�vȜ��^�~iH�2�3��d�4�B�:_�`�3�6����}o���Qw�Р�:���6����@q��qX���h�y�����xV�T� ���Y��Z�p
��<���1�w� �oi��\����qw�g���#a�Fu������}	�����9Y����ړ�,�FA�4��ܿa��K�Y�,%���k�_ORg��g�'Ν�$Z����OS��� �k��s)�T�$[� ��a3��-��D�E�6Ѯ)����.V�R�Y��F�d2�  6��쁓�v�(�=LI�#
3|���SUQk�W�1Bh!�O��:Աs���訰�ӓ�p0Q���9�s;�k/�{��H��'�<�5[�N����nk�Z ��G)�{\�Eġ��nxZ��i����3��)��R�޵��l����Ŗv��wylya{��`C�6L�_f|5h�ff�	E^]�I��u�����iN�w���q༲��O��1�Y)�u(��i]�L�{A��{]�"hѕ��g��]��0�M��u�+�f3�+R�mi��=G1�G,���W^��!+}�	!�qJM�-�]����e��9h�O��Ś=��g��ج!MB6L�т��`�9^M<S���T���?�x� 2vg���hF|"Nk����6}�<Hv�^?�� E�:����7��H�]vۄ���Ċ�Ō�ś0�IxС�,׶`�� X�1�>�>�P��i����/<����[�@$��g�Gv�A�3��e(*�����>q�ED�)E�q,Wւ��rIJ����V�`fK8]
�Z��7
�k�H�yɑ��k&o	qG$��2�.G�W����pt�Xň#2&�u�b�D�:s��+�:4��[߮k��!(�A���6aJ��䚘g�W����"R�z�z9s�ڷi����=Q9��0�$vi��cv	_�|�s����*X��y��F�;��r����y���7���X��h��-9��
e�U��������#�$������z��}�W��,eT���ߓ������M��`��z�KהD2Su��h��^��9�����
ƻfA����3]Z<["l�B��Q�L�R	%�i��"�% �&���83���u��}� WtZH��h�Fq0.��:�h\aI	��+������,p�ɽB�T�=�e{�w�&�~�E���r�.N����b;H���D��Q4W=��d������i3�~��UČ!x��VI*�`�s���>+�ӂ���r��1����` X�5��2܆�W������V�)��%�\����Љ����;>���5V��"
��~�#)���[t�#b�BElo��7�R\�z8u죈,D�T3A"����%ב�;d����a�U>�<;[�[��Y1�K][/�a���MO�r�^������&B���v��sO�p�Вk�˫��1�4�㭚�kyD��J  l2�-���i���OT;�.�� ���Q$�����	q�bt\"�f���\8�&>��7���h�\X�9�J������}c��1;j��.����j�s�U�u�r^-/Y�{<���ݪ:�D���W�X�4=��R!����I�ߑ�_�)���xuR���xJ|TW�~��\X���,�`�$"ij�bP|F�C{��tv����[k T4���P8$�s��������V�s5ʸ���8�Gg�Iԧ�ʤ�&J��e�ù}8�6�U��Xd%͐@z�͖s���n�Y�5�IpX o�y-��n,�W����Ii�O��VbO�>{]�nG�b�L��ר�Kަ؜����i����.�ʩ�@`鹋����$/�l�?�~���ւŷ-�������)9z�#��8�&d�_���䑽�."RL��(��}�EP�熫��h^��u�� �u��vg�Q,u���і4��ᢑǵ�1�������cL~�zwUJ_~�_)�(�T6�Au��޵�L}j�%~'�e�֥� �WE���և%j�5"+9I�K{o��6��-	N[��<-��:����z)�6�K�JPT?��7U���K����=�W���WX��w�ҹ����V�ٺ$5����p�yCn�R�� ع���κ�+��tM��˧���P &�-ș���רa"v`]�O�ې9uUĕ���K��.�]4*7�	ꗗe'�G3E$3�Ӆ٦3�M�G�FI�K;?�_[���98�b/�{�%��}H�������_C�5<��S�A���֔Q���4xU瑨�|5X�@V��\=E2K|S�,^�C�ܲ�m��:9�g�W�P�R�Rp?l����к�rޤ߶��Jy�9E�4+�R�s='�ذM�� U|����'D�w�i���t��Y��J�:��_���nS�on��o]�@D���5=}�+R�^����jF�-�c�������}3���r3���A`<+�kK��H(+�	�WtN����
N8�<<�(��O�2�<�x����Bq:P�|�K�휈��Xp�	�'̄[]��Gl�ON#8�j1�&o�?���x��͓���������`�U�!���!*n@�\mS�9u�����I�CޖZ�AOj�t%\�����p.�A*ܰ9�Ǭ���M1>q	�U*\������i�Zjv�V��Co�^U�0P��ם�l�k������}?c/��d�c�<�����	~��{�t����:0pϧq�q��6��m
*O�C&��H��9���!�<�X�,���Q54�*��&�x
�fԅ��HB�O&�KZ6�)/)���5�K�=�;��1l�ɉ�־����Bl[K�����:�;��5����y�;Z�#F 8��F;���O�&���"F(���B(������C��V*����؅���w%������v<�kT�Ia����q_:Q�YO�J����M��ܟ�j/�X�T4Z���ՙK���0��tb���6���4;91�V�ge�r|�qP",��&����̱�]~�2���'����G|�;oE���j��H �r��
#���V)����/�p�VW�V3 u��up�R�^�Jb��x�
%��b��78�ӇR�^M�<��(L-����aQf�e7�����,?xno��B��^q(�Ж�3�^j�)T�,�
x�3]�e�Ĕ3-�DYK�]��A� ݝ�_/�yihJ��fQD�PNv���NKj�����"b=�SBH0yo2̽%�z@z;�����z):II�5�V��#B�����Z�JDJ���ZUHl#�?���D��Zs�ط�u��}Z��Ш��Tq#"*���DPt4<A��J5�;u�+~�h��۴��a7E���]).C�������~��b��Bv��K_}1�C��f$���.g!�����-h�XD�$���S�T���Lk�1h��fG������(ƀ�n����u \P�E� �sy= /����%�&~�i���x;��6�T�t�>(^�b�cG���	��6#:��^���gK`{��E����RO2�4I��r�f��3�8��N����d���1-#4��=0���F,�{�T��]55%��p�AT�nx^Ǣ1�.��>N����"J�	��4�t�R �>`8^�<O<���`�y��� ���'ϰ(:UM��z���0�CT��l�͟�� �����������Q�$C?�HF����c��.�Eq���^�Ң�~LZ4�Ve�;��H2��h��KH ��4Fť-1�T}W���O�:U���C5�t�ڱ��5��C>O�/!����zt4�t�/�#����Za��M�0!e��$�D�0�������ת�~3����5����DPT-Ǒ�0u���M��-	ӏ�+��Ģ��Y�ӧ�����o�+Ʌ��z�3)X���}�P�BO~�2�t3�jk	A<�J��웳M'#�ɊM/`��AX��f�g���[<��CS�����ú���	-��*�U��z�4�1�G�ee�B���df�ÝEʒ,�O��z���A-���_�G�=������6�[�������#�p3*f�_�l����Ui��75�-*!w�M	�b�{��U���C��)c�Σ�:���k�u\U\�Eހ�쒢� �1�״���&��$d[�`b�G��k&_<^�!嶶A��dƍ0���%�u�l@�����Ҝ!T�=��R�Z�۔�kthʪMgN%'�� ��HN�wu9�z�u�Gt���z��PQ�����rU
0
	D6��>m�v��m��iJbu�:�.F�R���l��_�������&y��W���r�]c�����G�|��Ӷ���h�r�ƨ�G.��d:��q�����iw�hYi�٭ʩ/{o�jg+�z���� B��n�
ڮ�XȂz����&�������%�oH��e�E����Ц�gh�,0�#�m�6���yhO<��pܷe��.���a��$���!�"X���<	*�p?��gܸ	�	���d�"�]+�8�(.pO���#���+@B��j��� "�$dm��Aـm}7�9lB���d�cb�\��g/��e���M��a�������>ܙb��G�"l��{>R�"�j�5��M�n.�I������ Ek�M��B�	3�K)c�./4\��]��\�A9�ޫ�;ϔ�Rf{;W�BJ!�ޢ�ܸ)Y~6��Skp�oW5��zF���P�=vl�o�PW#;�PF^I�i���Ϭ����H���5�\��u`���|��ߴۺ����m,��՞ЖC�ު��j̠LXj��x7M�!�p�o!���k��{�V� �;c˹c��!�Z���<9�5��,����b�'���	��Y^ֲ�vW�O��jM�k�j�Z~�Aa覣USE-��FJ��"��(��R��R���"cE�y�*W�q���`�0��s2<��Tt7�I��q=~ѹ���$[������Hy*e��זY�� L7�ʶ+E�(��p]KTi�lʦ�h2j�i���gp~&�H���v���ҟ�{��I� MO �@���ӫ�E�^K�=Z����Qh��Y�p��
Rl;���ؿ����jf�K�%�LP��͟�w��ǘ�q���3������qQ�� U�$n�o7&h��N}�$�x�1�^���G� �?�y�>y��:�ӎ�I���i�P��Ԕ�ڡ��q��ׁR4!��]w?x�>0��є���Xo	
a��b ��40M.�`\z����LC��6�1i�%MfwY2'w�ѻ�=�ߘn�!�Iv��t��c̅��ĢQ%��~71k教�>���`o'��{i�)�����K|;nMZ=�DLL��F{��ED�ڰ�v��".��ך�A��\	d�� �F�=*T8��P���Ĥ�>T��1 ��D�4G�v����!첻Q�C�����'���������cC�0��*E�4t�i��$E���^pH'>L%-��0�7Fd�ט��-:tI��A@o��{N'���_r\���A��loҋ`�z��������� P�Z�;=���1d���f_Q,�Y�����O;4�A
XG�/%�G�UG���O��6�;�v/�C�8��B34��i����P|�i��%���V�iʾ�*JapS�];U|z"���n�w{Et*kT�Ie2��E���Uui9W>l�`����anv��e_p��@��&C�a |��R�{���p��G���J�*�RWЁ�?��:��6�;RNj��m���CR�y����@�
��8�o���6Բ�c�3�sЉ<Zޑf�4����o5�Ϋ�a��*��]��zڄ��_w���7AD/Y� B���	jؕ��D*��_�%x��Y�ῴWك�Y��؇�h���Ϩ�	BU�C�v�x�ɂgK7�hCm�-?�(Y�c��ED�A��Ēn4�9-ѽz���,���Ol��Q�h��w����>��V�����Ja{��t	���y�5��C�M�;��Z&@3��G/�����"�'��O���UQw�����)R���.�$��T��ǉ����_^|Lo�X�r��Hn�����h���=i���������P ���|J���9�EgтX-�O5_w��Y.JV�Mu�8��U�yt�T`�E�)p>M���G8��a7d�������#��fL�,��s��9ec��������Vp"KhQ�Q�.�9b�lRc��bv�8ˁ�n�{hVݔ7�����LG;E������`p��f�5�,�`��QW�,6H�6�d��ǻ~߸9@�k��R쩪�^'�\��ȁ6ZS��X*�!/!���=_/O~��Qx��G�p�.�&
Q����szc?�yܝ1���WҌ����kA��V�l�g�K����]#26>��}��ָ�u�V���t��s�(�T�_�v���U-\,ݡ������U�Jwo͟���N�MAM��pp��j+�ɳ�Il�D�_�	!d��s%�ۻ���dcHvuh͛z�y*߱���*�+�,�L>[�NLA�J�B�f�T̵��Gؿ���q��|cޔ������6�k+��xR�
�Q!�<���8/��_�
W�O�d�m2.@�Xa���1��p��_W:\�G�Q3�WS*�R�E�G���{��x�~�y�^�p=�M��e���-7s)a����Svs�$�3L��V8�'T���o:�&O�� ����Z�e����ݟ��0��v\8=��{^2"�Ԩ�}|�fk��J-�~	w?[�Oy#�{�\��M��I��6乜 `g��M�P�P��=߲�J��M@�s�_gS���\i���v���V��u,�{�A6J��_�P@��s�]�k����o�u��;>j`XƤ#�Њ�1ne"���"���$�G�YL����]��b�NU|��H�c;�k�7c�;��]�؟���p�s���U�?yl��9�a>��)�+�_5mS8R3����|��O��wI+Z���������6ek���i{�r[��P?�	0R����������J�JbN�N��&?�n���B֑���a$��P�zSr�/�9�)�v-6��V*���������a*�� &L�ha�/��� 1?~����@^�9%(V.W�����L�r�):U>'�	�"�������k���B}��į��[�3IP?2��Ϸ��Y���O�&r���a�R5pڰd���S"�`O,�S��_�)�|� A@��>d��+���a_41����^lz�B�v��a7�OyL����׮[n�?PPXޥd��|�=8�4��+��q�������z}G�S@1&�adm7J�����{�Y�"MZn��sw��!���������MC���i(c��3���CY���{�n��c�U�k�+e����dj���tk��Uڀ~aOD䷃�ٴ�Vb/�t���K�+��
����N�vu���H��~�E�.����0zR	 �9q.u�ͶrF׃�n�z0^��=�#+6l����ә}@I��;�6P���​�$z��Gx�שa��8��Ν�n�u����U�k�X.����
���N�O0Yd�K]��)]7m�J�FuOo �S���΂=�
�v����n�C��`j��"�R������������MX�۲��T�P+(/v��)�/�ml����g�1	Rf�$3g|�ʈ  UM���r�̑�٧yb�Ӱ/ %�B�	�t��^�K��W�^#y%�������BQ�C*��y����Q��FH��t˧s�J��n�a[Z]��PԞ]� �m1fB�Π�г�ߵL:��P�* 0�D6T+��җe=� ���j��p�P��:��J��k������H��[]A�R�N��������}uH"�R2�襐0Зl7������{���dmH:+y��A�^�5��U���ha':G*o��pT�u�E=<�3Ftڹ�)�f1�p;��iZ��p�3��]-BQI^PDg���p\�����g$b��N��{Iv���6$�TkJ�4�8A�&��*0S�.��zw�]�U�L����5/ȫ�U���#vĂ4S-(����1���7��o;�[s��\ܷl��WU��gER�EX�&"��%Y".��w�D���u����֑�٬���W�2iʄ�*��˯���c;p8ځ�eN���;�Z9�(tv�(�-݇��������סHZ�9]�a�J2m9��pܹxg=?4�����r6��T�k �g��v�gzF_(��:�y�IE��b�TWlK ��K�ܮ�K+�p�)�0f�6&`+���S&&1��:����~�9�;uH/��}�6����B�^��)�Sv=�jw� �:��+�yS��rQ4oh�ֶ$D�Y�IC��h�A�u�9U7��"��G�ԳG��l]Wu�e����J��|�Gl��u2E��1�t�:�����H�3�6��@�p��)��í���\����8�!>r�v���x���J�a��ԕT�X��������/P4.�,����J�S�R�ݧ&�}�ᶛr�^� ���O�Hˊ��?5�L�3�cf�N�7g�j	�3��P�Iv��&V�c{I~�O����5��,����G=J�Ԇ��D��X�ȱ�c���S��Y�~�c��c�Тq�~4�g�+����&��j"��e�`³��s��0�������g
]kj���jM�i����B	�>��o!L�c�c�D Ī�vL2�;a֠YTf9hlD��6��"�rlkJuG��t+��ֱv�6��c���#ﴔ��g��L�B��{Q�[ƹ��,"�Fo�|����U(�J���m��d��}�/�5����<,�j��|�m����c��}R[	k�ș�l��v�e�qF�h���|o�7햴�l"D���
�F]916؁[:���S	M����	6d@&��z��*�^�M/-���'B�47���N��]P#14RO�u�
٥1?	�����7�"�������?g���ɥX���(lLi��D���b�����ca�,پ!����j�l����DX���|�,\o�-�`��u	���<�Q �AH��ϩ�[�dC�g%� c5n������<���\C~:#ӡ�"P8`� s���@<��.���T���^O1W�?�SsIp������Vr5���V̟���L�&yn� N{Ѧ���a�ks��3��?��N�Y�.9��rv�E��j�.vIN-M�S+�)}�4L�9Ȇj:���.i0;���w��J٣��}-{�׊&�ɇ��)b�ӡ$}Wӥ�o貑=bm���x9�5����������8���O��@\+�!�.�AC|�JJ� )9w���nj�?��U|��oX�M9cE(jNdjDF'�{��!�����d�&��l7��H�]H�|sa�Khe>h�L �r�t$��<��ڒ@��rq�-3Q�����)l� g�f Gm\�&��ψ���<�j���������xf.��K��M�C�i:�V�l�*��'�����j�P}4�]�.�Gf��;q�9h}�!�6��P�<Fvh�+�ԁ7u~��>�g޵ϣ@�1D�����fq�!ذ���Q�wY.��Jɭ-��|��%Š�+��K���ܢ�]�~�����:�[��So�d���Ņ&%=yѨ|��������f,���2��4��X���cQ���Ŋ�ҝiU����׋5�c���B�n��P��z�[�ˠ�dP��-C\�W�ӚH��ѵ��Oۅ�%X�6�����"ue)�p�A���ǋ3)�u��LH�T5w�`k�	:�n_�^�
�-���V����m�����@�TH\l5Fm[�[�>��EL,�������v*Ogg��+L��FĄ}��=��m�#m���`��S�x�S�M��/H:*�H.\������
V�P�jO���̘��]��l����������=���)�g�fz��%��eݑ\$��k/Y��or��D��-�_�}ot�Ε]? ��x�?���0�N?33a��B�-���5{(��ݦ�g:B���,�k9�Z�s�Z�>%{�ȷ�3��R��ZF����12F������]��ᤵ�ǋ�����H��&���y�DK�ɼ�Z?k��hX��Z��=���ϭ��`��C��ЁW���)�-�/�ݫ(M m�X����y�����4�J�#"5qɚ�|�!������Һ�^�>�U��6����n"c��d��A��p�]�6�ߛ�N�3�{���(;~���6')Χ=4܀؀1�\_K�f-�'p��U�4��B�k���i��3V¿�H���я�Id=Vi
d�?��ES}J^ޣb�6�Q�!v67z��6�+�nf��ke���u4w�"�o �Y	��Y#���<�b���q�3�����+u���R�����)q�;F�����R���9�\ ��E!*�l%������Ic�=�d�nf�_Ù���n�m�=}*�"_]��t|9ɇ��f'�-�ǁ�j�lY���������xѫ��	�gwm�9En񫎛.�!�eUrW�C(���S絭	��IB�h��)�f_90sz���q�5&B<��ǏI)�+oE{��&��oB�Lh\���� ��� �R���׭`"�nY�iN��/ц��k	��.�9���I�ae��?�V5�zWw�5�t�l|�v�)�f�����O�/�
������&<.h(��wF�<�c������.����T�e�,Q��??�'䕰>�[����%�E�(����F�S�H�Y�9z�]�#���IiP~� ���WY4sa� ��������3!jS���Dx�w�Ă�1~N	{\K�4w��-q�.P��\G5�O+�QHq�D
XO�� _�l>�������.������5c�b4h�pE��Ƥ,^��ߝ��&����'�)ӝ��CО��m�O_.�B� ���g�2%��>ؑ�6�\���W��c�eGx�{����xNv�U���1&���J�^E���L�O؛(?V7��S�/
}�=��r1f��J��ۇ�W�D�E�L`9〺��@6>�d�����h��g��X��ܺd��]�d�L!�5��
�pH"`דq+V��s$��x1O����]h����Yw�9.X<?�To/����Z{x� OD��{M@�i�{�+�(7����X�ќd��6����ׅMQ.J�N"H�1k��x�ԗeZ"h5�c��N�4�DX�Լ��
��?-]G �b��oZj�>��t9�\�� �x^0V�5����A;�e���5�/Z�����B%W,.�c�$�#7$m�O�岊߽�)bX��^��\yH dCɱ�+bV�#�`_l$
'E��e�Kx�:� ��/>���^˨K�!^ �b��=Q~�Z���Ƙ�f�<��y��[�<���S"4%���א��j�/W.����R��И�;�3RaA�)�J�u�d��҇�C
dM^dHaުLP��g���a��=�_3�Z�L���W����K~�&g��i�%�ٙ2�t'h����-����NS�����[�
�x%��_�@�,��ʭ��|0:��:����Vq�+v�'���f�?�~=�V+�ո�
��Z�w������˅�v范�_9s��FY�a��I?佬��!;h�Q��0�Y�D���e- ������.���3�~9JG��]��E�[���U�/�R=~���u���1^JV��Fs�
�8�]��̻���Ha�,��ӝ�]mњ�ʶq�I���Z3�P{G�^��&�N�⼝h\;.Ȧ�I�D�:s  �*�"}�<N� "R-a�հ!�E��nG�H��w�R?�]IlV��=��$n���� ����|Uo�1�$�����k���b�ڸG����o��3�[k)��/�	��KR�Z������ݞ$l��K$b�7��c6����^]25/�;�sޑ��֒V���==Q߶>�<`�vu�8<�(�������x'!�O��M���&���hlP�ZC���H�C�.���7&�9t�;��VK��𾁾�
��3�J���h���Ҵ�8��+��<��,+1;
�KX��3�b�?��QE��O龎;@h�Aϋ�ٴA�|d]4�PB<Zyn2�;𙱹��D���[��!C�����4�n�PJx�Ƃ���a�j?,�A(¤Jj�	_Րʒ�P7�Ku����S���݈eՑmh%	��5��D2�ҧ�Bvߏz?>b��~�vߤ�7{wiq�-/��P���Bb�,���+�p��O�����[�e�C=�e�l���=��	r�_뾗K�5����%kL�`����(�HR=��ɝFہ��"Ϩm�=ZnE	�]��d��]?;��'�/O����%��&�cU�����w3�l�e�t�:巰*�}�Z���K[��B���v��? �B�;�^�LO�v��T\�D�:�zAдu����W�-y2�r�.�LnWȭYϥ�J2k��+���&�> �3��m�	����,z!�AY��VҾ�	e2!Kt�L��̱�sk�^f�Z>F,.35�E�C�w��ܹѭ�8%���$�7�s	�x�KŠ�
�9t�����;�>��tj�o�&��N|�ڽ}��s�  �
��X[%��Uc���DyD���[7��<���9��	����t�|�2B�AFd$΋	t���g� ��L�]%ɬ�wƅt$���
���H�t�/��}jP7)ÙB��ч�G���Q���߀��@W��V}H��g��BL3��X�4E
B�B����$R|(�T�{u���F��3=o%6~i���� f����/�j�&�P��K���Ӌ=I�?����r����������|�����05�te�݋s ���RSk{6�&M�	����YS o&TE�QG�]��~���d���I�D߳����o6h�a�G�nF�R�C˩ �l� �sJ㺼������W鬁<Y৥���B����ē��5w�:i��IhNy�J�=dfT�>ׄ���.����ո}Fd:l���|r�̶f{Ρ�S��=�����b���_�pC8�(o4Z��p|T�1ʏ�5��$��k�l� ��+l_��8�r%�$)����w򖜉E�����c���U�F�y��W�����P�dR�O5p�܇���`�K� �y�4�|���A�~��?�ݫ���s�f	O�]aE�CB�'P�-{��$X=K��\
�a�d.;*�r���\��V7�"���>�?1�10��s%�r��O����{��i�y�@��k!_7,)::�����3#�8�`l�^@�e�?s���ģ�M��n��g1L?R����Y�@�s�08{iU�n�,��*|��4�7�.�S{�1����1�Ƚ�[T����D�a`�j�( f�s
�jW���@���y��2f�է
ew��e������޶��˿ㆃ�fQ�R���p��� l'd�ۼ�K�7�L��3��`�Fۅ��#g�g�$N���9�Pm\jH���.���fa����|����~DI��ՀUk����ӛd��>��4.���}��z1�ב��4o����Ƣ4��J(g9B�
=A���6�uCӠ����/�%�1���ǥ� �hxkq��h�[��so!��qvmm�I����B�G��2��Ϧ��Ə�>;?>:��6]�}{ްv��7�3����>Daͼ.�\�Jġ5���h)��q��~4�R�p.�,}v�M�F͂[@�r�~C���h�6���c��Eؕ�.E!�cԥ`,��䁌#�qv�����}��3�y�?���g�RБ��ې�\S>����JR~,-�U��n�F_|�����<�=��R��LC�eF%=%x}����"!�Y���}	�*CA�D5��o�LƷI���b�bd����3:�hy깋a��H�}T�A{Պ�wP2� A��d	��ߎ���ɜk<^�M;�he��^�S}�,[���{�/K	��\㷥k�^��c�/�/n��!fM؇7y�jC�j�=�Xŉat׳B6w��6�*�æS��Q+�ܖ(�����|;��е����~��^h��<Z_C�1�舠��*�̰�<;	�%�����Gr���Yi�Z2	�H0�ʾ}��ҏz,�.uF��8�1{d�|���؄�Ӗ�	��|Вo�Ñȃ:Ȍh���}��ݵ�}�*J�,���r��z�
�S����}�^k"�@�UO�a���-!l	зpv�0�w�u�uQD�b�?�L��W:��qK@��&^������,2������o�R4��V1���n�-����Җb#�y ��H�S�z���bD�g�xW`jKi�"R��u<`������N�����YD��t�&T&�*]\R����vᵂt��{kU��&!����k�����9YA%$�6�Vn���,v�Ґ��/�$L$���m���5�n���	\;���N*�:ج��b-���?�P�y��)��(�����8M
��r<qʍ1���Β&�I}?��=K���9�}:�gʮ�� �n)�I�>i4红�'򆵅��nc�t��T������Hs㋰��H��+B�����F+/5�������)��Au�5�+bH��NV���*��!b��`	8��W�q8�)(Jn��̌���6�R�s�Ss88D����+s�Nm�@n��U��m���<Y1ڹ��
��O�R����7,�Ę�?��@���J$)>�.����u4������k՗V��'����z�d��C���E��q�E+T�XJ5��^/w�jq?���e+��㿸��l�F��!7�F����4ڊ����u�йY)i��L���(tH��?�L����Q�dW��4Vs)��٠Uc�m<�t�q�CX;�5� �*��yEU��O�<�H�Ш�|'�(b��=(���:ԟ�5�o�e���ru�?z����H����W�I6X�X	\��ī'l"�R�8֒mI����Z@oQ1�A�ή�
=��O ��^��ԉDrQ��⯘���9���<+�^�?��@R_=3���q]��M���K�o1�ъ]]��EY���h�I��8�Jm��Ǒ�ض&�a:��'׶��b�ĉ�A��\pS
�B$\1�%��8�p���7Y�*��b# /-c]e=f�n�k#{.��%��ɐϫ�@1����*V��)����֓B[�U��6t3Z��^*C������z�l"˂�����}f���.�X��D�Ȑ�g/��N��\<35
��+\p�X
���&��@����>��Z�9�|]Qj\�=j�d�Y°.���j����ab0�n7��  |�ϐ�֢���y�d�����fl�6�$���ʚ��diR���
R�ӛ��ߣv��c��kD4a$_��/�~��yX*f��3���ŷ6����-�xbF6��j��\�&�?�еu��t	�B	X��Fov����H�C�s��i�����K�ҹD��fB�Y'���PsU&*.%�2�jM�!~���΂ad��&���/d.����<�v���(�M|�$B}(n�/]�Ǉm�Y��绚����^���oY�T`_8���ȡn�d���7��y0kj�8����m~�ɣ5�BH���e�زR^�Ihǂ���⚗�ǜ�~�|�r��N{u���AI_}޳��Ve��a��M�ןO�SŞ$`����$g'}d���x۟[;��m��b��Y0�Hg�>��<�ѐ~��-Mk�8~PZ���"�&ց�����5{��Keà?��+�02�� q�2��\N{/3��I����k2X����T,=/�ѻ$՝PN�Y�����OR'�Q!�ƒ�q\�N&�氰=?�sTΧs���GOb����J�<�_<
L�0���YhjЙu~�~�:A8~^H�1�h�7>��1�NdLe�#i�r֫��欰����<���b{ͮ!*i?�#�X;�eH�^`0\��ѩe;ר53�_�� Z����&@��c����\�F�r\d>g�F��~E+}�&
 j��v��,�U��i0�����Q�̓L)ےd�]����X����Ů�n��[��$�@�v��ܛ���	]ant��3�H���QC"k*�lk�N��z�$ü%%�؛&�-� \�ØM�vfH��z����b>�ڟ��p��������*�ֳV*�a��/��ڷ�o��U�_@`�!�������}$e��ݶX�7kl�]���$n��$��8�ֱ�t����c��^g��S �֬S�^J�MS�ߢ�d��K��|#;������9�Ep"&���~�3�bg��!�j�k��m�'���,�}��[�cU�Ȯ�ú�7���6���򘶔kv��/��s���8���l�*��s���L�ݭ��ـ�~:�:Kv-��ѓy�ŭ$ݫ��ݣ=��5���my��/
����w�7� Z0��C�k�J��bI ������o+�q�ŷiG�DĬ]����hܔ�5��z�s޻�=�Y�Ώ�s����(�{����yƐ2�M�urce�2xl_T;��?�{G`���/&�9�b``7��Y:ϓ��[X���x�怰7�$£xa0 ���ƵI�m+�I����E���%CPI��nt���{8a���4%EADg�w�\}YfD���G,^n����@��: �u$�d���÷�����u8��2)[�j^�ƌpkU)M�+���4.���e f� �ͫ(�P�q��ӊ�36�k�)ᆅ���>�/�����r'7�oXN���B?�s�l�����o�@�R�� ��	�n�FY�tLk��V�D��5��k gs�*m����*��"���w��m�� ��������-�$N�:��ϊ0�\�諠W.��Y�oo�Gf���+�_��SI ��#H�����Ĕ1���']@J�e^j+G~A���)�B�4\-��k�Ėe���y�ɤ���v�dP�$���4|�I4�K�.��}[o���?�tﰉ�!B�~�r�lTTO��W��&v ?�:#�����+�AC
"`�yO/�@n��r�x恵��_�aq��Į/��O!��L��ʷ�����4&�h�g�;%M����4KgȮ�	��o�!���{�$�O���zSibލL-�Iz�=�����3'��d{=��q\V�����*z�mG�qx��n��Lw��5[��;����nh��u~��5K���INq�8H���/��zf�墣sy&2��h����2���܇ �)lZc�t~�Z��-�D$L)�/"�u*v�x76��z�oz�7��W�S���}�v���^'��_0�^���u�Q��"����u��cG��G>�����Z�bt6���eG8�oh��W;~w����m�c|N5"����L8}�g?�vdޢ��`��H۵���ꛠM<J��)C�C)�,�e2��w�1b�	-=��GP	x�qW<{��qI��z��+b6�/
�
��Y�	�� Ua�3&��]����0�?�ۨ9�[��d6�dh[�4`�L��w��9��>�.���w�D��r@�~�uH�=��ÆR�ͣp��9�y�a�1O4��96�7��|F���\��5��&'[$�x�?\V�����2(J�d���G�O��7��)�YY��[���g���9=6C�ײGeh̀�,�0o�3joE^�O�6M����WS D�\�����W�B���-��qh5�����@�J��u��R���Ԁd.T�G%�mYfa[%��a'o�����ޚ��b���6}5m�.�B��Q⮌��N�	ɔ␬��EE���`ܘ��Ƈ�	�RQ2���.�g�S�}��Ųv���ަc�c�r�	-�4<�v��1�^�S�^�)���%)�b*��oub���"G����T%�P�'��m/�яq�����#���;�Q;Hn�����^O�(`�`��:�T2�����~�I��k��L��O��W�2lE������5�mG�$}�t	?����q���Ӹz��~f�F�Y����E�*6�tA��j��wcs@Az0�<H9|�[�3��@��W�'�g̋��8)��/#fWǛ�S�M�`��^�1()�,�+7���m�ĭ�%�dX]�`�7.n8�?�0�Ad��s�G�F����^[P[]�<�7�(_�&�'�
��X��A���2=ۺ2���W�mxY<��3�H
��D1��ʠz�.6��1�&�Y�K
E�x�'��J���;��3�*19��	5�?�-@���������I�U,i�SL�eR�c��2.g�6%����Y�DB-�om�8�e%3�"�sξd�����!N��VΙ2��K��������g�n���5|�âƒ3��O���mH}�9�˄�Ѣum	$�|f��3*%H�>��X�5�ض5mĂo�4��r䪍�`��a1��LN�����f�y���m1��-Զ�k����{Ǽ�v�ؔ�_�^��'�p{�NN҆�>>oWH<�C@��Rs��d�� ��g����n��=��A0�T��?C.Hfb��z��9�����30��� ��I����#0s�3t�I�#^�Y�-ˬg[*��Ya�[5Wf�ª�j��H]ur�u�Why���!����oK��̨.�+�M�L%����j��_��i���/������4�X�Z����ua��c�'�_w����Tn�p��x�!�V�&ˍ͗���|1�4�\I���7T���%���(O6�7=u�.�����~�C�_0�My�6@#�[xy���/&go�/;�b9$G'zAH��ʬ�z�r��t�(K?�HY��/�� ��1^ʍ+wc�L,�_�Ԋs]9<�HS�r(�+�U,�4jXƾ�mFMA��7�0�nP]X�ҎT��'d���gO��t�ԥU���^=%*v��8��F����N�`AH�y�P��*�[[�&����R-�d����t?,U޽(�"F�s���:F�.��3��F��
���L����L)��������=�������XZv���i������g�~����m|O�0e�ʦ�����N-E�M/`	���Tu�&$%:�-hB�R��ۿ�	����M��=�-���kT]\a��������D�4���2��N�����@��	�&�T�_:��U��
|��M�>��rTr�Sq41}�L�.��*+o�P��* �]G.-��q���4�~�h%9�z)�s�L<f2������b�t��4��C,Z�[�v)��`�a3O�L�-��
���^�5�Ԑ�VhF�W7�adBD`L#zM��~d�8�K���v�k0��?��u�N�x,a�3�$�^�y�Zn�7�Jƕ/zS�r0t��-y R�x��z8�C�]`��,��@m_k��ǔ@��5 zc�q����7����i�C_�8p��=X�~�W�bD�s���Y��	�����S��>����x�9ؒ:�H
#�(��ve��:�*�W	��ѨP���r/&ge��$8�h߱�t��跚7�bݿ۟l-�S�K�	'0�ɝ���<7H0,6,i.��wY<n0�^^/�Z�z�>ܮ�N5Zt�s���ꌦ�P�Hu�M���3�Ԃ��W^}�㙜�b���������򫬤.�y�8sжj�O��x{	��$����.:���l0�������j҃֠0 Mp��M��/�<���*l��#�����|SV�MQ�hhQ�k�ة_�[�\�+���J��Ğ�w�)%�̺���k�.@�$8�J����W�� ���n�����U�&0uCs�Qm����L�;�FЦ ��5+�O����|G��c!+�?-�P��_��uB.�����6 
,�c��5#�Jr̘)O�����os�]k}|��}��%��4���3�|D��\3�>�rN,�2o�#ݹ�G�� �G������o1�˵��6ԏ�c�}tU�Z�$����$���-��W"b�L�yY��{8%�h^��'m-��çy!q��	ɝ\B���֨���z�MFj�2����	����'{0��!�(����]}�K@��P�G�o3F�ry5�������.��u[]C�J|��c	�t_
�YP��C��Kh�z�� �)]�8�%��Yy�f�P@������F}��z�lYq�NTr�}����e�Ɔ�MvR�t!��$Y�#}6�h|8���e��X���=��{ߢ�x\(q�+y<'�S��3Փ�z+YtB�E�oIq�4q�\hs����]�H�!���Q%A{5�IbG�AyN����Y�,��8�	�C���i���F���2}�Qf�/Uf��$[�TVZY�=���`�>`�n�˼����˃�h�z�����u�[is���"9��.UXpyL2c9�ܳG��r!� ⷐF�.7I9��P�i����~���y+�K
I v�(։�{'�<�*k��p��VEq�%=Y���D�;��$��&�AX>._�r�4��(��2dʲB��b�+��}^!c��2�D�_�����݌"]�wU4�u5�N�u�����s9�	*Fr�5I5��b�w޺�t/�/Fm��^g>W���(����yO�Sm��
��q��¢+zQ��t�xd5�M�Z�6kO��E w�E��%B,�d�R�:���@B��pO�ҹ�;YLj"�� ��������-Z#��J�����"�i'P	��m��姙�����r�j]���5�mة�t�2�z���@^"�$B �'
F(s�	�H�>�D�����`���ܵė��'�KQ�7�<
��X�҉��	F����"7�ɐ۸�lc��a�?� ,#�5���%�p�3��,����gI�KvE�]W�&B5�z�;z���o'��C �.T�.�82�gȁ>VGzz�Ɲ�"듰��O�V��K�k���(d�&)���2Rز��L�WO�E{;�PA҄~�H^P;,:����_W�&�2ȧ��jT�	�h����20D��q�rg��ipC�
�|��Փ�3n��|:����h;�Z\��H��gd���'��KZc�7"���h����GP̻#AK �`]�-�Vbj��V?Px[z�`G�����yV��]D�#'��nP����](�AJ�77�oW4 �Il{��Q�
9ATg�|~=���P��8���S�j<����q^��e��9%��/�d-{�JN�e;$k��k������G`��>>�tw�NHʵM����y�3�c70�aKy�Мh��bk�w��s�h���R���scC6���}.#|�;�b�zv�	,��݄�܆2���(�w��{y�5+��s%C�"d ���IU�谄�6�k�ڋ����(d]H92�d�Dv���j͎���`��K=��d�M�G;-\<��)��
�Ftb$.`�,�����}���f�h�8H���cD�e���9�O]V5{�ac��g}�G~���G�R�'���j��s�3�V��0p�e���P�MnZL6�l�5
��5�x�zY���s�[���^wP-A�P������Q{"� TL���{��jGɲ�u�u�l.�,���_�����ۊk�j���ȋ�"�K��zN={E�,�r�x�F9�� +wi(��T�{��!OGB�����Shw�[�zu]�5ҥ�0��K^M��\���ǅ�$���G�Mvt�̆+YFZ,2v���K7�&/Ϥ&�VC��>�Τ8�������9�?m���Z�7�����Űp	�E��3�pt\o/]'�	ܻ�<$�f��0�KŚ^��*^�>�M6c4���XPA��O���X�cB�52�E�s��gX6ŝ5Z2�mM"Bu�,�_���.o�
x2x!C��l�4�}ؑ�.��^l8Qr��B~O�
DD2��Pt�/��{��õ�sY�V7򚊎�7I �/��'Yz8,����H��p`|bn���T�� >��g����^f��?h`'�����\�&�Z��j�;O� 6�����M����{~���c��#�S-��l
�j;�̧(�W��Y��Q�N��y�_lWؿ(�s�i���Yt��p��dr��܏<qlF#2�� މ/�m+vxD��?���]������K\t:s�O�E�;n��=f�=K�$_�ЫwQ� �#���yi�x�ⷬD���]'mr�4wWS�֋�sQc��0VO��rTJh!�^�/O���[�� Ċh��DD��k�r�I��Y����^�=5��9m4�xxһ'���k�8){m�#H�����jX9�1��tF( �����*b���C�L�s��Y��Z���1�\�er" �u���t�� Kؠ��FAT�F�^>����-��VP>}��;���> ��IV$�ԐxY5�z�V�m�'���ܫ����v�ܗ"--z���MD}�ŋ"֍�c	���=�š�+e>���\l^���Vii��1D(�Sv��K����7eJ"��ǦyëJBFٝhG��r��κtޝ�r�;%��L���%.��	��楐�`hzsF����2*��-���J�H�����Xa����~�����|�t�d4��1П��c":��>;�O�)tK��	l����I���S��r���S��B2M�4­�*H�^�ߡ��Λ��2�p��L���1@G�1��Y�8Eeu�ü�"�0�8%]�0dfx��1%B��A�kV>K[��T��X#�P�	B��m/)6'4�{�=p-󗷲��h��L�Z��T%��nO�y���(h�-�LX�VS�ÿk������ �^�tOҥ_@7�Rbd���̿��GK�s͹��J���9^�-�}�:i��~���}��1�g�*Nvn�Kh�4��W��������6�*�ɴq�3t@X�e�4V���#��$YϬ��;�\ݵ��F���'PV�t�(ِ���V/d��)}��7� Wjm�6n���[����(�{h=�����x�9�G��^�0����p*B>��㵬yv��
*jv����G�u*�V�� �3������Z�|!O�W���偃
���פ���Rx_0ef'������~��YT����E*4/�[�$�><�W܈(Q����"�&(�z,du?�f�$�ڣ�I�kNp����m�*����?��[��������w�tZM0i��/���ٱ�$o$C ��>�꺰:��#�� ��O��UWpnd_�i��Xq�8W�� �DV�NW�hď�t:XK'j9\2B���cB�I�6��4����F.���e�L����}6C|7��)�h
�n�|߷LEo���/�9� �������%��-L��|٘r���#@8H\5/�$N����M�J�˩:к�)���5�'
�-�l�:��2�|�S��.�{ ��,�r[�B��Y����m�)�K�S�Ƨ�*
l�+6�05�HZ�6}����ȼ*B�zс
��~8Ⱥ
�"1������) �aw1�[<0��=$\��.�H �~8��y��y��R��(%�����jw0��k�t�oQ�s��v����3=݉9�d��e��Nc>+�c�#�Xv��E<=��� �K1�_�qdI,j쀃�t�Ii|\ifB��-��I�S<p����� �ۡh �>!�0���8��΃4x=h�-��n&�|(L�w�U��y��	F%�e|&�#��n�Y�_H܁z�y��ü������	��Hw7����8b_�l�CʆT�M��.X7�	w �"a�K5u��"����1B��A�{�*��@�>8N��%��¤�f�bh�[��;X)�~sMy����R��>�(G�(�m*�C}#/�3	יd?|�-�\O�ͪ���]��m���ڔG�?��l��E�� ���s�~J<d�z�.�%H���1N̓4:>&ѓ��h$s�p�9��lS��'ף�����9H����Th1�9Q���y���X[�X������*�Ğ��Ҹ?�G�Y�J3�A��L�M�M���	]9�9D�J�E`�v�~��M/�4��vˋy�BZ��[��I@	�K�
(00���SG�;�2���	�C"���ڮ���i����!"*3L`]��s��k���t�vvm)���H��S	�!�d�y�G�`׭L_/�����t����Z>�pk��a9��ؑ���*�!ɬ[�/$���f��8�b*��9<��I���$ u��`.ՑQ�SW��F.�ٷDk%��R?� R"HSEX��᪟5$dG�6���b���v: �F�M�2��h�K�:��k;I��<�fU�H��C� �ҞY�_NUN����n;R��}�˴��$[��[�0T�v�\G���<�e���קL�+��Qc$ FM�r��d�O;iO�d!��7zV�� 5������sh;�Pl�<us�U��!C��J��d���I�U;t�ώ��΅e!�'a����~?��9�jH#�Ɉ�9�]�l�Le������c\�iI����!����P��� ��w�ȯ�s��>Z��Ɉ�6	�|� oJw�}9�vO�R��Ƌ�f�1�o��<"����{Up�x��Vq�W�A��#߃����J�fH��]H�:V���̣Tat@'�(�&j�usgP��Z]N���k+��ב�6n�{�,H#L�h�ݻd���3�J2��#Jha�49q~Oq�*�&MO��k���E.5>G}�A_���!��g.�qg�,Gu*���2� �0��C��K�i�/rE��(�a�Qno_�׵>�����r�e����({�e�E]e?A�M���`���e��B��Zi/��J?fǆ�%YnR�PM}->�$W$C[?��,
J�'8�,�N���Y�� ����;}��ۭ��Tn�Ԝ9%q�w�(��~'Ԩy-5����l�oV���J�-���73�?S�JRؾ��w�������m%�(����F)��1!����$��Y����՗ş3���d�:]��Xx5�"sI�ӫR��xʕ�����D>����󼫷�4y��
>t�|�ߢ?� a�(���n-�@8��bc�.��2��+���w�5�J��+@�G~�6�]���L4��S�W`�����h`�"�@"WHҶ�q{�Zu ��(k��,�iC6_#��s��\�$&3��4Rg0� :�P�8uJ��*-�a��׿�ז��yD�R�H׊b~��r�e��;O�>�Z��6�_����`��j�#BI�-3:�k�ؙ7�c�4|����.W���/�|���Y�*9[�J�k�ڇy�u��w�_Yϕ�b�� �Z���O�ޓ&{,<�?��_	P����A�dz�b8O�P��%H�0a�}!s����h^YP���,��HtIUd'�ͅ����3OY������F ��y&U���i��c��W\L�Y�,����Z6����#�k��!�Dc����Ñ���o� �[���,@W��4m��	r+�v�lJVcSJ�����6(�]Z��N;� ��s��q���6������F���/�95^a�|)B���Jq!�J΀_\�]A��w��Gk��m�Z��'��1�f^;d{���Γ�|��Os;s@P��T�}.4�7��V�����c���Y�0
��,�3�k�Dh��d�;\f�ſ7�8�/���aҲ?41d����F['`�9��z�Bɾ�%{���L�G>��t^L�׎Hv���U�჈�Tn@�ǪQSp�P���V-�W�DF6Ҷ˂/�ZF�|����.�F���Vt���e�(�%, =��N��s�}��LP*�(��,��c�4e�m0�n|�s�R��fX�����Fdb��@��1m�N���%˛��T9��Ǝ����|���0�T�
S��g��w���+2�����̘4Yzڲ3[���W��C[Y�o�7��C�%|���H��K�N<�ʅ$���yF%șF��3Ӎ:�D&�j�ώ�R`�˨�~L%�0A&�^Q�Cks����#�b��p
�����gfKc�}�[���mMzW�3���U����E�3�J��`�!c������X|�mJ��u�	�峚�"�F����܇ ����Y,�m~|P,,NI<	?[�S1k��q�R\��3�1�5j��I�3�w�H���-���V�v�٭/Z<�L.��ƟQ�l5�������q�Dn��譟K��S@��QQ��{��y�Ձ��ԯ��)|}�(ɞN-������䶆�<Q����
@�6)ʭE����������=�ھ�m���Y�?w\((0H|��Ȑuzv����)��c�![�t:�j���J+����?n��<2�+�@�詾Yz������K�i	~]b
�7�"��ex)z��kG�5��"�A=�r�ŵ��m\?�˅�b�8�뱮��-�gD-P������7Jb�����=��!%���L�������	�H���Xh�zLI���<�v�[T�w�9�]˜R��$�%ޣ���1�C�BC<X8�@���/�ҵ랴��]�._�	0�?ܯi�qڙ%|##��.g9�<K�{/�zFC��{�h
��q�V�5���F|�����.l�xe(	��K
�8l �6�ii���29�ܷ��kl��ĉ@�������:n�������br���	���.�Qs2P%�6z[۱�͊���இ�B�r�'��E��<���=N���	8�	����&�Fu�or0;Iݙ$:n�u�O�_%b���~�r��#�٧Ι�\��Ow���o���MÏ����v
H�Ϗx�FY���R�շ|�����+�q�%]�Z�Dp�?hF�m����r�������D�l��QB�h�P�r%(vP~���	#Fܳ��#���4�^G�E6�i�1����1�����b�H],k'�a����@L�0�o�AvE��]簎�Ng�Y��)f�J��raߍ!D��tZM�3����`��M�ۜ����C
/�<8k=w�k����l�6��V��n�cp�P�`�F��)�[擿y;���;��#��c�[u���[�a�+����D�}����4ka��#��0ę�(�0�9� y$ᵂ�G� ɢ�%��k�@\g��qJ�K�����)�)i�^h�g��d>"�,�t�GvT�v;��|k����f��`u~�)	��]Kw���M{�D��NE�@8p��jL�r4�Dv�u��1�ąs9�4��EԚ������*KFP�mKy{�{�Q,+�>e �r��_����s�Pŭ��,���&>� �Ĺ�����h��0��1�Eˢ���J�#J���>d��1.�x`G�u�Jʨ
��f��_g�����,��{|�����a*ֱu�^�Ldi�N�`�w��9������e�����r�=r䌅��y��e.
�I��Żl�汀���q+xHD�9ة�$�?oä�{3��0��j�.'�R�}Н�yè�0MV�JX��O� �[I,0�<�[�,�2K����b�]{�h��;��h�/g����`�8ݔ�K8=�'^�r8kD1��Ņ�o�NE�q|�p�K3���YD����~e��(/�l�j@C��"#4���TM[�ܾ��x����*u\�9�&7�|�;ѰB�2};ː�>5�T���;�h0U;i'�Մ��y
�$�XG4�a��F�����'Ow�k)�a�n�<0��=�,~g@�O/Fs0�j��]���ܫ,&T�ލ�0هH�C�R����T��k$���E��Hج0��:���ތmڬ�q�n�@]��e8]���&�tkDX��7d�@���kMD[Q,���\�xa.D��#-��0����dҽ�V�YH��r}�<^+�~�B���3���:m��@�%bE�T��7�_;lOd+ I�A+�2��]R/ԯr\�=�y��k�xxB��`�E%�	�w��
�a���j@�]y�,��.T#8O&�O���� ��F�||Y"�`����8�g�k};�����)?��X�E�9쐕�Ӂ�i��,�h0D��W�jp��"�E;֝l�󋨂F�`���}���Y�;{;����w�W
�P):cd�RU 1�T���*憷hjU�n%$����������u؜*u��!��'�V.xa�a�r�D?����Y��trZ�ܙ�	�H�<#-|�N�
������O��=Fe�t�M]��&]�ӆ���8X���K�"��S��:5�N���K_��Q�vH�.����ąx�S��6�2�[�����GN�&�5>�<��|������8�`��^�RR7R����!�)I"�(&�!�]4��Vn ]���ڭ$��V�!<��܈��a�W�؉��s0��W�z.��n�NN5+;
3����G�zcW>��1�������&�|���q�(��$Y��t�9���Q�u%��%�%X}ٍ�!HT^��*6�C2L����;I!#ۖ���Jَ� oz�T@`��4~�5�x��������w-D��q��L��4�0/B�x/���E1�3\ؾ���\����W ��ڪu��ݒ��� Ӝ}�9���w�?wտI�H����!��Ϭʧ2�a�� ���2�κ���D�F��Ul%V�*��b�ǳo]�.�$�%뀈��;<R���(~�ek���Ȯtd�6�����L�j��U�'D0���r�v�o��w�f2� @��zk�1�ƀ\��%=�o�dԉ�C�A8��p��������T�o���e
�nn΀)UU�d�.�g�	E�Y���0���N � 䔎2#yF=P%�ZOI�c�X\�Ń?�R_Bqإ�N��% 2�����)S���oY�El��O,�T�گ6�@�n�3�@||${yl�������-O��� C�:����k�wz��*2�&XvO�Jnه�9&im���Dy��j�#g�c%!�(={),�����5�%��Xk����@��03�6 ��f,�9&|<c3q���>.��3*����w��¼��d󳡺/���Y��@5�fZY�`�O�J�Rk�x�����һ�]�1�v���rE��#(�]��Oz��Y)1�S2@s�P�JH�F�n�W,A>�X翮)䋾�I�F/'���A\��J��x�4����e<��n� �W�f:sW��}u�U��[�b�\���`���ϝ�_���Y�{��ps�p�c�����9g쏪i-T��ć~z&��9�5��[�VP�7h�0���6/`�֩(��������4mCݭ���Y�b���K`P��x|������89��#��V��
��o�bC����q�jkɔP��h�?v����o�vZ�������'����Ǯ+�����;�h;�<�?��B�p$���;o ����CE)���4>t<�a����@͐��7���ޚhȕٵ���9���������@��ǉ�|��\O`����v���j�?�x6
�cՌ¨a�Aq��Q[2����G[RB�ui�`eAf����p�.9�+4xb?n���R�9:ѳ �.>�7�d�^� t=l��#��$����E�FѾ�&0�
{\ t��6�� �K�:� >���=��4�7���8iC��v�&����V�������ʬ�M]�x'��l漭���=q'���f��-�ۯ�cm��|$z
����<�X����6��&�|F��`$;*芼�if2�P�&�͑�}^������N�����I�̽��#����˹M��_~ ���XC�H�
� G���W�ڪh�
��?�6���ީ?�}�s� ��2j�РFc[��Dк�� ����.FC�V��$����ˋ�T�=x�e룸��H��\ـ/ʏ�����3u ��N�l���M{�S��ӡV�q�M/�O�V*�G�}��Q�<\�ˈf_���L�d��\�M~N�V6���oH���T_+��⣜���L�������¿K&|4%$���fZPÅ�$�t�z�$3�J˖&8�	i��2��w�_�{@��4:��}��� ���h��G;�i�w�J(���5+�B^���n���9ʴO9U��|�'��ct���9�i��o��/��%��iCʩYK9T͝q�J��	?�����B}��p�57)�NИ�y���%P�O�G�P,��*zi��ï`Ǎ2Y�T��G;�S��^y�P��C�ڞ�uG����XL��?I
w{I���:E�zV��g�Ж�$���t����I��veQ���h5��2��vC���E��n��b>�س���	 �*e�4�	��+*�%7�mc�7*�ݦ�H�x���y�:{��y�,5���h��ь�t��N%J �&Z�c�w�3b&�A:c�:t��؛�i$h;x��o�W��3ʿ�[H<�c�<@�ZŒz<�:�B[HG ���=�7�����e�rԡ�(�r���S鸡�ܿø�j���M�"-1�� Q|֢�t���|EVEX���xϘz�x�n4}s��ݳ�k�F!{��"�ʠhc:�T��t�+d�X�ݻ����OJB�Q��r=������=�[�F�6��^s�s�x���cT,��òe�@�E�#W��7���"�Z�8<����:�DmQ�ת<�CωҥR����j��&�x62w8�����w���P��mB[�!Bf���M�@A3���|�z�tS�����.��V��B����$/�AِF��������@�"�jA O��L�`n�X���c��RZ�����6>�� �������%E���G��*=<�*Li�v�n�:J�®K4�Z{� ���לL����{PB��̈́�1�"����*'����G.KG�K���j��[E�ߛ�%���sl�1q`ځt�Q�_�(6�|P���鮎���%|9��5�sB��Ee���Q�	�o�����)Լ�`�Y�W�%�Lf�3��z��ڱU��A��=�Q�?�n�����AgK�-��E�xV1v����6��B���`Wr�M=0TNI�����h�w�A���Tdp}�{��gG��u���R��(�n�!V\i/�Y�����q)+"��FB鄢h��N3� a�j�2*W��;Yӷv��;��a�p)�{���e��g�'��`��=k��d����	d�8��B��6d��ĭ����N�{$h�W,4�~]q����?��b,��YN$j��7��.���@VA2��l8���ʌ��'�&�@u;fq����:u\�v'�6�]��%��wa��l{��j� ��'��ǔ=�����]"F�H���:gV-�^BwB0n��di�<�|۽�]%?�ᎀ8Ӕ��r�]��ě��x<�eй!Bh�zJM���I�R��rG��?ܧ���O����МJ���=�-B�WH'9y�d�|����p][�y���ը���f&�WD���Hh,sW�p:,ͱ�:�Pvu!��	�����i3k(h�\(lt�L#D�OT��d�
��(��-~j�P�Ă��wrA�� M�X�@$|����ԃN��Q����͠������DzB��5�8����]!��iU����I����˹G��3�gj4v��˄�OT�F��y#Ӭh���C��S�Pn8V���g�۬�N	Iø�`t'�֏В����0h�eq֯E0�Q�GP_��X͓����)�y^X{��<c�� ��"�8�"mx��YB��R�*�M�r������9�W<�������SDЛ�*Mm̏Y�I�c�u���	ʤ�o\�78�rO7R��@un�E�}Az<�ߣu�B	�ٌܗqd���_F?�n��1ڎ�T������e���i�>�<9�|�^΅t?��>���&Ix9��cf��H�e�]�[�:�Ϊ"��#xߒ��_{�5��t{t����¢J����>;8Ƭ�'�T�AZ��i�-�9�<�+ƫC�L�(�IҮ�i�L���k߃N5"W�w�$� %�
{�p�Ǣ�嚇7Ԩ8�R=A,�Ɨ{�SF��Wπj �pη'��w��v�@��O�d�\�i �������T�=�oe{��!�.���/�Gt���j� �kӊ]�z<qr�g���ĉJ�7��Z�h�e���[�T�"p�GܒqkB��u,&���G1��L߉U��y�k+
C���'����6�ny���н��~<:�v��N=�n'Z��X%�Z@��Ʒ�;͡S�?%���s��?~���h9���Fv�x��S�9RMK����L�~B>�ɦ���T�ih���eś�Q(��˘X吘6~hYa<�Y�A��
�7O K��"#�]�O��������5�評n���I��9Z!Hr����2�]��x���ah���|��ʪ��ڸ���?�z�D^�M��1v"F?��*�����J���d�y>h`�L�u���P��)�"���K�VZ���q�"���_N6P]��"�H����-d{�=����E�ח������eX$��2ŋ{a&K�A���ϦXR�V=Y�(s�/�ѫO�������yY��(�ê�8��\D��U�-ClN�6z�$d	k���(����S��������vl�i�f�\�Ú��]���I��Pc����M̸d�f�7��s�TP3�����߸�셹�3m���[�#YA��r5G�euH��#��D��dJ���)�,?����2J����f�[v���$G�B.� ���a����<5�^ɜ�Z�8L�uX/<M��l2��2�)3�	.����ސ ��c}m��,��7��||{8b�'���!V0l֪��IA��]��A?�7h6������"��2�r9܄R<�D�J�X�\0��*����t�YZ2��ʫ5AV�j�m���z�Ī>.`�OT�f���G��i�=������qh��o7�*z�:Gg�r����қ��n.%J�!v˩r
3ū/�����nnn�^��z�=�2�,ɘ��9�w�f�3��'DG��Ȩ�nO��u�c�x�̚�'C��Gs7�1ݶ����X@�����S��#lj�5�/G�SZڵ��|ɴ�t��庯�#4x�Ȕ3 %SJೊ$nR�-��7#4F!,��]���PU<�I�����:g��,����fA�M�:3$�ǋ*:>��oav���٣oSKy�8P[���Z$���k���D�b��7đ3k4��{kg�cWz����8	�K?����n��)�[ ����h��uq`Tkf�g�Jv�sކXx�+��>C��+C�w�8���W��1���c>�aǝ��L����@�nl{oK��z4&)�W5�g�� �d�Eү���dג�pv����+�B#x��&��u�I�����e�Yu|vfw�L{X+w3�j��3Ϝj�Z����{gv�A͌M�t�Э�(�����e��J�󓿼VRI�,�p� $C�Yo��w(;ԣ��g�z��?jǫ�q��e��b��쉠���0<�s�X5Q~�R����;�UO�r��z9㸳����/b��8Bp�|��R�-��r�|�	=$X
")���>OPk�ZH[�t�iR͡�¿=�.��Q\�zw��#{u������8�]��Ñ*wf��e2$�Mŵq�$>ч�/Y���0�8�д�E���J��ib���Y�r��x��OY�+�4�EI�B�5M�e�V��H��v�T�)�R3��;k���>x�U�����c�(ȌJ)f�z~m�֏� (8kS�[?�R����^��z.����s�6T�,ت+�,������������%�)�����U��\�y�����A�
�{��E�Zi��T�;����>��_���{8A(�������Z;dI`z9|p^r���Ǖ�DnΦ!�ilæ>3�ƪ��DO�A3��I22��H>P���z�0�����|��(�����g/c��"�8 e�Z<<3�97mR�cmy8$9W%LC��'�<�� �� �#%�SK�Ov$W�����W���H�I��S�4�>��O�$ 9��?H,ɂg:J/���`B�v�� ��֖�Wӄ��S{.8���"1-e���ʸ��D��3�q�L��/3f8�0���|�uT<������)T�)(N�.v���!-������hɟ�uhA������F�<LV�>93����B���X���E?gz�����<7�b�P�fz�b�	�)��^���i1�2k�*����Rݬ�͆��BgI� �������oƉ�B������ i"��`1/�4�w1^�!��Fni���bQgf�50T�[�j���O��Q0���nT�����?	���(������pQI>�8�CrU =
5�"sj0�Kށƿ(x�iWV�W��jB<{W`��
��ʦi\���[Iޮ���l�p�H���SK���*s�yaLuz�V��j�t/��{�R�\>b�����,��h��0�*�8���p���cw�Yٹ��qhH�N7��|Dk���L��8�AD9[�_�<�\Ƭ5��?#�c�5�Voz����	6`����`s>#�-f�gc��ut�^����ѥ~�08om�j/D�u��ɒ4���+�ш}��{�6��9_(��~2J�n-z��C�׫�BkǻI�U_6u:�Щ݄�u/��c�k�ni	�B7r���(C� ����F���c���BS��z��J�U�� 6oGڎ��= -��6��$�ۦB^�S<�8��mб0�{��,�Ak���^�c�_�]�*�1'�n�B�>y��S�xh���gZ�X�^R��t5�Hs�K�g�>�7�z�������ҫ@���(J���#���M�G�9ʠ���V��~,���2�����䬈L�#�XP�O���}�+� 4�m����d�)H�3O(߬�����ZJ#�[�v��]_92*�y�O�xn8:q�}a�D���7���m����~[I��o�
IL]��/dة��%�pP�?�h~?yC���7��ֶ:n' ���-���^�*\g�F�U�%�aH�����%�������v�5cA῾Tl�#~v|��ݿ�ϵ}�-���Q��`@�S�lV`��3�y's���밶�nA�a��WN�MȩX�MZ-����րZ��.u��F4�ٶ,o��i/s��paܳO*U���ܷ�f䧽+&��P�(��/_�����Ò��G���7�i�_^?�i���w����W������50 �B��@�pM�5."o�0J�B��Z�T(�_��uaY�X�?a7�Q�V��B�}�H*�'��E)?�C��Q���ϔA�Ʈ<��aZ^븒�|m�S��ͬ7������X�<��Rq�[?x=�/1��r�} H�Qj���'0���g*�s*� ����J���i�U����\��Xd�/�&*+�+���&�@��J����+�n'��{��wַ�g�/���,���N
���eZ�"|��X3�N�&���)Ke2��۵G���N���o�i]�!�s*�P6��sOo���O��v�?��I�z+�|dBw��Ɏ�k�*��tM�}�~8lm�m���hSW�Đ�����c8�lH}:|��!r� �2�ųf��9]�����{��[z}(Ĩu���;5@J	s��\}��u`/N�M�7W3v}�c�����xy?*�}�i��P��n+?�����	c�CD\E�D&e�@����3���XS�����.�E�� �ZxI"�\e������	��]xTj2u@�Eʤk�8< ����:kc'E�W��'��$%F���a�-Y�g=޼��ڕ�L���x��df}�&p_1�##��I�n���ۙ��/U8�{Ϛ�Y���O�f�F���4�ߓ���iz�W�d�ͮSЉ�h�6��UT"�e7��;*�����n��_��ˬ4���i�^�6Y��a�e�D��3��؀2
��k�/t+5�yCC��	����ƹ��)"��S��8�����YV�/q��B�@���"��ѫC�Q�T<p8�0�{�A��6o!BN�MҫcL1�_!6T��i���Ze�LX.=6fO��k6A��0�'s,�@X3�}�I�	6��C9$��q���w�Dn�1�+欎/y�O�`c��~��¼���������1=e��&ס�Q�C����z.1AH�$�������͝q�O�j�*����j���4U�|.V=����F��?^Zw�!w���X���i��6��o��Ӕ/�����"���嬡�����1���J3����Fmmw�+�}3,�Ɏ�#����U��V�R}�XR���ng�������"J!�t���n���c�0���Ƈ�M�uޢ8fG{K'��� ��R�&�S�CuN�iР?��]]֙p�v/�g�?:�S'`�����<����5��:�{��e�%Ju�P�^5Z_E8(>�Ҳ��W���~ �3	h��I4��48�j����k�s#��զ9��SO+�[X�LGN�!��ro~��?���D�n�&�MC�Y��!	a�_���lh���
�!@�ťRy�RT0B�� k�ҜldY�eN(�\x�ʝ�R����n��� c�����t@�yHA0(�M	�c�|SS����|�l�]�d�� /P2-�dj%T�1эh!�T��as��V2�Z�AmV�T}�c�>
�a=̡T#����h�����qe�����=ͳN�^�f@��/�.��]}U<2L_�j�v*��I�5��s�`ca.�˜B_��}pHlh�mIY	�m,.+�?��T�s��*_
���7C�T��^x�e����N����\���٘?- J�4�^WӘĢ�T�I��^5I-�R>��
��b��#�u�<B�T����f������"5��DY\{�T�u�Wa$�/�c�)����õ�Ļ���'O-��FKi���ƉG	l�qq����L�.�s&�,:Ά�5'j#�}�$��q_\������<jN=��UGݲ������⵲�G�W"�>�y�?l^��B k?-��o���vG���*�cB���~�(~!��p~������J
ݗ�$5zWd�� 5k_�\�H���$�Bh��-������I]�����D8<_�!����^̇PL����s�T�Hwv��w�k�
9�_�}4���z-�*1�3�3y�'g�-��m��1�'�IR�A��-�h-H%@7`s�j؜1ϧENU̱�_q�y|nO��X��*>Y�#{1	�.HM�7�p��ҩ'�	y�"��m6$Xd��qϳQ0�_Ôwf���VV>��1��/���̪w� mr��EEa��c���?];M�|X�V����}E�(!M�p���ȉ�_�����3�ˏH�hc��F<�^�.��O��=!���ٮ������
:��W���I�h�j��4���b����8щbi�����&�W����//�@6ce���"�}}�AV7j�����1���ͺ�k���S�wo��Y�({�r;*���eR�m��JV�m��(dpN1��3d�Ys�-o���=ǿD[=�z��J�֢��-=N/:�/�K�b	�=A��3���7���4��(�jA��&�:-[�	R��}>�F��~�,��I����Y	�g0�F�e���[	Y�Εn�,I�"��6j��������v@�m��.d�F�?FoR���]S��Yš���Z���׭)|N���{Ib(�O�&�oBa5Ø:�n<�j,c�媷�B�"��UyL)D,;�iX��uƯ (m+Z�-9!�4�MT����N�����7�����U�8.�!����8�2��O�E���SK:$:�������/�F~��/rnޘQ{�-0L�S+�D�u���c�bHmk(�<�=��%e�r��jmk��^(�ݟ{����`kuGo��vTHU�4���φ?y�z�:]D��y�2N�Ӊ��+^��~�a<��Q���R�v���g"�+�rg�[yd�p|+��Q.��4]qM�\"P����(��i�"k���4�Y��0���ЀH�|��G�(�J��уsh�RITB�_v��g5��Hh��,!6��a���;���E�>��2hWf ��O�Y+�� #����h{�0�W1��8i9[�kE�7%�>�1F����|/:WB�����r��ô�?x*��F-\��Bݺ�Z�>���N��.Lm�w�>b�w/���M��7���j�����$"���O��s��w�{����T���������c���漆r��]1�� �b�EÞ��!L �Q��$�9�5�H���8���
�W�b�	��)�|�gA���I��Ə��B+WH0�?��J�8��rĳ���z�������ȱt�w�F�!�6DH���	��^9 b �����e�Е���E�l��ы��;�]�?���BA���(wˈ�  +���2?��fk��V+�e�p��|g��Q.��9"���:����sOSF�ܓ���;�fi(��B��B���������ɉ�>�\�n7`M9cz�_���*n]Φ�dYs-�T?u�����33�������D��υ�J������-��G`��@%�/�#?���P�Z����U:�"�J�<���NJ�!6��OOn�k�	<0KQ.�P�̾�y���I8d�
�Z��&�J�w�ۿ�
��/�Y"��iؙ�Vt3�9��a*��SJ�6澩�?�=�v�+ݶ����$��l�ޞ �$V�i���D\�9�V��(}��4���g'�h��]y6��n�p�.9��E���WGPP����UnŰ�Q)��,�5�W-M��p{��D�%��RK�����A�r���e{�,k�2�AV��������C�F(ذG�&�h��t�bB| ��:SƏ��x�0�� Z	������6�	��oY������I~9�j��L���������E��ȑ8��m|���SǦ��C���`�g��=�Nb��5�g���~3�ȿ?k�Q����ev!4a�#͵��YSnl���l��E��痻���oh�n���N��<��,u����.a�p����ܿ]0��6N/�v�H��F���!n��` �b�B��g�Z��H��e�:�
=r3�bg�-�ϡ"���5w�o{��A�N�y.{Q0��:(d :��U ���e�j5Ja�������nq�&�����C�s���5Yc U�HPh�
OQ-J�yB1�����F�ϲ1�˳կ	
5j�F}�'�D�I�=&��_�0�k��	�~�IHq�����J�l�c|���A�3��Qv�=L��d�����F��q��"M K�A�+�gvW۹��Q���)�N��?��3�m#�.�C���i��,؂�
���jW;���S:2C�<���e��P���3��e��F��:�Y�j���9,H��au�/��<I���SH�
p���	��:A	d��2����??���"ѫ��d���79%tV���<F���>f,&�?Xk��qU䷦ic%���|}�
���вzK(�Q��(1�>ݚ�_P��'�@~0�`���L �b�~>��^�gɷ�����r7�4��k�[�2af͌k�a�I�U����儓o��5���扨A�_�'�_�-Ҋ�,�v���� �4u����mRc_%��b_���p�8�T�H�~[���K:��k�'Q~�C��;�T�b=�=/���cD���` S&kqCf��~��c<�G)�����{���F�>ē���Ee�{���[qo��3�?5��1�0K�[��:�W*-���r6��ê���<5?�v�����.�����*��
m�.A�ʺ{���[�(�$M�1qݣ�Τn�?0Baɺ;��a��P��\!����!A=��h�e����Q� ���F{�������dYMA	ڲI��F��Yt�CRr�CU��ބM7��ِi�ڨ+�(��ǯ)�^�n��*mמCA���UHߛR�Ԭ�ם����*��E�qܭt2�pT�.q2�����(��e��mi�>2���"��P_�4?�s�/�ң�z}��Q��;��A���;xa����c�$%}lD�qNSx�z�B�mz5��b���M�ݹԻa�~y@�S�u��.�eׂ�X�PA�ڤ�~�0���*����%�
����hdǄ�_�|�Z��Z
�J�&���d��
�x],�m�b�W$k��.�_�|�M�Qx� 67��Z���]v��р��
F/�����3���=��w���~�J˃'N3*�C:��QC��D�a�8�
�>]Qj^@�a�]��*��4�UKg���C�ى�0��������٧b"d��t@�'�3�3�����[iE>��� FP#� Z����ZE�Q4,��NK�E���W`7VD�ׇ����?Vo������s5(h�1��kM%�8,7b=�b�+x wr(aU1���G&�sH{�+���Ѡn}���1O�|.�[��%�d��桙}$H�Z�i��o��Bh$�>��7[�?TY���������}�C����r��)����c ,���ϳ#G,w8#�~���q�"�B@<{b%nA�L�,箮8+���/Wb&ND�#���/g&��m��Z+m������ٺ\��1�tC?E���z��%�<��3�aEKC�$;�7fu��&�D.NM��0:�G���xkiZ��[���(��p�+���u���u�ߥ�uQ��w�v�H�`�X�p��2�ɍ�ǗO���0�J)!4����{�\��1]�%�4������d��fe}�������D��.ef�*aa�]���Vu�L�'X�nV��_��:XzQ�i���שB���^aQ�1��� � 8�E�ӿ������t0E��[��co�,{C���¼-5~]a�D�`��˽�d��J����"G�+��:�{3
Pl3.�m�y�\��\��n�_&o�.r)�2@(�������7a�=BvE�7�}9����'��𝠶�
�<Jb�k��"B�`X�c�7�L�d�#�VS�js�N�Hd<T�3u��9�p���%jشi���3�?6�3�X�ߑ=�_$�^�s"�H���O:Z@�zLW9&l�S;��H�a��tL���1������I���o���G�Ғ�L��W�7�����W���w���"���S�eo�b�v�Ι�x����	+i����{��S� 캏$$�Ňj53&4/o&b��M)\���Mk�)Ɣ�z�wT�F�wa�m�Kh�2ejb��u1$��cB��L1:;k�Yz?��G�-��b��F/$	�q>�/�[�ܚ���Xg��#60��)+��^��M#�#rYj�>G�]�\�����{�a`�|��J�dJ���}cLr m������]�ˠ#�>����J����PWgt�
�*��@�a]��Op�X���1��,��ݯ�Yf���i'U�qg����ć`n.��O�9�Z.��P~*�{!p���A���҅�ָ�;Z6��=}��S7���9ns�����G�4t;�mФO�@�x���C�Aǫմ#�4hX�Q	Г���S�+�ağ/.�~�����eg�$^	~�fM!���ɘ^-V\�����ۙ=���C��hA C�w�Q�$.k��ƈ��	��K�gz�t��g?;\m�u����������	.WHpcik��������P�0���c�eT&�����L�9|�֡-�+���UX����x�V�Fl)F�CL%�L�J
�Htg8�=����qU�i�
�3H&ߑùK����5��iGc��T.�X�I7����2��o�� W��X5c�a�_�;���܁7] @SI���h��oy��y��k���7���L�
�<�3F�q2ͱaP�����Cs9�?��oz�3���`��1eG�p����t�q�i�����H�h�<6`#�"��D�����7�­5�Ƶ+^/�H��������s�R�����F�d�"�7pc�0<o L壧Md�x��Q�<��B=2�kyaҤ���	#DG巁4�����R�i�,�ۅ�]��[�d���sӌ���;�*}�ëIW?��X �0��\&��g�\`���o��]���Xv�z'��+�c�r-"TR,Gn�CQR����*�b������U�8;�%(k�N�ѹ��H� [R�c_��j�U:@*H��ӧ����x�]Bj���{����}`�kl����8~}�@�FT`C0�&�6�x���G�����=q.����V�7S�����'Nx�$<9���YcG!�П,�N���&Q�ٜfH�#�sR�;�S�}\�>� x1*l��b������t>����U^�{D�ޔk|�e��(O�6�]��:V�C����9� <�ǊSm�W.�N�4���{'=e>�Pe��W���E��$AEXv/��;ʗ<,>���!vq X>�=����~:�ۆ�nyG�a �!t�t�B�%�OC{e�5Y��f֍"�c!�Ծ�a�L��p�KeaZSt���OY1G7��A�y8r�1=������Xr �\.B�<�Qwe�G���+�8����iVlore!o�a�~Z����:/ꌉ�an󼅇����:vlh���#��~�d�q_w�Е��X�(M���T����}���n�>��������,�&�����N~6<�T;
R;��$>��o��?��<�"Y�g[$a��8���4Jv�Xdq\(��U#6q�sj:ahc7i;
°}!O�/Jtd�=���u�{ �TU��J%��<��֨qƅ���Q\+�ؾ>��X������X�ijk�� ��P�/}��ڬ��j��I�V�ϗy#��T3� {�Q�S<��9��e`X�4m�1��4��4xk{����	 <n���h
��R0���y�$kp-lk�l5�I��c�+<v�^��{�I�O�9BSsM����)���V���-���{B����(d#]�)��&���i�<��&���I�a�>�t�a2&��>��ݢ4o*`X8�,��nOsP& ��<)��	��̷����\�V��R�2���C��ճlK�gEe�2n4���jߕ+t
�D}'���w���XwC@'X��)�=҆,�_�ܐ�sH'������&���C����'�w/ǈe�R+4���:By5��ˀ�7�uˠ��wB�"���(���M��Џ�Tu\�8�",�)r�j}��X�Q���G�*�	ܖ�V!�08�)+��HU�@�,l焜�{83RЁ13�lj�&��t��e#4�W���'�&��&�/����ܢƊ\��|?�d;=|�!�9�Ԭ)��x���:�r�H�K�y����H6��

M�b;9�COƋK�Hhlz����P�eLa�S��B��?��L!��i�:����4-���O	�~�2}���yg�k�Z�����H�G���v��g@1T<FWl�q]��>`��}����9� Ջ��� ��/��C��=��;�&So�-�)~���:Y��r2'��1������GlH��	�בL�&3ʡ�9u��2"SYF%�i�m�������>��HM��>�)�(��!�(�Dn����>��P��i鸏�M��j��2=��dx�4]��.����k�nC@�ov~�Yl����	���#8`w���~�/��ڑ�7��W��w�o�E���u�UZ�T),r��!X�
���<�R�\1t'��
��V�7�(���)�h,������ڷ��A'�u���B�e� `�iSX���Rv��W��)���D?2F������6rx4��Ȃ �@pڳ/��C���sU�#o�[��5���P�h�,��3/t4���
;di�8I���~!��؁�a�u)�y�#^!��{_��0�|��%���A��	���ʎ�L���g"�Ju�����\�w"f�=�Ɠ㚱���7��k%}��QVf%5��_��pM_Z��q����oL=�銯*gR%��<��
�G�c�(��9N�g�[VK�����£�~8	�����1OY��
?��I��p�6Z,)v�_K.���0�H�ȍ�פa�(�(S�L��RP��%�9�E�G(_�r�&�,��.v� v3��jrS���R6����F�D�]�?�C1��2�L*��'��g:1=Dh�zŸ5Z�)��޼'��n�^��ܗ�X�k�D�*W���4` '�x�_�˨^1p*bi����n��9�eyo�r���*���{`g��e0�f%e����g� ��1+�q\zM���I�4ClI�H���L�������E�<���UO��z�L������Z�8�eliq�<;jr�#~�tA�����+����D��Alk!jp�m^cX�>`=N"���4�J�/xE�A�Ch�V&mH�I�u��r����y�������|���b��a-�?%�ߚ��<8Α�}�xq�И��(w;��q(����^����GE]��_F4T���é��e�E�����,�X���mu<���D�  �Lg��m��4B��r��-���Κz���f��L|�;`Ζ&,;��'�[�&G��Fs����n{�Du�Z49.SW˒J*5�Ƈ�����&�����<R�d�t�.w�lg��;g��f+1�ի����g�	��s=��[+��������K;	� ��w�k�dxS�!`��֣�L8R���D�!��E���i�r%�ϯ�J��2_������4����eK�^�	�����oSY��=���:v�W��ĮI�����E��RWH16r�Pi:��1�� �ۍ*�U��;r����{���NJ��ָ	����td�k�Ӡi//�t'�#��Ǐx�:B�
�8��@"��i'��	�#c9-K_t]� ���k_�W�ugI���On��i���s��(N��Z����Z�cŭ����ZL{�CX��娤6��վ��xf��������a���bm�^'!�U�!����:�[��������|�b��e�,�0���r�'�&��+�]k�bɖ����:�+�o������9"O<��`ɔ�)����vG��M �u�0u���+8����Zj6es~��7�^5��rr]�;ڛ�ǯt�3�u�i�Tu"��"�{޶�5�/*��D����ZF����t�.� ��h�GU��Y�Z���p��8��� ]��`�[�-��j��`l���`�&���2{{.~�
o:I�T�$,�٨��-��hu��r9M���� I��]�A����"�/��
��<fz�����:�\;w�eFuv���bD���g��F�g�]:/����9J�+!u�p�<�q�f��~a�����[�� Tyd� ߯�zS��<�kx���V�@� �v�|i�1�B��)e�U/d�Z�7Y�u��XR�wXQu�|��Ǒ��,x�ڿ$����}�>V��REꊷ�O��4���=\��	.5�$�������8V�����qcUp膮�� �y�VMc�`Ć��@�|#lwH��aV��l�R#���!L���"�$)��$xҫ�}��1�R2�����r)��2#� ��q-zB���Z��ԏ���.���+��h�{����(�ܡy��Z�xV��L����R����r�\~��)�'U|^���껺F�iM�Ko����.���7N�U�9&�n�-Į��|_x6�&�(��]����C�.[n%����������𖪗�<\�.�F�И�:�/v-v�&d�����8V�~���,s񄑬�I����>س竢��Y�2T��������:��ff�e��(k��[(��rm`�|Tq��m�˄A�r�ӊ�{u�M
���t�ǩg�2N x���?gE����(�
�@�x:��l}ۉ�-a�߇wlA\���[O��ˁhѨ��`��&^��-��n�+<Q(h��2Z�{���E$U�U��
=�_�����P�_ѨF~k��CWnZ�<)��9@V%H�y��6�-4�2{U`��맄l���`CЭBpl�ˍ�E�,��Kߣ��c>����`'����פ�����0'�ET��#�����-�8��)��U�ۑ 8/��f{z�r{�xg��(��LS��qeR�y.i��}�!��9�\�1�˱��A@��p��OT�o`��6n�����%���K�k�"��	*?n���(���c�
J|�'Ϋ���]_/󼁼Gi���滧�T'n8�D O����7v��!ۺ���=�[9"㤥N�ʯ��	��rh���ͽ�0�n���2�8�Ik�g��2���U�m��_����=�����b��Xr�1��'��J�w��Є�|
���hu���Ï���J�)���O
?��7��4����H�6��An�SS��Z�6�#��������`e%���7EF�㥨X���73��t��e�۹��^�����q�ʬ �D[����A�ϲգ��5�fE賫���չF�i�w{�寤������c�O?U��yO�w��s�V-{.��"�,����p��ņ�.�A09i�����������0�T-��N�&��|[���ԥnD��c��
����{��&eCc��Qk���_���ӗ�����3�"�����p>�T�A�DV�ߍ�f���忟�y<�4�}Q�r}s�]�+J�5G�/	DZ.��(ά�~��Bw%�  �E�Uƞ/����g�|M�^ʤ�&��ʋ	���i}0���`@L"h�۟��QK82��l%�zbӽ�VI�8��8�4���)���6R�2�
����(8�%�&�E�iK�V�����Z5����V[�'D"�IQ�mr��).�����ۇ�G*q�{��y)�	~Yf�r���<
�L��Ǩn�ѯ����B�`U�zU(���>g�1�%��Z.���*�u�^����cM���y;�S�Ǚ~[�����P֌a�EEV�nP~�S�N�8�P�ͤB��R~�mΦ�ED���Ȕف<�<�LS�vn�/��w�����,�:�2����-7"�%]�SJ��(z��a,���`#mR�e�>�Qv��yz�+��|TdDG���\���6��ta �*�j�	u���L.�Y��B|ؿ|+?�
�,	Oɿ�j��{�ME;h�;�\���N/nϊ�ޯT4�x�x� �I�~k�a�+)����'t��ÞI}�};Y��?P���]E���.6�67�@򴼹��H ƀ���nt�; zb^pi�
����v]a@�}���-n�KIxo�<� �[V�tmYf�$�ȋ�L,�՟�(r�܏n��mG�9����g�����e֯�D6�}��T�>l5��K}\�1Ibk�ߦ�_���	���MXIʹ��4�}����f��=���� �21�9�� n�BX�fr�^���0������>kQ��oo�[�Y��-�4�rhT����ţš��_^8K��7!I�/�=��w�����'���7�C�Ij��[��ݶ<�v�P��oi�ľ���\(\wzF���U\�ͬ�I�9i��5C!)�*Ku�3a篾�W���7��4�_�B�W��\�턛���]*�����Ol�*�Gn�\�c�J+��/��St��V�QD6}W����_m�3�6_���>n�Vo�+��ML/Ƙ��܃#���̀����1`#k�ʘbԎA��pY��RL�jxy�q��P2><�mK�s�X\�_AxWwt���T�7ߤ4���<�s�Mҟ��#*o��Z+�uA�d��o#��髗�>�<�7���^��>�>��2G���-�kԳs��=5G�I�����᣶l*�I���~���e��_�6��
L���U�PߠgC�|x��h�iOV�y[#c`��~�^c!-ۀ(�A�ooM� �Z����L�5MqАB���T��+S�f��<;��ٲX]A,�P�/0�3��mM�o�PQp��zP��,~�\"y��wW2E������Ʌ=����̖��y�H��B���r1�Z�U���)g��s����z �l&�-��}x�r�/����̓�1�m�x�>�ji���go����s�j�EǇ�Ϟ�Hn��BQ��c�1����w���?�az�2��}{ ų=1*-��y�"�N���1���n��g�ģ����Q�á��?|��vnU��\��w��o��\�_���e��>��GK����[�]M�v�Q��ə����f���c��C�x��H�rp.	F��̊u���W����t�"�#������d�5e�Y�
�2�T~�7>�tAR�%�fƔ���AM�����"-f�I�=��!rыy��>*f��&��Y߷&