��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���2�U�z�[B`�#�� 3�����E��R�=R��1��TH�G��N�����` �۠���<q��c}�޼Y%�(�"�sڙ�AӛXG�{|��AT��x�PL(�]������r�@�h=n�O�^����	�{K�*�q�a�T�FV���:`��Q�օ�H�m�Z<A�=p�Y3������ϭ�;�jHz�#D(-������Γ�Qk��c����{p������y�q�K�Ʌ&�o՗Vy��P�N�*��}f�G��g��&�W��$�R
����a��㯅�Z^<9:�G��S�kUZ($�%��]&�A��Q_�+�\�~�4�Z�:��iI��`I���E�G�&d;���;u�A���|����"n���П�d��D��+Bӏ�}��r4:җ��	���OR7$�j�P�˫T��=YǪ��'Sx|�:��W�����[�Y������$���̀�Р!�b7+�F8������ yB�E�G,!
^~��zW	ly� ��:��֬��ȣP�/]ZW���D|�jb�P�L�\d|P��	�O܊�]V�G�M�2ʨo��������)�|���p.2Ī�Mf�5*(N�i�E�J���6fi�c�d)*��eq"TuKAeb��ܨ�܈0'G���t߈�pz9?>2�e�=i���#n���(�)�9c�"y/��-�
����.��V�־���"L��dX�c�(����e�r�]�SgE���3 ɮw;�a^���j�q,;1TZ�3�L��2Q�-�XްC(�6x	�%|��4�ŭ|$�1�p2x�5��		m��8k<��q��*��c�9�y��+D� ���}�,���t
�� ��\� �7@���K6�\���(�"�ʐ����@����NrD�I�7�ݟ�̻�κ�q�Uu\vwB��5����I�pp����BeE\�{]./`+�q.	�˒~�<q��n��]�<~K�|�z깪��?n�LC�r�|�������}��4�T��|�e����0V�Q��~
���Ӭ^P��7� �*��)��N�w����V�V��`� �請�(q}��ΓR��!s�|'6�7$�E�ձb�p0����P��2�N��D�2�2�u�/��b�B�vs�P��
�%��2ِ�H�]:X��QOF��g� !�Q;�GQ*W/�o�F��=� Sln�]xd�e��9Sݎ=���W'�yvd��sL��8ڥ��j��4���T�,b��h&�
������W�;���;�Ώ42ŕ�?��o��ې�8l�2b �)���ٵ��U�wZ3��A8Br��歆�k��~˥ڃ0�p���L �t�M��U�v��&^%��K@�2a�r�H�w)�c�qi�=;�|:�og�<�:�Q���A��9��_�6�YYɔi'l5L���G�Ӛ9�a�қٗ�A�wU�d[���0o1_dK��`8���oe����U'FJ��n���~<�%�o�U~Ӌ�d��%�©x��*���ϟma���w��ٲ�f��,�L���$&b�S9_R���� �c�o*t��<���3F𥔚勬�C%~z�m?��8?�Ï�4LU~���k�/�C����%T�W#��h���:6ة�~�#�^�SR���	�PO�:'F�@b1E`<�m��3���Z��z��liQ&:���ϘC[$�/�}�*��Xş\�H6���oќV ��TN��1��R`t���
u]^�
NTp�1�T�sZ�_��Ü�"p��7b��X�%S!ʥc\v�ۜ�z�N/�S@��;俎r�
7ٿ�~Z?�:�1���<�b�Y��T%w.��ճZ�H�+�W�+�����8!^�F]"r�s^��1�烷�U�n��6��.�L0ղ^���l�ܨ��'�}�Pg�1�Dʘ�e���-�wa����B����o*$U��=e�b�������F��7��4�<��Q8��>V�C�����f|�˩�%!�}Ts��6fZ����پ�CD�����{�"�8�� ��5��U�4o���ܿ%4�ƌGY�w���L��dn Z�b���T��\ܽsn�;s�*����D��)�aR��7#N?y��װ
]����6��G�ŭۮ�`�Tֽ���١�l)%%'q����Vk2��x���Eq�� ��5�{�C�}�K�]9Up>�װ�4�]#+�H���}����� �X6��l�xB��e�a��Qv\�(`�Cn.��p��}Z&q�6-����5��d���p�%5�'B��,4z���λ��{h�'����Ć����F��#=ǵ���j��l�=���y�l=�w�T���m���uPW��o�qDP�PU�X�j+�i�/g5K|�������	���H~!�@���sLͻ�� 
f�|����fD��=J¡�A�z�J��-g"5~��N�	��K>ygy@�7�L��kRf�m��I܄�i좗�������7q��l�"��8�<k�=d&���N�}3��3�HL_J�����C�d���ֿ�l�eP��+}H5�O;��~$��T��2^���F�����Qo�6�#�J��J�?e��y��\���Ƶ�g���jT�T�N�xcz%��l8����W���*Ohd�t�ݻ܀�QeL�&�c.2�sk�y�;��#���ȫR�/ñ:]�줿%��\��/�Ц�z4%�q�4��?�P߾��0��YY�ou��C�г�9
# I���pl���Z"��Y�a�ÆS9���WW����Q[�iجyW���PɇiAo]׊_�)b�My������畹��Z�h�a���Ɛ�s�Z6�H��$�{��ձEQ�9��h,�\G�REH�Td`�??e3LVV�Q��j�^��|׆tk�s]�PqE�Y�6��ԏyZ�ऊ�PO�]:�_�l�M�$W�a�!�̲s�uLP��w�6����!�Ԟ���:	|X��R��/*��y�:����'��!� Ï�2js2|��r�o��V���QN�o����@��۾�.�,?x�n���GX�_X�s/j=ċv�����'��_�Q.��E��-;}
�)����y������@�2̒��,DO�gx�6"��F����$Ss?�����1�Y�-{�	��sr��B��Fi��oS➋Rtd�oٷ>
��Ya���U��[e�*����4.L�L�T��JZ�2�D������ϰ�Ϥa���!|8�^"�f��m?H�_J}��@�kp�[q���tO&�G�0��"���G��(�]KQ�5�sE�iW��X�4���Ԍ�;�L׸'!�#%/�$ׁ�5�X[H�ְ�J��p�ϯE1���*�
\KGB�q��bo!ڏ�+ٿ��l��B���k%u��jMau���8��pk�n��G2�͘#����"�S<�$�m��/��x�!bW����myL��j~�.Ԅ$gG����Y�`�ٗb���c�� v��<ё镔�`�U�X�4���d9�F�i[H,$e�<}��~�,φ%�&ڟt��W2����rA�dU�dQ�g�
�c�KE�(�AI8)�E��m�'��}!�fj���w�}�tO�~�ˊI�_�#V_%=�Je)e�li���ع���%U��y���4B�V��q*�Vݨ�)��<bH�Hlp��v9�P��m��=����̣����P�Y�cad��b�)��ʟX�i�mL�X���Ӡ1H9nU���͂�"W'��v��M����@W��2�5�'�z��m_5D�^ɂ좁�5�n�?v{ ��S��R�g���3E���m!��$Wޭ4��4RS��(:�s��VŘzǲ�>b܋�7|�5�����^sχ������`���N����$ʹ7�0ַ�=�ܗ�C3E"ʫ�!�j�Z3kF��]�}�YXv�W���I��6�p��3�V�O��UJ��=��b�Q4n�7��h�����*�ɧJD�7 �{4z�.���xF�J��l���O��F2���L��P�y�qR�dX��r�$-����i���l���~X�����d$��� ,���4���`��ꜝ��|F�X���m���4Ɏ�'��~.��{���o���3�YSI����j_��tu�����%���ϵ�\7����F�K�?N;���=�æ��Ji:��3�1Au��A
�M=�����i�+Ȍ�D�PM�5�b?�X ���[�#.@dѩ�!>������)�����Q�ѭv6����%�J��%��?��g���sl���n�d����u����zȻ�:é�>d�5�yLF�6���%�V�Q�\qfa� ��qQ0%G�� ����ˀ�*����A�����U���-@8ݳF�65�к�E�տ[\�ϘG@D��:����;b[�^|��pL�(�0��d�M9�����جR�;��i��.������7_�jo���&�@,�D�u���a�ާAy�=�Mb��hE�ߴ]�y� �K�L��$��)�e�zK���Hޥe��\�L�CS�ؐS�DP�Tʥ��6v'=I�u&��ǿ]���y�|f*W['��2��x�a��#ꉎ��1�큄1a�z���ѭ\P�a&�*(����B�;G���=W �;B#-mK����\.���� �mDUD�	�&L`(��d�����w*����:k�9m>�f�o�?������_z���P������w�����'����a6���_��_�˩.o����M���� �W��^�� ���#�!����h]�`���.�������?	Z�@R_��@�i�}��3�+�XDu�"��*�[>o�����<v�8��wŽX��5rH����CY:y�ɰ�����~#�.H��d�mp�U�(�b5��q<����6�n��Ҟ%�4��b����������!�(�$�ucC�}�Л�B�T�VzK>��,K���>��4�@���SD⡡� ���£é8�3p��+���vM+ád;���L�(���׎�F_M�n�d����Kx d�-ݕ*����S�)���b��/)���m�r�`����3f"`�Lk��6(.!:�>-e�E�������'4� v���-2��h�����c����6+�_�=�3$��{�4-y/+�x�W�id:)�:��2V	�������=��^	�4>�P��@�(8�����\Y�zb�Ƕ+�$����۴��`�j
��e��.-�OVjS^�k�ۮ�d`����u{Dx��z�=��9��j�m庅��>�l�݈)���>�3�B��a��0�����
��d`��|.ɔ�pwl�P��\��{�YZ@���#�9[V۵x��������
�zl�_�Ǣ
�����ӟb`r��V��7��p��aC�P���Z"�o�6q7:�I���žC;[B�<[a������������}�f�m���9���B�{=��m�����u���@��\ ƳD �3w��P�͘��1ξ�c��RZ!{<w&:��$Zј�l�s�Ӥ�%�ٙ��z�ޝ����7nc��'� �V���������P�L��v�����������v���4�F�0�5Ƶ�R�QJ��?�t%�,r�����@,Ɛ,S
�I�A�Y]����d�C���8����u�
G?��
 �爛f���~�	�̍[�� qah,� �i�
��	��>�{T�ZEJ�$��2�RnW����`Q�óuÑ�d��j/��Z ��aV�Y'䛩%��i���^������y�d����ʤ
b\�5z�o�=+HY����a�7�Fi���Ye�A�h,_��+��+R.��Pv�U���ZX�6�h���E��oA��`̵�:���S5��:m���[P��ݽ���j������8��"%t��0�k<���i����m�.�#/�.���F�}�xHqQ��Є���F}�?�ψV���[J��	>nn�UK��R22z���� N�(k�p�Y#��!�8�v-�X�f�eg{�h�dyb6j�W �<L��w������N�=��O��4�����JgZn�x�D|���qe��\|�Y����/^���@�&.�%�F�wW��J\y�\��|���:�/ro��#~��d�w@Bho��+w{g_ȉ1��5�aY:B���st�{ٕ�Po� ��[{����ub���ct�І9w'4y��Csg`.NN�|'���|�'q��_N�$�%�(z�T>����;�}	�Ci�dw�)��XC%A�0�Ŀ�5ķ���č'�P����1����O���}7H��2�Ͻ��>}��Fd�\�z��)�o�0�<��.�R�Pe�QrR\���A�Ƞ�V�e���x�,G���g-��Oɖ����܍����}�3�ޖFbx��_��MG�:CFcS�2b`��cˇ<����uh��	�]��曖 `ָ�v�֪��Ď�tS'�CJzBG4�(�B(0@�	.���F�G&�M�7��q���U��J����Ͼ���3��U�_��ᨼ[�}-�)�"s�r_�3Z�c��1>b>UvL�P���Sh>; ���L��g�Q����!�O8�3�\|�4ݞ��ᚪD�a�9�	�����*f�JL55�F+�#���C�-���*Llky����F��(����ƉHx�(Ӻ�ٖO�r�?��l��@;b�L\�!^��E@,!� )M���kL&y�����Ԋ)�i����R�;�����G�kOh���*U���=�u2ј��:���6@����l�F�x����	X�B�]�A��w݇|W���j��^����]i���=�Bn�Ȳ�����CK��h̗6�� H��c,%g�)L�i�%:��ȒQOR8qp�����H�q"���D\��S����l,vBΆB�&&<�݃.�6���:�F��6,e现������ݖնn�5;a\.+݆�-���	2�X�.�j!��~�����񐘿9Z��ǵɣ(s`F�bǟ�Z�5�`He���T��$Z����KZKKQ��8"l([?~	;5�Pc��ȸ+��1���V^Q��һb��;�B9��|uk�a ��&������#�oOoj�Gt:�Sm��i��*�b���*�_NeP�),Mnb���+�-�v}>�����������}	���<K �рý����0�:oc�����;��]p�ל7�ԛk�3P:���l]W�^#�K��F�
��-[�;U��|�hGk�~�W��t��ə�����ޯ�} ��4,�;Y<pP��5لe�������O�jk�m�.�r�D��b��1��Wmyx4
B�
��Z����g���a�ӏn!����I�r^�T�#~��Ȁ��ft�S���|竀7�ݖ<|	j�~��k�t}���c�a4s��va(�
�6��
��i�%S�+���`:�C�0�Þn�q^tc��ʹ�^y��y������g�3aFmiw%�M��� Hal6fY�g���f�����aD+�,��x]����r�'+O0JD+��n��2ȧd]>7m�R$��&��W��>�믊��s��K�u� �u���1��
���G��`=PEy�� �/d��>/���k�?��+/�ǐ�DH�~s�5���l	x�(&n�4��A�>O��@��<Ju�Wx=�Z�s��E��-}�\�	��q��2�PU��0��(:�e��z���69?F ��A��ܫ$��$��v�)��`UM�?���j�A�JwJ��`��$3���Q'+�Փ��)H��kYc�� ���2��P��z������6z��m�ٓ��o
���?%��х�V�XlY�3a�j~�W���&�c�aY��2�Cs^֖��y"Ԛnw{�� 촲{C3��知�gB1*��D0�Z�{�Ur�gM��m�Z�B�S��E�_�����1�
�¦�y�&��𢘌��#OT�I�?�BM|���?�	wchYe�H���U�&���^��^�c�dۏ���N#��]T8!JTK/v�."��5�|������޽	�Y����v�0�%�@��+Xh�Vf�$�n����ٗ8�� ��|��/�tE�2;�2vC�Gӳ:wL�����Qe	����?P��{�un�P�G3���gnMΓ�n]^^!Pet'|���ː�o%���q�������^iA�O�����."y��BI	�ѳ0�p��s�ذ/�]:�v�Ė�`��F����`�8#J4�5�sp���p��j_��k�޵*;���GW//��H�V6�����h]_:x���Փ�X���ol�5�Nx� L��o��� �p�F$b�w��n�D(ϛN%^�+���_���B��t+xm�g�J�քG�̗�TVr��nĶqM�2�4s��i��h�Q㸼m�]�s��e�Մ�G����)�o��Sj؍�$���I��`>�/�z'�d���ЭK�����tQ9t �a��f�a81�B�G��T�B���䤰���At9�4.������X�ڰ汣�b����xl�)o���^zsWv�tݳ��r�{D>�xN5\�H��7��n[;��[��	P��!4H(�;�ir�;q
av(R1�u������7s��`G�������o@> 4�fP쳀z�gd��0�d' ;[-�-u�玒i�K)IE��5�RDʕ�	ah�`�tz�s������G����F����-ȁ�i7����?�勪�Z��{���"J���5��[��� ���ޅ��O9����"c&�$�$�k���9��3��T�!]���ˍp]�#]���q���/�	}�$���Q�Xj1Ľs(2=��r��H91If���*��I27���K�ߧ�G+��7f�x�~����F� ��e7C5�um�,v:���r�<~[�����L��B-���o���e����:��D�ML!�_i1e3gU�,ȵ�rJ�8me=��iQ�s����m��,��ړLqJ�p9�r�}�ҟ�E�ZB�P�ʹ�:�~!Ћ��ΞJ�7�{���Ȥ�~l{GM��Ap�zdmp�L�G����*E�K^y�x��NE[%T�"����)�)T(A��< 1m�l�=�Ǥ[^9twL~�<B1��J��u�z���ˮ3��j@�
�� \kΒ�,[���@ �����,���p6T�����s��}��UQ��� ��1V�#s.��15}R�'�yS� k�)��x��_��HG���s�M���N8��:�BM��fej?��{�N��P���C�0��ͪ͋���׶��gX-b�W	H�1ʐ��ډ�=3mu��������>9Ψ�� �<04x$�5
�~��I�n�����t<#Q�$�dJ�g.3P�#��{��$�nJ��YHp�� ���O�i>tx�������Q����uGDr	�\vOB% ^�:t/�ڗ�:4Q>	�&:oPl4>쯬u`@�fv6�F܆N|���������r��=�{�z]pE�yg1'i-��D�E�8@O*G�8��>�(F��įV��ӕN9�<s��Й�������DQ�V����vR��x�]}Gf�2߾�e5�>(�g����\���!�m5v���Ux){���&Z�0���_Km�+����}@'�b�ҏ��+4`ު��I���Gb���	�C�sF8|�aϱ��-��xq�(�C�M�ɡ�r��;�:����UT�+\Ng_#S]��_��^��g�FO:�0PA��� �4�L�]V�F����ǌ� ��}ɎJ��^�w�鲄i�4��{�#  4����l��5LqV��%}��
�Dko�Z�ݜФ��������7 ���m���	h�i)C?x��6�|0�<q�XUlPrї,O]�n��_���(��Sb�RI�N��W��]�Á8�������婞Y���sXU):��\G��n�{��'�mg��Ŀ��� 9�����I���F�U�t�NK`o��A���{Bi@ԿGRcΒ��>�y�q��0�B-Ѣ�����,��b�s/��UHR��}'���^��j��CGG��&�I;��(GA�%��]B��{|���PO���+Q�����E�~:&�3�Ꜿ�Sު��^�x�y��L��B
:Jɷ�Ey}��N���`p�(ka3k�E��*
���pmĤ^@5-�uPf��@��H�//��'_��T�Q'�����K!�LBg�$i/�c���"�}{���Ė�DW��v�Ǜ���Գ�z�kYiT��?�q�`� �8�w{/���Di�R�KH*��9RSYT��8��8"��W���I�5�=͑Rҁ%^����: ����6���'5����w�CX^(t0�� ���I�j=�=}Z��~u��,r�s����>�d�A��ݴ gv�Tq�4��N\X�*����I�ƒ��ٌ"aru^�.��.�����#���J�~��M&U+��N�5?7��0�U�<���z&�~#���� ���X�t�~��0������sX�����<��b�	�蕜2i+ts�J�A�1Ze-ޅԀ��"{�����x���ޟǕ�W��e3aD|g�����W�'f�Qmϲ���ocݩʣ��׆��M�6��
��)�E"��Gd70Q0�f%�&pӖ{�R���5J� ��=�(!����P|9C
�]���iB1��3��I��:� ^vcES
����.T\A���G��P2�	��R0:L���i�!/Qk��^�24fY	�����w9#��eY!Ӓ~����H��^�!�q�kұ�m"�Y���:V��.��E͝H��l0?ڞ�8��s��=��"�N�9e�1��f6{^1@.'$(f�.f��wD��挚]�}d���U �K�� ��N��1����?U�$q֭����1^|W����z�|�4(b}�3�:,�7��ȓ��0s6�+�Н0��˾�9X;��<�d�{�����Z�)�����E��z.�"�t���B����Z���I��5Ah��ւ*��<�����A���	]�S�FfT>3j9�㍶�nt����Չ��)���zAw0�Rh&KG2�����̲/�߼R.����8�T�H��5=�)�Y���S�;��z����EOW�����2�Yn�����kT]��-�[�T^8k�s����ĸ�z����~̅��a�T��,�ë�p�"%��U��t;y�V����l���=�Q�^s�	����>z��E�!�-����O&܅v�����V�4:��߷90љ" �>w�Ν�Q�ɇ7�Ƙ��I̽J��N���ɖHsZL�x|,z7E�J�u�BB�f�xE���x�cS��X��O
�1�_
��2����H�&��E38��(����+�#zf鮯�g	��vd�Nv ?��K��zV���ɠ��v�Db>@�`-�3�D�W|X���q����бゖW�z:���-�c��Y�G�j�^-�I<�X$X�KU��eT�����
�!�����?ʫv�R<H%�雱�����ߨ�2����#<�īO�����碪N5��Ho2q�5\JX	��^j�@��V�Ħ�.�����(�X�Z+�Xt]'K��2�k=IDKCE��:���
�b?�]�,ƫ)�+�t����ks)��Qb��\2T����W�v�Sԕj5p��~���o �r�F٪WQ�j�F�]�c���yy�,��5<Z���u�7�k��w`���޵A^��̒-�1"���zs%���1�ӛ�8�JY��[�.�N���Z,H�*+[dZsc3��RkV�
���Z��H{����3�˷�(���X����t;���E�Q���j)�܌$��Q���e.�%�Vr;c-�0����kY����m �9]1��%!��{�X���]3Y�H��qwf�bW��?������?�C��)I�v�p�7F�<� lZ׍�#QnvA%�C��	^\��y��yg@)Y��/X�UR(����|��n�SR�l���R�6��T7�Ա»ӕe�d�&e_�dw�(z���p�0T�<=گ�v8(U�l����]�n_E��yg��Q��R6��a�F���z���%�6 �X�&�w��7��P'�¼]��
H�<	���$~W8c�=��T�~��Pn�zIv�f�I�8�p�(FY�^�g���](Dm�!0ro��݌���3;���]z�?S�	
�[�x"8��K��3�O�[E<�7�:��������˱ÿ���.Ө,�tH�� \j�Z��%v��0�	��4V��$�?����"o�v�I������Q-�h߿��&�S���:w+XR9��e�閚�Yۯb��p���4����y�Mv$v���L
V����<3A2�O���^PX�ˊ�Q��e}ۨ�[l8����G�\��o��d͎G��_�S�՞A)H1 ����J(�$��~�nϳ��;i4��?��"m��)*����Mg�!q��L��6.��[�?B��9�¸r���:��䍢�U):�n�|Aj���/�L$4_N��)ֶRGXuڲ>�sNn�@?i�n��0E���9��q��/$@�F����$�R��6I�(���� j�dw̰�V���f.,�2Ώ�bYy�Y¨%[B�|���k���U�LON+#7�/����eD�$ak�1�s��b{�� �4��&����Es��H2S��TF��d��H�eU���1����4k��M5�ݴ�$풓j:4�I�b��R�",U-��7��lcg�G{�Ҏkr�Y�nD�u���"����������B����t.����T[�:�F-�L�/J���P����D���\�����4W�hk'E�}ƍ�����}4R��Cf�0�M~�1	v+��I]^R��!G��,'�Y�@�>���,������*Wϯ��ulH&����0���?g��O�
ܛ�\iP�� .��w~�h(�U����A*��^0'to'��霑T�/�H̬��_Ҹ~�PZ�`���U�ڡX/�D���)�ZI��cfC_��1��6$Sd�Pb�W���8�آ�9A�]!�<��?j��aL"����3\�0� ��rV(�س��e�k���,HI<�=��c��z�� y_u̪�x@(;��ܧ�xp��K�8�z�%�������@ ~?�2�O.,%Vu��N{H�hsμ|����^�/3	�^
������¹Lq���d:Z���f�����0����~�`TY^�u�P�;�"���WY"�P�\ �H���A��Y�[`���e>h�a['���b$ ��h�̛�ޫ���D�$9����d��.a��)�?m/��1_�z��ú6�b⇸�f�T�l̔��`b�ͣ#�z�j��i�b>ͼ�����Q(鋐㙖60h>"������0�6˪L�*bg���2��P�,I�͚��S � �����N҃�����-k>&I�
M�����;�i�"��s�1��]B��b�QG7��&������9�Y��pƐH�(&=}��� �̱O0���nsr������$��`��U����m��6�\��n
�� X.SS�.�����ָCgX��e����K̄��8�b� Uҿ%�Tҏ��Cf��nFms(�"jx^i�W��6X��q��Y^�&.
�D�I h��:���؜yD��{�7lᅵ���˘��f�L(8���70�nC��|�SeD5������'�C�Mӿȓ�Ӂ�����{�y$I޾��K��٣:r��Xj��aI���K҄FS�E+���u����w� �i�vu� �i%e'��̮g~%-��>.�#,�=��N��H�V�(���KS>�M��#��͹��$���\*&�ߴ������q�6-;Bօ�NQ�=�k�������/�X�m���v�=6J��ޗ��T �8�k����^�J��W�WR@e_�����`�~�׽��j7W��1z��Mg�#������Ib� NN�GH��C�WLbA���b���Z�`���m�4�#�'%.�&�wJ�P۾�p��cwέ|k��k2���\Y�=
\1�������>��ZT*
e��$In��r𶯘Nb�_f[�}�R�q�5���?������'{�ٮ7璡2�w����CZ��}������l5&�]��G������0�1>��w�,�:f^�e�.{g�-ɔ�����*��5��L�^=%��̚P�n����k��$ep���jAsc����]��p���*�)G��~;C_PWsB��hO>�#\"sM��t�a%�;fD��z�ؓ1��W�=���L)�:8���&A��V?
��0�t:ˍ��*z��V	��Ę]�$n����v{�o��m�0�su�5A�.Er3�iIj.�g���Jw���Kz�Ga�V�3�b{�'<?��f�6�,���r'ePnl�"�Q���
T{���9����rY�_��&��,:���)�X�nV�f�$5J[%�C����K��3~���S+]y������+��	BAU����@'�DHXq�΢�H�:���&��91i�W5�k.2ַ���N�b�2�|�0ܙ~0�Ѡ����:{[w���R_�p�
%�)e!�[���"�Ǔ���j����5�p��=E��@Ȫ��{�}��m���&�E��.9$
}J�)={�կpj��'L���{60���?�����S(�$�02�1S< *��񩹻�'��3f7�5����]���	KO%��X7V���M9�� �'/ˆ56�E�KG�݁���<��s�ff ,$dנ���3媥}c=n�׆���!ug��ߺ��Q�����$If���`�0mpݱz I� ��~^����i5ɲ��wr���g�v�v�b���;m�`�$P��|e{��'�?"��5��]�`r�=ԃ����ϲ��CQ����h9����R�4k�%$'�RC7b���.�d�0��0~1��HPo�2�3����YJ��ՠjuB��m�#0����=�pa���$��|`ޕ���7$��sh���̨#�&uWU^�Ť�u�S�QuR�i@����������|�x����P4�S,m�Nv�$)^(ֻ���y	��iJ���
c=G�ɜ�y�٘a2�f�#Lx���ء�%�f�/�1�|�7�[;Ojж֜��px��L��'�a,�2N�|C&\s��Tg=�t��� cK�m%��زM-�]�>�9�ͤԘR�zQr;:��^
k���	���o�i���9`\����~�e���X~0���җU}����D��A�,��VzyF��KsKR�/�{���iB����,��p�75�'YmWC�d�UZcO6�ɷ6��֦�쮉�ɫ̹p���7�ə�<�7��&�;;���on���_�@-�y�8�\�e�e#;�$����)"�Wa�����fe��o�}�ɕց���e��&�v8�J��
bz��V'�g��&��< ��JO�0���?��M���DhS"����F�-���c�N��.40�
��@M2�7�4����ړхoBq&FX�3A�[��T1lT3 �;�О����B�Ԛ�S&|p,>"qSu�kv��|!�h d�옙����eA��ƅ�MMB�BK�G���e��p>Y+yG��N^[�I�0����|�m�%f�K˒�~��W�����.�Z���{(FI[��w�����w����P6� u<�s�6��v]Y,�N�� ;�	��^����<��\"��J�	����ؾyY�fI�1V���%�n���9?FI���n����c�`�$�}�~s��K������wi�؋�aڥ4�P��?�up�:��ej�T�����f�&�<�`��2�}�:��5�h�T�Z[�8 ]��>D��� �#�+z�x1p&��gY�����g&���9�i������5Q�f7�t^���/�^��g�C��w�Z��I��c���
m��ǉ��Os[馄���S���Q"�-�K�7����a��:#��S%�l��DHX��'싀���|Y,#�1�a zT��j]�Ap�I��w����ED�%�S�B��[3�jl?[���a��4rV�~��I9_��b����ر߽հyYD�M�]NE�)��i0�����S��T-K�O�0h��j��#/�7�1�̲��-5KȠ�7u�����N8�-���r��2��6��.�8z��7���0���r;� Ot�]8�R�4�g���Y�_�Y>5�����h��&�N������	6�:e�b���#�+x�+�kN"@X����L���-+bM.$����ny���SW��޲��ҹ�#P�|�Pl	$���zu��r=K�mb�Tq?��](2�	�"�+w��4	A�e��� �T݀��������PZ�x��-���
=;l�	�����${������Pau�o$o�h(�,�,?JЗ;)@���k�.���Yuf����TS���S����Xs��MO�U!����9���j��ZufkC��K��Þ3�P�����#�篼�ni���!�0��`���˺�N(��:��z6�l�!��E�����h�	��*���Ņ����5 �"�^�N�3h}�)y!�+j��[O$^�Ԕie�I�P`� �Ǔ�B���1�6k�tM���ዘZ��%b�_�'¢���UZs�S,
��|�G� �,J�Zz�[�]评�݇��p~��v�v�ǳC�JF&bhN��6��d�w���'����q��贊fY�jۘ�t�X��e��oܐ��ڧ�Be�q\�#-[.j����c;��[U�a���_���y��FŨ������;ݿSHM�خ���KG�����̞@�=�I��l�-��I���8�� ӟNS����4�?8�k���tw}b�s�0�����\�$���T��D3i��/�
��?���㗵1O�����%4��O���Lk^��֜� �f����N"x0 "�SؿP�QK�[��o�r�cF��Rd�ʏ�	qR�7+�:���x7P�e���M卛lEC�vނcQ�|׎Ǔa~*$ԋ�k�I��J���AUT�����8s�r�76d�� �Ѐ�N�n$�v;�k(�%}��i�mɶ�ݏ� ����N]5<`V6���@�L�(����X��9����! ���| �Zy�u�����j!�Ң�~LDp�(8��iu1�K�p�X��w�s�*�f�ʡ�|\m�| �7��A�>[d�.�)��{u0��x��R��Dr�ǐsm� ����E��<|
���.�{��8o�f0X\� �97�ϥ���q�Ŝ�̆wRg�'Z:_3�N���z`�	m�w�Xu<T�2�\y��{Ҹ6���2\xG�V��B���2`8�g�u���7�m��Bf����tY��������fA����J(�@���V��̏�+l~�q`�eH�hb�h�I�Ԕ!Ԩ5
�kP-��MC���{���8�|uh%Q9�}K6�V={��M3��4<1K�8e.(+|��^I�r>]@2B%��
EJ�'b���с��ճ�3��\)k�R���@�=s2G{�����Qj�ڱgz�������|�{v0;��L�l
L�SH�H���}UtK�G�D����^j���E}�A�qy��K�گ��v�6^�N�n�+��Gs������P�v�e2)!���K��JÄkU`�;]�[ �܋��6W`�XY����L�d�����S��G�(���1Z��U�\����a�jX�m����T�*�fp\湔io���ؖ�g؁Ĭ���Kҟ6h� �*�bI����.̑� Ɇ���gO�F@����G��nY`��?���I��S4dY@r�S��`�Fl�����u=R�Y�|����U�h9x:���9)�c���R�o}���)$�ДDH���)��tmO���N
�2�eQ4�ѥ��j��z��.5��i�[v��;�9@�%e�=�I��w#hGU����tH�>؅9U�0m^���ݑ~���W��-�kb���"�����q�*�'V�	��p1R]>msW��H�U�����s�x�"��Ҏ�W���1M��Bd�q<�D����.�6�"�+�'�d2��ϵp���z�ٗ�[�6oK
)C�gI����Y��Dس���%
�y;�L��#���{��d���|a�q�e����<>gF���.H��R[�����?�J�+��M��v$9�e�`�ɎO_��.&@��w�k���1�$2�E��xΚ�w�]�K����՟"�϶2�t��0)�$�(:�&�!��?���ژCN�աrH��8h%���zD�"��C(.�S��\������9 *�V��*O$t��[>�Q�{�����D_8��˪�ػ���_�UJ���ʕ���R�5�L��*}��C�B�)e"!g����cW8��MIP�%c'ڐF�@�Ty�ȉ�l��:���(�Ő��q�9:���$o��N�ED�s��W�I����L��6M��`��	׍>ˇ@�"�f���'orBC�
� y+N�Z$
�
gY;x$i �(��(��O�J�L�e�0�+Զ.�Y�7��a��$d8���L}�~T<�w �ͱm������b�U��<�ɺj��]99�P�9kxE�|�C�A8�>�P<>�O��8.�Hl�i�+�n?���Ғ�a��Q8��yপ�{��"寎�_����$�Nn���#��OS��
����U@z�0ln}�=X�:ժkFϳ�z/e������I�*�0SM�J��t���ð듇=����AdS���_nƠ�w�E�������l���� �H�z'؛pO�Q���Xƾ�{]]?���a_�����	���6Q"��0�"n~1�`�����n�tBs?����F%�K*Vx�j#�?x�I����Մv��t_Kr�ׂ�����"����ka���$+�8���EqLW? =P�ى�A�+)�o�,��s^�����O��`q5�����O�m~���y����]�� <������A�,���.���$�Q}uN㕏�}{p2���`RVa���h������i�V�ę��G�r��� b&?�"�@�0�ϣsn�� r[���A���m;�>X,g��з�h�ڽ�NS%��a�_�
����U�ʂ�a#��݄g��> �N$�8sh��Q�uhF���^�:���
1��!��Ԡ�֖<RՑ�h#��M��7I�鷱ecY3���Y���9�QT@�0�+�J�~�S�ԣ�$-��α7S���]O��%K���6�wm�E����Pϊ���Fz�����:�/�^*���I�puj����Sm�<A@;$pѕ�k(f �]
]c�'�%"N���)U�ZK�G�'I�Z{gPM�I�����l�4r'���.�P���U�0I�>��?*������f*o#�&�?IU����rǋ�ߝ�U$��ս����0��^/'.K��yK�9�U/�q��h�B��>{f����ǀ�w�ДM�����B�To#jہ���kgȢ=�΍��uT�R��Zg	�2�[k;���y��Hh�A��kc&�8$a.v�+��J0]���u�Z��rF@4�s��U�}Q��#��0&���X���s����Zr�g��xJ8����rc$;�!��0�l�i#��p�"Oq�/���{�W�S�#mq��|�a�Ҋ+�k��S���&�k͆���XP���>7V"���r�����%����j�iZj��%�j@5%� ��	�>ά9/,@<O���(�2W�L8�2_Z�x��
��%B3������%0�EsXO�� ���5�Çf7k�7.�4�9n���/��i��lL�u�5`�����o��)@�cN5�]�Te[��'P*�s������>��'/��7� "X�5���|�p稜Z�93m2�٠�{�ȳ�]�O�{7¿MԼ@��|�놟,E���]�~2f��Rp�q��_T���e����(̕�x����/U���P��6+��i�$��_�6	�x��;*E�q�ucX'H�@�ũ�q���r>��
0��hH(p�q[<ӧ��E>��'k����I#q�͍�!�;��b���}�cE{�L]S��}�Xl��.�t�1�1c�0���X7�ܧ����{ǥ�0��*r�y�� �J,�ӌvPFB�9Ƽ\q�O�
7��x�^�a:>:������<��Ao"~��MT�-nte�Χ���"�7�������Vʬ��(y�0�qߛo�S\��eÎ ��&:W*�ܹQ<ue|����N���l�*��� l��Rx��7W_��;���ɚ,��@c��'>{^�lO-�����j9��e�Y���g~��I�W�0��y�j����H�Zk��=	�QR�pen�5� �н�m�e]ܽYn}�cw����f�pڥ��&)�)����;צ��iכD첿�ӆ�e�Ś���i���v�ݬ��C$������_j)۟©�i�f#w�,ұ6�k�	p�T�1�bU��:�5��y�u0qyP�'�$�A�tN'o�����_��Srr��w *�l�5|�.��	�?ߴm:i?��_6`U���t���kB���+�Et�2~��%K�����
Ȟ��n�mVy��f�s'��I�"H�ƷB��,�jJ�4c����\G��T;�I���z���'`��̂��D�W���gv�m���}� .,����JB��M�ޖ����[E��h0%S
Hw��$��}����k:>�o�TN�l-8�,h2���p%�bW�R� fz�<���1�yd�c�&��*e+9��N����T� )�y�x��}�{�4��U��$�X���A$�GV�� �G���y�����v�-cy'�6���3m+�n!�����Z��3�l�M��K�fp$8Ʃ����3u�(z$���S~@�jU	Li��p[�l	k
�B���m5jVӏ�����ǜ;��U�l1pd���F6�ѥ%)������Ҟ����u��+��%��Ě}���P�̐��g�q~1��e6aPT{۔�� �7�SJ���W|l=sb�FgG��zC.���?�G{�J'XS	_d�ڜ��V�<�4�㪫�lL�����a�^��wJ���pp�/��ñ�(UL�E]m��k��B�>0.��B-!k�]�t��O�6(74GQ�˃�1B��G�G�>I�fy�WӖ�S"�����#��s��/�	�`��gѻq9���/���Ƈ�T��2���`6Z�QA��ٷ3\��m�����xՂ�c��9h=��_I�Y�L������]F�%�#ђ����,%O�v�P�|`!&w�zđ�leZ�{�kk����4i�{�턕,V��d1(�D��	vo�`uS��X��i�Fr~n�R�	���c�x���H��2�o����z�����o���>5�{�N�9k���oZ+6�����u^e�m��=�TO��S�g���M�ZÔu3�W���3%�E���}v�i|ܳS-�O�f�:�˷�~�[�b8�x��T���Z�w68�_�A�HYAulp/-���0d^dw���L�xΚ���i+�k P������S�$' 7Fʻc�S�a�� #xU:�讹&Q�r!j����5.�1o�f����ЁE��I]�3~���6n��qgz���K�E��l�R�-g�<�ɰ���5�>�)����|��8e$���.C�wkjZ���9�O{�����?aA����ҋ���Nn�g�$�j� ��i�̗	�����1��Ip�!86Ͽ������ޫ�h�aR���o�]W��|��:��bY�Qaa��I�����T�Qȧ\���Bg&�
]������Y�q�Y��R�{�z���P�Ԣ»�JV����(�����C:��H;��0�v�h,+��u4�Sm7�xQDbP�8�\��Rm�b���@�PV�dy(�ݕ�K��Z��%"�7c/�z��y���Ox5��H�3{��¼��U��p�↍F����^C/��ԠR��"�LU����C��"�-���������w_�✡̈́Uj�J��Oe-ɪ���,L��� �����L�l���P2#[<�{W��x�vp-�Qqrd�3�s�h���/B�{�{�I0��J�6t�8$�%'��J2�<���*��u��W���Z���oH"�k7ĕm�����լu��t�s��x�q�,2W�hr-]�V�3�8�.n-fxs��oZ�/����BB(���������&`İ�VJ0������+�,"^qG�13���� &k�q��}6^���6O�w2���H/�m��$�܊V+AեF-���l���OA�����alf]��.�U�N�0 I�?�����7�J���9�|MwW5?�2��y�1�v�wܖ Q���
v��,�:�W;>uG~�ю�u�b�QM蛊啠 
ȭ�H�v_Qn��w;`���x�A�& ��ϿikJl�������)�ccK=J�2��Fa��n�$�;���ߔR-8��D�_	~V��ޗ�\�9Ӑ���w�+�v�/E<ǭ�D��\��R�sr8�0������UW8�+T��#nJR�RC�$��V��<[������ț")���t�#Y/&�Ի|�Dw�u9�	������V��e���oJ$[<^k��o��E7�����oRH����}����rT����1��������}�vJ�J��%L�5�--Ǭ��\X\{����^ �b����]�\A�z2ߙ|&��5�~�����;
�� ���P�����F��0����v�װ��Dh����Ɣ����(�6E�ʀ��Zs���d/k�VY<�Ξ+y*{w��+��!]����9L�|ށ���׆/4>6�}��IM��,<����;v�9�I2ۏ���!g�dز*-�d&1\�u9���l�VS^�#Z���}|��
�<���2@��lv��G�y<����� 6m޽UrwS���GҚާͱ���pK�|@V�@�����#�;^
4�	�R7gi��.�l?�%)��І ���.G`�_�J0�_�`�.h~N�Z��`~��L���kϛ�vҭ���2F����4 �u#�=������p�őu�9ģ5T�~�'�vp�kh]���80���|��fX��8���f�HVy03\�F����;<�n��6���0)ꎢ�����.&�Ix�M8~��H��������Ts���)\<T�{aP�	M �e�t�&g"&�CF�	�[`)'��M��1�����[��<����7�G}�]!�R2s���lpxa���1F̡S�?����Zğ�pP��q?<��=��GM�<�s2mC"C���V�}[���!w%��zO�W��@ug�����0o���4�.@}�5��"Cm|"7di�姭��82�,��[S�`��p�?:3/Dآ.x�=+|`+�A:Y������ezN�Ͻ��دs��hd}C������� �Ea� �,�x"vĂb��<�a8�%�G���d2���^P��%�� ՘�0�����xַ�Y�d�2N�
�ۃ?o��iI��ˀ;J���4�,&5��d�i�I��&�e�0��8@�K�~��K��Բ��l���w�
��p�r�ht����S����"n�s{� ��3��@�"2[��Cpȼ%ck(̩�[�R��؂܅Bs,�;6�J7���&��8��AI��TI�>up�e��&.d!�Ʌe�����}y�y�D�l��Z' _�F�}nl���I�Ҩhc��F�S1�2��>���#�	h��V�m���fz�!T�y<��O��ȏ�4�(X��mv��"���B��|u~����6��$\�5g�@M:1
��P�+VsGiu8iE�=�to=���lB�~ E*�Օ6�M�O�>IS}��N#����2!p���Rl^��CI5Q����SV��rN&R�s@?je�t�H!��)�� ăG��&|U�.듐I����q=&g�S��z�Bw��q�*�,��T�+C��l*B����4����2���k�s��sG�X�� Ӝ�����
?��e� �|���!-���d�-EL�EY��t!5{ɲj�ǎ#PY�@���To�c_����S��|6��?����>%k��s�<e�K�_倐�>��%,�C5no����f��@v'���!�K����ˈA��J�M�9�"s�*�i�'�ߡ@���种ؓ��R]y}l���i������Z#��c ��=����
*8��#OO�磵�'��y��c_m�/��.��l�ݔ���皙�:���%a\]h?��Ǌ�0&l�ܐn�=bV�v�l�G-gN7ool���%��	_�l�m7R��viQ�j�󾧉T� ~�Z�́�|�������p�w��a��$������VO��!��(��L�	j%e[�D�Ƴa_%��rI1F���U�+[����Ǘ��k5��k< �5�f��s�`���?�
V;�gB�B"^�'E�C���<I�J ���ľ"<�_��6�k�"�%E�Z^YƉV��Ѭ�Pd�y�('D��^��؟�?��-k>1~�X����I��\���"��T|7[�?A����l�mQ!�pŻq����|˳%Zҿ���(��j�	w����8�����A�o�r��5�Y����w�;�3H��w?�2ܮ�z{���1K��5²D�$-���urpÿ��[���
��Uf��I+4��Gu�{�tP�Fw4�By�h�w{,;����8����?�� �=ͼʲ�&�G�����&�̠=�mQ\_��;�X��r�F��D�=��/q�!j\��o+D*1tZ����T�^��෡܉=���˝*�`�|E�'�����M�@et̹����,Iaon���Љ���`�*���p#{���@EtG�ֆ4�
��Ut1%�<������>����4���v:��L82Xw�q_2u����1�(_��v�8U��U�7�/Z�̚5����:�ӯ�ܴj��/�FRs0�3t��Ѽ�x��"��j�; �v���/f� �PHLTG�W`�mP��6FF��d�X-d�c��/Y=���Q})��{84��v��l\le�_�3r����,2e�Ź^f;��Y��j��I�q�T��:��&�P�]ɕꈏ:#�s`�&�pȶ�a��������������u9��\���-���ˍ�9f�I�9��bp�_��O��:��;O���j%����Ź�v�8\헇�v:��[Mݒ%bzC������[��ƄA��"���^F�
�&�����<��%Q�r��C�'�Mjat���P܉���ޑ��-�k�����& K�]�q�2QF�SD`1!e�{7v�CyC�|�U,$\}=�8
�b4)m��u�+���^o�8���W���h�BΈ+�\	T��jR%1w�ω�d��S���M�d�h��b ��!A�gp�����H����-�p���bS�1+0��r��V9�j��##�B�w�2<ז��dBy��Do��H3�%L����T������;�H��] �_M>
��F�^�h*S��ΖD2���d��vǘ�TVO��/���(��X���%=�g��V˚�s�>�� ��yoZRx�x��4�m�
�^�Ta�� ���Wz~�oJ~�Z��Q�:�)�uǤxV��B�B3˽�}�b+Q�J�J�W��U{Uh��*P��@�O�S��u��&>���i�E^����K�e��Č���UC���`�kP��6����
��s�u��!�t8�Aƅ��#?�j,��qI�dn�4���j���;q��E<��8Rc��>[?�en��i�+����j;*a��X�(��P��o�������Jޒ���ڎ7Y��xҢ���"�Y����wM��c?�Z-�@f���ժ!�qUڱa�`��T��/�X�jan�[��ZsO����*�����c��(�/fW3�H�gW�E��9F��؋��m21�;C�����e��y4#'n���==�B����W[T��\T���{u?��覭�d�^#q]��⍓��j���o�2�+����Z�45���/����!�?�2��u>����Z��W�MHR>]���4��!ׄn�Jq�k�c}��f�,���0T�l�M;Ϲ�H�mt0�u�<E�PH����H�Zg�E��'&gG�d�"���5�2�B��'S��RP �c�����3H�}2M2��u��;��A�Ֆ��	a�5j�N�-5���{O���K���%9Hre��e��gԩe*�Lr��á7��$������c;�W�y�r_�$8����4bj	#���r��()?�Ys�����GmPP�B�9>aW�xo�P��u_J���3���W���Ab��,�k���4j#a����ؤʗl�L*�EL/ƹ>���~��g�V�=&�l���GГ��o��r��h-�������2,S���)�9�����+�IƵ3EM,�#&,g�u+�5� (t�K)rL^q��_V�$�Y�����I�n�\K��H�~�)��R�OG��eMUN�u=K�/�r�Z�"���:LV��/�?MB�f����E+��'R�����(��sw7�j�*�?��Ɇ:U�%V���>+R�e�7%�u0�1��G7B �ʪ���99�3�:�z��L�pJ��'��|
�ƍ\~ԋE�t�C���F���q��NO����nY���z@�e�-Ņ��i5��yt��1�#�f���d����#	�p֍�'�ojo�~E4�ȷ��W���Ǉ{����	��o7���_3����k��N�A���S�y�v^�b�dN܂kZ��#��<ب�F獭)Q.!9<�{��8�A9�e�4 �>��"���K�M�r��,��ݾ 	2�N<Y��x����&qu��HEA�b'��
S+?1ṳ� ���v�����^��Y���[��̈bN%�s��0���s5;��&����j��*�g�0�(�3*���g6ӯ�q�fo��.@�e�l�-�jU�{�D�WSSo��ۨ�x�`���x��+�C{(��'Τ���oBni�2l~����êp`.���?c9�zx��s�fJpV��uݒ|@.�C	r�%��4P��F�fa��
�HenT�xׅ�*�8����t�$tk3V�"�gE����#�Z��������a�:x4~���~�Z:��d�0�Eg�(~����}��&4ʖ��[sjY���K�o�r��F��z�\�l����A����֫
�9SR�^���k��y.�X-HU0[�
RnJ3�����Re&�o#�~��s�Y.,�A��(��B�pl4�+E���X�n�;=��iL�X���V}����jߡ@K9�.�5��4�� w8�l�{��O��h�L�d�q�����InZk���6n��-�%Ϟ�#�h{�bhT�|17s�H���v9�����4��K�p2u�9,�a;�Q��5�;��'�g���CV���`��b�oi��ޜ�0gF鞙v�۰W�Ѹ���G��Le��������Lڞ���WW��W5�U�"�6Zrjk���~ɤ��_���)8ζȈ׽��h-��U��ap�D䏵�[�~^�i�NBN� M9O������[����Ա�O+k4m�`��m-������֓�v��㺆�ԌVb&��tm8å����TX
�:���F�QNLQ�?��� U�5�24���&ܴ9vn��%�G�y�y4��$�����@ѲIDއ�Wz=E�X�+��?c�=�� �t2����V-���m4�T�.4��+�A���u$�X�ZէJvz,dy�P���h�`;�z,�}�*���Q,����Q}d�2�;n��b���P� Ȟ�}�\�=�T�Tf��ݸ´km5��Q�C�$m(79[R$� ����@Y��j��؁c��6J�&;m��Y|^��2�P���=�	��3��$��|W��%TI�#��%�M�O��?�;wz��5�C�n�qg?�)�`������JFe�%'������*P���<��4*��2M��I0�SЬ*�)��Qa�O���H�ElrĠҾ�
��M����j[[�=f�E� �Փ�)$K0+��N�k�_���s�&�ɐ��UBd�/K�l�I+
q+�[������j-�M�+�&�{�3X�u�Gq������;6vW�_���Uz�1�CrNq�x���w��]�����b��ܰS�3�h�.�����+��4�a$H���i~K�(GEd.��F�����d�*�u�g�S~�����Mcnn��
!�`.H��l�0��[�^�9��ڗ�T#wQ�Y�S��)Jn� �a&^NP��gl�@|/Y�c�w�Pѝ��>P"�M���;�sb��cRt����0��6kM�E�9��J��