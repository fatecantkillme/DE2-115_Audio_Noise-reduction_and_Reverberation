��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��/��Q�w���a5P��B�~�/�'̙���S{���^�qѝz��'�hřD~dVr�F�!5�=��[�\�bYzy��d�(5���*������j M����J����Cw&�u����Dg��>_�,��o��3�9=]�sn��5���A<�-��Y�,���AU�G���̻N�	�Ϩ�g�ϵ�w�Ω�k���R�9HO�o�u�(v�W�T�yVL �q^�Q�0/�����)1�cڵ�E
�W�D�t/�Ș���~x��R�X7�]0|��?ͭ�m׭��e��%\rN���H�i��8A(_�P��0];�ű
�0�"��(bJ��OV�[�0h��ɛ�}<pB���oUq%�9�,��Z�SwC����c�J����*X���BH���	U�25���ZcIa��$A���@#�_�*}��n�z�TɋU �6&�S=��a�E��C֦Wr�O�/!M�4��4 u���k:�dėw�X���')}��+�9}U5��=w|-��Ijo�i���s��'�4n�A�>�@D��Җ5&P�	}ҭ>�r�'(�r�F=��/+-�n��H�'[��6���qm;A�d�p�@��@�/�D{>�څ�b �GXϔ-�M�D~�)݊�ks�����~i�6៨��4�2��4�T�?�S�Ԫ��͸�������w�|���3e.��@�W�kx<2��
��A�eFyjP#u�?�����A�����	w�������K���#����V}s;H����vr��5�r~���,2��5k�����r����Bd�����՚�����Ms������U	�˽"��ѐ�C��ď���10����3��JL�V��[.p���h²rG�x	�Wn�����i5?#����y�K1�d !j2���җ�<��GB���s�_\'�ص'�[�;��O�Mݴ�	��ws?�a�k2�=�ۉ��r�=���e�ZJ��\��Ȝak�ȓ#?�b�&ES�t.[c?
i��g�.wи���W{5t֯�ݨ~x,ӄ� 3MnʁWF~��#�XT E�{���L
w�|f�G��GϨ�8.(����+�O�G�jj"iˏ0�\S��o�ug�L��A��+s�GI&��f>D�v>g����.�Z0˫F�ɭ��V�s���R��kfhc���T�F���8�n�����yC�ݭ�!9���XӪ`��MA�O%V��<�	�{��r�43�r���C�f{�&@����&�9B��c�`��vw���ޙ�����Q�6c��M�%���l\ޛICbX	h�n8,,��Q���qC�#Ls��o���W�7�w:�F)h�g�U�����+�F��vϮ�h9r�������g�N�|&-�X��mrt�J��� ��S��͋AX���6�l ƨ�^ZG��Vl���Ps��*_�~p���eˆ)i� ϸ
x�[O6�9���6�P����W���:g��p�/}Υ�ȢA�&@����;-�CV����@�ϔH/[궥r��V��������ϑ�3���3����b�sU*�f��NHG��D~�m�0:�x}�MR	aRb�Ss�DL/�^�aa���_�n]�i�d 0���k��7 N�J��}Ɗ��f8��Bm��6�<Yzh�����
�����Z���- i�7�AS�F��pX@��������S�lA���⎁�LT�f��I	F���P8G�oL󌨫��[��S��H�-�P;�²���XK�W���_"���Z2���.�&���R6B�H�{�(�<��Glc�y{^�"�G0�Hѕ�R׍#� $��2O^؂�s�l-ilB.��/z�� �~�Aq����\v�í���������ԓ�����b��Q&t$K��n����l&R���)�M,*0�O\�q ��쀸��EE%2�u�g�r��ĝ�0qǕ�x�nN20L��\���1+�0u��L�<(Q���ߦ0��{t+�ִ�q^�m��|�R/m�3��ȧzU�v��Ug״�)�_R�Vy�i@t�;���k�(�F�t��v�.]���wut�fZ,������Z����g)'������kB^�I�Ŵ�RX�up��Ȟw��AO��I5s#|׭�f��/y�ya���+��"ߵ�z��9g��C�'�'���8�;���F7E�<=��5� 4�j�}�Տ��-Ɋ��#��kR�0F�p��z���i�Q������<��5d.�q��=�禬[���Z}�8t;��<O�bsz�ضO����/.jz��`)��O�B��Vwd��P��b3��R+i����)�v�B��=��ܲ�mYx�F}ޙ�[R>�>*�7"H�)�
�������Q���G:�ZLRQ_i��@��Sp�(�� �ή*��ȡ�
��5M6�#��Q�r�0�O��0�X[�t��Mz����� �thj�M/��{oy�����syZm���X��Z� �Q��=D��?��E��$(2��w:�Ct�=��GK"�ߒU&���ѐ�qǾ��)4�yc�E��n};Y�(�"�48�he۵���[��z����c�N�k�>�X
ތ�|�6ii��m��s?��ܪb	K3Iо��n�<�kz �wN��!3Y�ۃ��f�ddd��YjT{�BzQ^	\`(%7����^C��)��x>
@�i �a�ֳ�H���w�Dҿ>���,yq,69vvv��7>}���d��iGR��b����弻��@��@��#=ߩw�4ұ�8�\��&���N͵��D�g�����J�[�Y��O�M���!g�`��k޸���G����J,����yx~wr��*-�Zh�>��wd��� @���$ߦ%�4�� ��]'��F}�����H%yJzR�Y�&�H�L����^=��5��fd���]"�5F�6 �}A_5#}��{h狺
�{�`�=�bm�����:g�x��u?�9%[po�I���+�0��\;�S���aV*���C"��`P_�"�,)~��dӹ�{.�!�:��HmYGT�ct�n�����i�Ŝ�Ӫ�3�������p�0����ID�u6k�M4��e�Q
����e������ƻj��������
ۅ�Iܚ�
�4�ġ�$6;����]�d+f���'�A
��IB��6�V�����5|��D%E.��jDҷ�J:��"��2�S��~���A�	�(�t�H�ö�TwH*�t��[�����*Y?\��l��ΝO�)�w�����i��GL�6��-z�i4�z���Q5��౺��JQRD��8�4{�U�Zv�Z8�&�
j����fBC�.����L~��ݮ�K�:�u���9�x�!B���a*�1��֮o�R��=̖--���}G�;ed(�	�FA���߻;P૵g��FU2Q�i�@�k���9�,�{�G �~���WOT$Ԇj�|�J��w�v��w�O��31���Wᡕ �PU��gpw7]˔o;1�m�i��u/�����/i�"�ي�,�Z��s�2i;w��oxp���}:O��=��R���a�5u�����l���}s/��6>@I�����D�BĈ
`���|��A � �#@��M��Jd�
��kM?�=�~/�Wa���~��jV�?.�K�ҸA_�ܽRң8m���Be�����(Cu-Mey��Ƣ�zђU�Dtp���T%;�2����yk��D?�4���Ӌ�R_*����P�Q�

�ϕ���^��S瘀�@��:8>;9;�_��������#�i�H+�V�V�5ٹ|sk�aktA 
�s�c� ����D.'�FȎ=

4t^P�<��������Y�~��2�ҷ#�~���V��P��<ˮ��AYW ��	�,���2!�֦��ET����RqN�[`��H�*
�2o)���nk%����
���է��܄gE���%�X�J4t��(����״i��|�Q~�gO
o�U�~��(��|���T��?d��
7�fJ�Z,,0{ȍ'۞|����]D�sw�3��O,���~�!zua�XH��<�	���w���c��=�ZNDH�h��r��ʊ#�zV���H+<�F��n�u�̀�!;7=�;ŗ�:)�0d���V�Cy��>g����o�y��<W�2JA�o��[��M� �#oƎ��D�ؠ�0/�ѝn��Ԃ�C������mY����٫��������v�����4�n�/)�"8���累��
��T���CJ��`1����w�K�a��M�%�8E�B����ز>����eDٟ����<�<���b���%	�+��H���E7HP��x{',��x���
���pM�Y~��S���8R��D�T�bm
JD��Vb[D>�����y�L,���2T���.�78'Y><���ƇF�<"_��DB��{� [Z߻��|�V5��n��������u�&P'D}&kZ�@~�@���M��`�›H戮<`gf̜��|x�?�p�	�����o3L,��(�<�j�w&�2�4^Z�Y0�C�H)кB'��αyS�bfkǪf|��E�^���"�=���;�
Q��sDt�n��*�	3�9"���HT�S
\nS'��a��'�K_g�o�k5CR�����J�Hy�t�wZ4��C.tr�"5H��I0�m��5����gLg�Ў����=h���c���7�K��R��Z���-��o�L���-ʘ[A��3f���t���3�B.V�r�h����b��JmET��W�w�g%�����:|,����n��84�L� �U��Q6@�:OL���p��s�b�^�w?�݉�')������c�����L$&��ug��4s0��hM���tӎ�b�W\얿j�]Kfk��c@J�����qQƾ����Z�)�;6�֚�u���Y4�'����bz�,?�l���ѐg���e��:�
0�=�w��2�-��'��ޫ��/+:H�@�������ew�Q��7����"�ZuxYfC��]�����}��l�+5�������d�20�4�>�PZ�?M�[͈)5#t+3Fw� Nx��M7�.Z�;�w�JP} h;��+i��3�������J4-�R]��N^�5Mr��/�hzx��VB��#���e[���#��ᦼ��}}��Iv�������髹���G��thT�UQWvN�+���J�R0I�ǌ�r_@
�Y�/��^�ې�}���I��#4o_7�e W���ş�V��_�f��%�3���*GY�_�7��E��o��$4��
�� �Z8�RU�|��+�*h���O��#"BEb*��q��Þ3���A2����#%��V�2�C6�����N��e�t�͇��n�֨6޾��TU��ʐ�R�4�䑪�b�_A�Z�M{���U��<=Њ���(bS$�5-���*XP��:�j�����2\�[����A��m<1�:.���>hzK�Z�kz��Z�P��&Jmr�eHT�D͛��zmv�����`o�O&J�)Vc��֔��P������c�A��PD�0)l��)��F��2���s�]e۪�a��_��#i����Q'�6h���#���ض���YzU�������X���l #���s�7P��Μ��r�f����ho�7����[W��A�:b�ǀCp$�(��W7W�I
��C�ݒ��H9/j/"F ~����MTr�G�`�ޖ�]��}�UV��#^����8~��d�l6����t�
U����)���S�2�s\�f'բ`M9�����	��B�;MM2�tݽ��fcn��	}���~ uT��.�^+��w�v:Sy�3\����K����q�d���ۢjDC�!::z�#E�2�MF9Q�vs�Qq��l@��b&��#u�w3�e1`'��?�(^Cͬ�����4�nS�YZ7�UZР�n�'=(�X�޽��Rn2gţ��k�$�U�g���:�`�*i �x�V_���I�aӋ�D�����#����;ҵ��D
T�5�k*�４���/7î~d(�Ц�����#j<�D�띈E#�5|�����AG�eN�b��Hp�v�6V��n	h�
��v"���y���#N\B��� �H_K�I!�K�o|�_oKxd�����ڟ�R)i�O)m��� �%$ݫ}^v�&G\yE��e�ӆǗ�D�:��FW�yw���xt:�?2w�?�z�8������|Q���_%	��9�����[R�`>	c~L(e�	�|I�iJ�}� (@O�6|$;����,�����lO��8��^Co�`�c��j��p�ǋ��K�à-�R)�����]5N��a�/L�*T���g��s��@ %�2��:��Y�T/���O����A~����i���
����YvÊ��U}4 d��[�����*D���	^3��i��q<B��|ě��0�T^��MC��X�[�т�PO
�hc������}�,յ?w���`�X����o)�O��皉c"�P�t���u�'5�]8/�bڨӰK�f�ҵ�;<sG�&�q#��q㋷��?�
�g*~��L�dK$O

\�p�����D0p�
�}Cn��i�{��5ĥjΉ=m�M��|�I�X���8j1��۞�({��/�}�W:D���Qͧ2�9��%Q`q�V�t�n���hh~�_�z�'���M��B��u0�&��ei��rã�v�WR�+���rk%~š�� M��/7�χ�����j�����M�A'�	xcI��DCW3��0���7�4�*Q�H�����E.�9��{5�N=�@C�d��w��h�N�Y!N������;,�₦����a[��t,�J���lOX��2����N֌���X��eqʬ���ol�r�e��X�և.�TN�Y
w�\!�� �V?MY���~R2>��V�r�����0v`�c�E�r6�R�����2y�ʅ���E�v����}����|������t� '�V��/���#�oD\�eJy�B��c��NN���ښ���U{W;�(%�!~5 �D����uON='���2,�����0����]��<(#�0O�nMYvê� �j�Z�j��5b#LC���Pd=�_lq+�o�m�u�	�`��g��c��1"�2\��V�e ������-�9��6��e>�*xh ]�.mU�EW;�5X�h�=}��_�u�(�I�(�x��b�9�V�4F�1�+Gm�ˈ�8�� ����.�p(���]�f̰x(0 \#R�8WP�Д_K,4ӑuT���L爦=Ļ�]%?�<�W2���P��L�z
�9�{$��5�#8�A0[*gĬ@C,�e�}��=*��-.���C�}!:�Hh���g���y�`6�%t���b�k� ~=�L����n{�6I\�xص�ء���mkAJ�y��zf���ўN(��Z�#C���W��� �2��s��,��V�s=������A�|F���	���e;�rU�5�3�R��Ĝ��[�KΗЉ������1X�t�`s�� ��#�qGVK�� '��7�o�ӡ���9綃��N��I*������k��nm��N�qV?�� �I֙�N�c
�ԏs�}ve��K��xH���a?	�P�Z�	�{���=!��w���{,�,0���im�Z8���b�?�&#$��<�8���{�xE�%H��5�`��p�V�"���0^�]˂�c�h�V�����U�y<�Bg<e�����q�{���I ޵-������4)Sk�7�:�Kk���rճ\�E#� �U�b'Nh��HG3?Ţ�"�
~C���:5�O�G�fؗ\��RN{��V��zg��9����͠������s�a�쥉�w��}i?��Ccx�_�Ӡ�sql^n�5��/������?��'���(�u�혱�{2��̐��2=�b��D��)#��;��m8�So�,��|��M