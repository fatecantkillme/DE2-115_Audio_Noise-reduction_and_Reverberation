��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<�w��Bk��J��3�Z5��� %>\	�H�� �`�z�.?'��l�<'�U(ן��Y��d��ւ�)���p�C��K���2y�Dt�Yo�&��V�7Z�:��^io�,��0\o��\�Tj�g�M����|��<�X�E�#���u4h��$��8��3�I�����hS$Z�̭9*�t(�-f�_�*8�M����F?��[�v8m�}���cEn� �>�O�б������~�Z��ޫ��ÉɈi�,�2�7��T$�d��.Mf��]0����┙Ȕ �:������N�A��1ċ�+F�K�Bf��h��n�hC1��2�_Gً�R^dz頂�70�����eqP� %�d��p���',��5��hK���(�z��g�.#�4��B_N`�.��X�\ � S��#�̡1.P��]�"կ��ɟs?E���m�u��}�(���]�"������ز-hЉu�������'v�Vn�����GZ&�/���e c�������n���=�|ΏuI��iO
��Z��A\�1�\;�.��~y��k�fç���w��'����UҨ���_A��a4p�Ne`���2M_2�+&^rݙ�P3��xlȠ^u�-G�ѳ��:��#¿{5�19�g�<m�5K~Gp�-!X�ϰ�W��{��	���j����+G_$�>}�!&����m*�?�rpE�?�9կ��P���cq��%C�C�����֤g[����ٱ�mI�F��#<&З�q���W�j�{�jrԄ1����ьs�P��Y��{�d]���am��"��@T-t�}���w�W7��<�s�?۶�}<�`:��
��`�R�����^� �wF����w����A�-�g�����-�,d��xͩ8w�⦟c5q
�
b"��^�EY�Y�=�P�$T����� q�D=r��mj���m����J��,���`�s���D3������HS/���dO勏/T�Z��	��c�����ik]��aq��%S�o�^�lSr�����*:�C��q���:H��K6�r}��ʝ},�G�z�����V�"f��a<Oe�����F�c~�Ų����oMXt���l��O�֭�W���s'�F��J#N�U�a؇E�o�%�ħ��k9�3����y@��W�����O(�����������$Z���26B�Ƈ=	c���3��?l��n�+�����u����P�ח3m�)��o;�~���^�4X�oѫl��l� �󳭩%i�����ܞ7�/j�W%۞����W.}�m�x�{h+f����&�֑v�*Nj�>x�^��ab�N��^T@��e��6���\�V^�����>��N��M���c�X��˥pEB�'~Փ����^��څE-�SUC"�*�v��������ipH�K{�:��.>#KyJ�����m�f�@Ҕ@.aDeq����A!"ݍ�%>_\ 7c��Ǣ"}QH�S��`��P�g�X �NH��4S�R�Γ�/3-1�Y��nγ�%����5��>]��OohG��QI�8��1Z���uU2�K�F�lwl,�|C�X�F+��G/mR�B#T�ڨXo�C��S[`VQ?�P������6���8�ʕ-��ˠb!C��͖�L���w�������
��yW�79&�3�;��J��Բ�v���@8��w��h�mP6܆���q	����챚]ϦGw��U"�7��rOwF/���@�">���F&J��~cSN�B�-�w��4�sx^�D��	��4�З-�x��·q�Yj�砜�r���4��M���	�?�*KQN��ј�����]_ _��J�#�$�/�3�ҒЛ�5E��o阶����R�=�,Sy�T��֍�TpՍ�y��O��+�&���I"��-l(�>:J{퍬��i[n�B�gР��q�j���M���hG08�>�Mh�g���h{-�Ņ�=�-+�L�䔱gi��7���$/ɉ���P��ӈ5-�8�[1v4��`!!|�!�������z������M-Mb�Ux���Z*/�e�ñ�ͨ��2��ӳ�191��O$���
�̩��c���x��nA��d��)'��c��q�9àY��ЕFx��`�ȳQ,D�Q�Z�Cw?n�V�;�,������b�B��3:}�l��5��e��1N�كG3i`�{�8%������ݠYݵ�?Fp�Yk���J?HE[p��N�����_n&�w�2Uz� X_u��w�����e�^/���|aSkG�����c�L��z��p�M@��� "��8o`Z
�&$ӠQì�B2/���>"��p��©^~��6�k�xS��jl02nX�~�O�`�'�U:��=�E�4�H�ɏ'�����I��.�i��'����:�xC��0���!��>�f���J���zt��&�ޞ[}�+��1Z`��������4�[��Tt*�T�y��v҆D��"f�,�c%!Xo��� �v.�4���������HzϤ*QI���Q`i����Z4�>����Q��ܞ�0��<S�^6{`W��N���sa�B�v��e7�v������^T�v{Mc��C�>נ�H���?���hYƦy�%�#���
ly�z����\�;��0	�и��8f�zA��j�nݜ\�쨊?>*��Պ�xU�G!ؗ�W�5�r��%U3l���҈T�����׍�WP�*�x��5g�𺣢��j���_���R��;��>�s��o8���`��
���h�MqʹR,�&�#�*<��(ĺ=W��ګ��?�*nWA�����}���P!�=>��T���=�>#��zع��(t��|���o�����e�a�'|�F����2�F�eZ{,����މ=}��#`��gp����������)L�^w_��h��[{��'��ԏļ���ӳ������,�`����2��Ah����k'>d�㼗y�����*���.�#<��`�W�{� �8	���T*֘V}�g ek�H�"���(���.�w-;���':�m��O�G�*m��"�N�K_��_s�;��x��8���$3����W�[�4�d3���v���'/�33v����Yױ�#�z�D�v,�4��@�V�)봦U�?�4=_ʲ�1j��@��oSԎsY�j��'����C� �5�2�b�R��ᦏ)�n,L�� =��RN������f�`(Rl���w�
]��/�<�T�Ϙ�=	���uֿC������3����u�i�y�+���̂�c�<�|��l���~r�8��`����͞���FUL��+D�8+��8� ��� TIkD2�uj�5������I��@����W���hn�voռF��>ϦLW���K�pG�0���	V��'�i]�,�Vg���XD�i��ba�:~.a(��6��Y�UJ�a�����C�Վ %�g�q ]_`u�� ���/�� ��_��F�5�+e��@���8X�!���B'����3�Fa����� ^�=^�K�zHf���*��d���o6��Һq�� q��l �K�k�-@"����ֲ�=`Q�C1���>&Kt����*Y���
@�-���lde�Z�[�{�c��\�n�iKk�n�P �
|����3�L�����.w��j�i7��{xI�kg5�Bn/gq���gP.F~���.�����P��3-~��oP6W8o��gU��y2���v�*Y7i��^![G�!�+��m�]\x���~�Yq.�!+�+e��C�@c:ȡ12~��,~!ǽ��� q��?-H�y�K ��+EE�-DJ�����jFZfz���x�Gw�]U��"��yŢ�u����_��g!�"�����9
 W��.��8-�
 ����ԚN:���h�n�#ހ�3-��~��-�f
�=�5�d���|��nos���f�"�!I2��l��g.�`�FEf��3S���2�82�:*j� �����#��pQ$�鄕��iF��w=���D��Q��qr&�L�Z$(��#g�U�W��	�����A��+g��< �%B����8?d�|6*���,A�n�CO|rAp�������Y�j�ֆ�]�)o��9�,:�Z�\,���c�ϛ��3,N����հj43f��]�c:=8q����g��c�:���
�&��WyC݈T��<(j�ń��n6��*͓�[7�Y�4<��mz�����/�˰�5�^|O��vb3�UՓ���y�����5B��F$S����aDςv*�R�v��j/��=�)X���C{@w��n����Ôle���_ɀN�
GUY+��3M��od���d��~�R�͢2[:����W��Dǎ�����1d6�&f1}�����yt[1��ⶰ�yvP���h�ȡ��55�k�!��g۾���Ӵ�$���n����[rWt��!xk�e��%$ӄ-h	>Wp�P�%�� m�D�e�Q�ŧD<�%SmTmS��s��4�Y�}��8-�����}ɧ+�C����\ݼ��>+����-r�c�w�-9E\��G;��3��z#���Ž�3H�졀U�۹,'BIe��f�ޏx�=3cw�J�)�e�WXA_�;����gd�!u�W�<���CޖO��%�Y<���N�V<�������s2�I���P���o�0�@��!U�%�0 ��8���):�%�y$3')��ܽ4i�3��8m }�F:������V��U���}d�p�!�֣wj�w�'Zq"�/�)u>���6/8\;�V���4|6iJ��*��?Og��)�0�
G�~�U�mW*]��+ 1���	ՆcX�X������K�!��I�=d�ar��ecS�ql쉓\��H����3���/�c"%��^-%���R�[|���|Q��;��Ǻ�Җ��r�k$�'���?�V��?c(]@x���Z�:���#�Dh:P5YY���g���߀O�|��17�c��[�ew��󯯩�02�\�z��	��
H��#H[!k5�^U�,��%�ځn���Q�Ć����`���X7G�d�r�J������^�tM1n��ۣ�)V�#�x��g�=:�$m�9 #��\@\��+ҋ�r*Ǐa(ǌ��,����0����SN��X_*�-���p�ͲT ;��O�'��rr2�UPɫ2-�$������<�X�b�\t7�M9*�`��{"bI�©����Io���ЯC��|�ff��Yn-�¢H�{4���W��� I]+�hUsD8a��Hkݐ*B<V��,�j���uc5F� .J��Q�a����)�����	g�穣CP����ݗ�����<7�7�s%�ħTܯ���7P͸sX��D�u�X~�%�N~���P��~_�ėk�;jEv�ۮ��g���jS^��ϲ
��Mܾn��V����n�� i�;]��A��2���>�"��h����зv�����G�!�K:\s���]n�S��ˊqjFX�:ϭԷ���� �&�U�����)��D��z�ot�;�:�O��u;�V*��]��wI�w�:�F�@\=V݅����2�+ .��z�:�^����L��Ґ>��;�s��ȑ�k�U�a��R�4׫6�]�|9/���P9n$��3U� �}��f@8�dO	��
 ��%�S` ���0K�=��u8�������j���<^��!��k�^���>�C��H`�Z�׫�שw�gZ�~B+� �m�a����{�6�Q�����8n�8D��K���rWI.��ǆUwqǮk�d�@PQvd���~-/�p�������8Kʐ�	B3$�J�{1ɺ�+5��H��**y~��7��/���X��i�)k\�,
F�n�׀'�z^m/����,-x�S�r��\u��?f�R�1��S2x����UL y���iz7�'����ؓ%X�c���h?&R��l ����L�H/��6�g�M�c�>�1U��Yhs���NL�e?�� ��o|���m��$�������F�����9��L\pv�蔇\���H8D`��G��6��q M��>�'��Ԑ��}��v�8�v���<��x�%�=�VW_/�Ml����nseً���܎��\R��/�.#ۍ܀�J?q?%�����޿�LMB���i����0�5���9��`l6K�;˴�^�"�B#�uU<. Z���*\Ǒ�٫��ޝg�Y�c��	���a��e�9���>�=���Kj���A�	��6Udx����F����4	�n�9W,Z3ku��\{�����M�·%bc�Ci2g��,Ǔ45��@��G�L�%�y<�=@�[�%�������h�	�D5�7��R�(ߝ!�����ŋ�~U!�O$����gy�u\����9I�Ԧќ�W�H�������rf�%�f	���`��@d|0��H_>�ƶ�B�?��I`Ϯi�eR� ���s���>�fp�/ 3 ��q� ��$]�b`M_#%'qY��t!'�fy������[�j&F׆��R��@5�Q��a�x��хl�_�-ر��؟"��+���v ZH��ɞd'wH�=�uTV���J�����-v��(����E�_y>/8�֎i������R{u���R IZbE�=��K��'������D��ت��1��q3���T�w,�	������g��GA��Q8ڌ̙g�A�_-��/�ʘ�Z��ޘ��7qp�di'�}�C)�~����������x�RY�V��� �����IG��YK�a����K� %��}�
U7z@�p��qy��
.pv�i ����.4p9P謩e�:k/��y׻݉�����<���<NB`ӟc�fZ2��(���������ͬq�,Px-��{�T{��r�+ڽR;��y	���\��H��,yl���WRgaoFs�4i�y�e��QH��y�K�B�|D��SX�"���pK��=t��._�fX����[��v�в��7.�!���ŭ2��J�x_i
Y�肄�55�vO��=�Q���S9|Ù��bY��a��gf�>Ù>b��L�oGثAM�M��{L�Z�gܺ���Q>��<���\��i;��6	37}q�+����=��]U���W��c�s�A���ճ�����)z!Z������R�����H��X��h��������{�Y!��� Fu���0T��*��_�i��c����0�#�H[�S:����G������xU�B�h�*�%���V�!/�\��%&�l��cѬ�w4�l>�0�Ӿ�a�(k΍e���V=h�f/����C`��^��It��o�В)��sE��1��Z���\�΁�k?���'�׎�d�X�@t�b�",��Ls�W=�|~�I(ʈ�ͮ"�;��b�\�)�iL�FT��d
��a�A�i����^�L�Ɣ��@��ҳ�?��U1�+-��<#N�%������4]��Žgn�;+��rG_��N����z2�b�I���%�
iaS�ƫ�\f�O$����f���D���k��
Oxv2nb�9ʟ�Q�����r]o�͞�5�l/14Q� ���O~ �7���i��3��S��׮[*����T�tW�E��?��7�pZ�5���p��&�4��ՠW�~��l�^<6m��RP[���}O{��|2��wv65���O^�}��24��h�Q.�n�7j8�ۯh�"�.GA�~���-�668�.��Z�Ա[c��:����YVk
h>eZyM�{�08�"��y�����O����Ns|�6�=?��v��W��I�kD\z�e�#3�W�o�H�C$0���-4Y���X��n���ʾI�㪝��V���k�I-�º�e�Y�]M�G�d�T�<�?i~8� �i��7|/�dX;����n ,Z�Ω�"_�Ch�r�&a�"�R$PN
��T�C~a��ߪ��*� S�r�9����jR� d#ĩ�h�����K�1�萚��s<��A�6��2I�%��}Wt�8����%�[q�B*�]_����A�ڐ��k~�%��ef��'�12�c�	f�P�@m#���R�ci�aI|�|N�YVۤA��͝��x�up�[����>�rY2\��h���3���Hf�'[��Θ���9H!M�0��D�d �!r/PIZ���|h��U���Z,� w����' �_��=�1S� �n�t�4_���:k�+��᫲����8�?��!�ě�T8<��k��Wu=�w�7;���*��~-"m��5���p&g�bq�1K�0	���Rn�-���p/:� ���O*��Aݷ�J�H�&�ArMp�ϩ���"w�F�Bk|�7v
�)O�q?�ēђ�!� :�4q29ڑ��v�?�w�b��1����fT�q⵳\ӝb���t$!�6u��Y`.��Ou��3��=�X۾��?}�"P����� ��#�<tx;�@Z���\�.X�O7�0p�ic����X�MX�
вG�7���H�^e!�g2�hׂ��A���uWd[��D5v��3�D�������i���'r��#�8D���.?;�`���$eB�D�
`�R�V�R����泻�$��*Y��W�f�g!�.$���_w�\��te6�g�~a��@���:ӿ���-��<�I���i�uCvm��A�I����~�d	����b�E�m!�Q�c�����E5�ZC�.`z����SVnH��ݳl\m���j��3P��p���2�x3"�M��q���ЖzDY��D(�y��s�֯.�rØ�~Ⱥ�:�δV���kD��ݳ�@���%�����\��Bmq\�c�N��n5�j�xp�	���j����ЬΓ��V��R�_(���ӝA"�M�{���T�皱m�o!,��9W���@�'@��7w����I�e�`�T`M�U鱛� ͽ��ݤ�D�#컺�9����eEE��wUTP:uǻ`�<��J�57�~�bjɅ��xCǉ����lI ��P�H'c��8���n�v�9|`�b.��j�3o����H��e]A�ta��j|���BJY�\S��}�X��8��*��@��z��վ��Ƹ|DQ��\q��-�(9.��>k[���(��7Ԑ������3���+)��~Wȷ���f�Hx���;��^�+oϺ�o�q�o?RB�o�rp�S7��%VW�nR�\[�cVDv�8�p[_O��M	 d��+�,3�B'���a�ş����$Q�"��n$�	�ye�3R�m�+5��/�g��x�r�Rj�"��l����f�n0|XE-�Km����a�<%l��{Ҹ�[�t+�m��h|�ј~��Wp���`G�FG��~H?5�����s�#��;���x�l/��1˟��=⣲?�+�Y|�d�/��[>�*�LOqB`p�w��Y�����c�M9$�>ܫ�K�Gݞ:��1�d��N��f;Zc��:'Gʋ%1K	�\
?d+����^3l�����/����[�-J�͈��p��ֿ<��rR�Dkd���� �jT������úz�ʕ��<G�8<"��Y���h��x�����[�<VP�F��y�<x�I��e�������Ҫ��,���2ņ�jM�vHm������ 4����	3Ҳqh����*4��@������AD0�NP��A5�+1���ĳ����*0��EB�v[Ֆ�H�i?�#z�=R��ab)�Ί�Q�-�2m��YpL#�(+�[J��q����Kn��N���Ȁ���������fЌ`4f�ͩ!k�����kE����o=z ���?(��/�e��k���à#,;��/tCBy��͈�E�Ix��N��Fޙ���!�f��+Z����s��9=���c�g�c��q:I+dC+Np�G��-�Q���0ο<_����۰@�H ��d�}11�h+w��P��b�+@�i���R�̰gp��[���|��WV@GD�/n�����͢g��њ�F���rT�}Ya!n�V��Fiҋ�g��]�,	'>��o�