��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<i 0*j�_噰i�E֠X%9��
�Lj��4�?��!π�0�g��W!�J��损�Qn��������!��c���!�=�>8܁�� S՘(�Kw�Є���W�ڃ�1ﱕO�޸�xb��.g�~w!t��h�9jȇ~�i*��D���2i��p�x���BX��q?��ꞩ��}˕�og��J\�m�9���k7��6���Co�3<�`{NӔ��)�Y�a�;��	��e��7�4=+ʲ#b ͪCm�}�l2�~�&1�tN�s�%�FΑ��[a�Ͷ�{|a�A']��^g�$����`� 8�}��ym��,!Ek�vv��X_���t"c����8J����vs��bCW37�<u�b̀\}�_�;$t���[� �4�K����$p���a+��"�:�T�������[�eR)|4���hׂ��(.�M�^��PW��ͱGZ%i����o�ȸL}����o��_`-�m�K~�A���2{{�a��'�I�[Q�������;L��"NR}�7�}��Є�(a�[�I��s�Ҩ�mM�L��-W��Q��������׊� bIYU��	��APȓ|5�G*��`�t!$�'l��jMj0�P�-+<��R�;p���s��?qҟr�'W�.�WőM?N�j<�*K��hv-�Y�?��Q��1I>�»:�����U�N��Gy7��mQ�ɉ����E��Qܣ�|�Y,���U�.��UG��f�by�������#Z��2Y�l���mС�}�gy��DU#�(Q�+��.����zц1 X�P�A�2��s��@${(qȒ��wh����� �@ٷ 嘵���;Q�=[Ѯ��W!����?4��W�ûv�=p�#)F}��16�n���`��;Ұ��̔�7c7D��7B�w|î:�vU-�m�ା��J�n�U�^�5���`��Wr����c��;��8� ,��d��V*�oAAM~���4��Y�+m@5eAO��V��'ņ?0H�D�j��y��ƹ��(W|�4�'OQIP����.^��֪_=lK������Y����;�%������S��m���V���$'׸�R}GY�}]Hr�Er��)�^u؁4uc����(��]�Ώ[��,��+u�jC��\���
��2F���*�cF>�-K�2��N�/, '�$u�Sb'�0gx�� o��\ \�D�K:̷G�x�x���.���4_�ew�&&dR������~|_;?$�Ցq�kQM�^�k�/��ݨ�:[3\��l�z���>G`�C�����0�~�u�d���&%��~�՜5�[���x�&+d�T�yEI����]4j���_�fFΟ��w���W��p4))�-,8�OEP���U���C�u��vA�6*��
V�	ο�~�f����Rx}�I7g�����.|�ҋ}3ӂp0���6�_aji}���v�ò�1+3b�K���Y8,{{��[:.�2�[�o�C�ښT��]�h�w8n��?�n��XiTK9)�����;�� ELd�w���P�_H@��ً���-\l�S�&οk���Aa5ɑ��pJ�Q4�G�9�5�h|��fʸ
�E�O�)���pg����h�T��u� X)�wfb`�{Uix����	2�J�>�B�۵m��t�ve-�'�c!�U	�]�[���ä�����ш���N�ٟ
��K�,�g�(��	]3�L����K߿�-�����%�A����W��K0�l��l~����y�F�A�<�2y����k��@/[��P��:��F��m�`��WD��7�����z����i�h������Y��ǀU��O��h�Ҭ)�L<*b�x���G4�!@����wB�xݣ�s�f�KLd�����N���DZ�.��c|$�}-#��!�l�Y+��SQ�w�l��=	1Ik�M(�-k��i�V̝/����O;�q�46��k���u�OH�xL���*ޥ�a��a<6"S/1�$�֧gn �M�v߹͜�F�ŋ�_D�21-����B ���ϥ��\�1�X�5���G˨�о��̬}ZR GDc�`%c���̏���.��8�>Ij�cu9�l�e�1xj�b�?�?b�p!��TgwL-�y���V�f�p^g�r8�p�!H�L��=ܟ��{���/��j~K��#:���v�zz���yL�ݦ��_s��V��W �M��X!-��.��&�	8����]T	�1�E�	�Y5\�v��+r���	<w��]���So�F���}l���{{�4�M,�6Y��$��!����H
E��S���~,�& 0kl��l*8jLZ-Y�I�;|IS�$�h���ïU;~�m�+)+d_cE�����1����&} ���!���f��t�"��f�#��҇���%�{�b��*
R��n=�(`�m_�BVdoJ�79[x�UЎvg�J��E�Ze�}ɱ��O�R/�|�̓�[���u�85[�ϐ�Eٿ#�[�� D�>@�UQ�ؑ݇�������� ���/?�͈�0��\Z�<Y�я@"���J�M��^g������՜C��8�0(�q߂��
�y�s��S��V�'�q����E܉�R�>vmXܼ��fvf*�59����%�ECn�S�R�׈�s�~k�4S���@�i�d�
˟l՜��Z�A���ˏ��?ͦ-�&(
	��w�|:Ur�r���Y+�RGiv+��Y|�J����8h�p���".�6َ���H=��$�/9g&��[Om�Q0f����$k#X؃3d|�4����щ�$�S���жN��C긾ÄI���:M�r��t;��J��OCy�~�+S�����#��9e�w?3e��u2X�M�@�ܕ���+�<���&��=He�pEW�݀�5ۈ��p��RR����o�� }2u��M�.6�bad�y�u��Y���(E`U�H��+7�S���1+e�m�%�?��'�t����P:���J ��c6�kF��"F����g\�EX�ZS�*��j���>Z'��ӭ��C�/Ւ_40�я`	��S��Ιq�z�'�/a�e��hxE/�Rg��%�=xJ9-���5$~<�^5��Rә���PF�� @f�)��Lj��K�Ƿ�(^\@�G��L��y͜�@����N��MC���cn�˂�����TwZr�8&�@�  �LK��L�g��q��}��@־�N��m�o
�ڬX�1�T ?�A�U/�E��L6�4��p�S���\8�|>�0����X�p�Z�:\�9Ao�{�z�O׾�NCI^�V�~u��ͽ�d���h��z>uL�P��~���IDӢLj"^�s�F���z���{q��d�F�_P$���Ss'H��P�4���Sr���/`|%�m��s���^������5S��we�o�	�+�X�KZɹ$�$2�$��~���,ctJƤPğ�FR};�z������(�A}�&���7�9�
s�a�+����]*z��vO�
ܜ��ͷF�h����,���cw����m��4�s ����uE�oVJ;��j���d�I��{����d����D�?]A	u�_�'@�t��o5��$ڻ��Ǭ���4QJ" ��<��9f�M����Ӟ��o[<�W�ĸe����������H���8��q��~ƟU/B��Њ���NfdE�h.��uC�����R�z$C	�}�C�tw�z��@���^ �G�#�9������:^N5ھz�^)��,��
Xt�T(�`.P�sj!t�����7��*\�.N�I�BME��yy�E/����;�>��.�1Ĕ��B�\�1e�0w��F�����#�6���w_���E���9��-e� Nq�ˌhhj��&��i��+"t��)=�ؗ�ܰ��	����r N��|����s�*PW ��Ո�|�����e#z����;�4�k�u����>�"mj���A�-�h΁,Ⱦ]�%���#�`���2��gA�*&֚�_�����SZ���\�ސJ��	�f�����Ѧ����+ȏ<��*<���XV���SJ�� �)��5�|v������+
օr:+-��e����[��5Z�[�om�
4|�p�n����`0���d�����p��%��f�� H�![�G,��h���� �sn����yLo�^���L�n�z������9�`c�Zy'���j���/Rʈ��A~gR|��m>���9��^�Z5��p���J�[�-�)cq�������<����K'�Z�Q�����viK��Z�TTқ^p���x���&��/��i�`�wg��Ӈ����3�/�gLtQ���:���NC�P,�Dc��a�W�q��;E$d!?}T���َu��ɴ왰?���v�l^�4�������= ͊7N�G�X}-�+t,Gf�BZ~����ٳ|���;�0R��#o$�tlnYρ9q�϶m2�Jɹ���Βuҫ����Rl2w�s�������/��W�~)�QMye���eBi�,w��4`�NDn�ow�go���'���^�#FI�P�H�H�s�X<&7��������݃��T�"��48Oqì7��C5w!S�kt,0Ɔ����H͢z�yP>�b(��,W�]-�H�|Ъ����E����jf�`�hK�	?���eDW��*"���ʉxZ������q���fd�2�[���T_�BMAՅ�����2K�G�C��P;��U�A#)xu�\�F+�����Z��0���EY�_x=��>��I���>��|-X}���h"����{�4��fr��sWK� ��g��NI��Ĝ�R"�HÁ�Uɑm�<r����Z��c�^T2�q�OPSV����#��2Fv�m��в�6Dځ�e�v�I�]�޸P�t��
���T�v8[�@�U���d�ПU�~t�L�'�;����A��&r���>-���������\����E�����WK�&D��u�Гp�
1�';D��L�@��֨!9�ƒR��3�m%[*T�Ȩ�c�<�R���X���'��D�e������� 
eT@Q!aS��(xa��F�"�10Pk"�������P�����L�SU���x���'��v���.d��g�Wk�w�Ӹ#7�a���4%f:W?�1�?K{���ܵ��淴��$��{����=����:RL!M���J4{��W��ْ~��]�T��l,�I�E�b��D�k��}����cC�b��ױ6��������g<E.պ+�jG�6����<-�`���dc"�5=û}禛�kqV�����N�-�X�!��5�p윳�'�XM"�8[?�q|��"t�𧈡�t�}�n��*�dZ�)='�+��:'�m�:w<�,�)ސ��	�q��A�)iY�r){üѺ�A�>��j�U�L#��6jQ�,K�=ӭ��f>��!V?a��F�,A�$�f�a�B<��y�����k��#y��k��Cl$+�􋓶�tfD��wMv#_ 8Ј�
C�p���:V��Ø
�9��t���j@0�h��=��>�e	QrCñ�����K8�eQy��\ZG"k��X����&��4�^�Z�#����<�ys��v��<�^)�%�����8W�I���Y�C$��^z�2,�w�P7���XI:�X��:tu�БBƥ6�e+.B���X�"�џA�I�P_���Px��4v����b%��\e���~!������@�yC���d�B��\����$�r��'�ŀ�L�^���AA���K��܌Ŵd6)l���@��Cv��%�=z֘�w�FЬ��	��b�!,t�u�W�A�׀"���
79jt	T���X+W��f̘:P�ľۂ���m6b�� ��2��wl�$t�s?��l�:����-[�  �UD�_��;�K6<����Ih� X���s�b!�;ϙ��:��f� `�\_)���)��rԨ	k�=�NDrRL�͑W�h6Zb]B�s�ۓh��|_A�X�p<�5����d���[q���`�@�5��>4�ׁ�:���_>�T�Ʋ�+W�����x;N�X��H�r*L�G�(oe��1�S�1n��ͫ�r~�sY=���Z���5o[qŏ@'xZ{���=R׬�Ht�ʌ�X��A8�G[,�����U�7E�ia�{��)nMkh��*�`J�Q�,�j��7�)���b;�����K�D^+��XVb.���%G}9�5�?V��|�;7+�Y�0:��*yl�ClU� �,�1�$7�{	6_lL��%�޷
��w���p����،"Nvs�؈�X� *�g!5�[Y(9���\c:)R�v�Jv���d���a!��JC��d��*Ѣ	p����Nע��[�=�8@;/�٫11��n�>��4�bD^@MU �7��{�T�km+��yImW�Vz�T��b�����v��q�Ag�&4߸�R�T:�
#:����L�;����+�Vc�BU	�Kb�F9�ό?G��_��)v��Ny�ȻWH�7�7T�l_<))D�7~����HGa��iF��/�]Rd1~�d
V�@��X����}5�8�Q �{R�#�����n�xW�3�
R �='Q�B$j5t����QP���
��2��pCR�D�* f�{�O�z�6�x�X�����ԍ�S�W����I�K33JE��#PO]A�|Z+Ӑa����NZ�/�x�1�������2[���gR7��2�h4�����S��^����A��t�kf�}��N�i�n��g�|�P���#�dtkR�ߧz���Q��C��$�-&�+�\��U�P�6	o�W>=�Z��ba������!�����v�<[�lX��r��T�� X*Wd���@�Q�X�J��t��7*ꮺ��� ;�����xp(�����lC�P��,�ٿ�k�[��� &�3 �໵��L������iMyA�����k��7�޶�(8	r���N��H��~���x�Կ����/�F�D��m��zHB�<�Gٴ�"�#�ܞ�ƛP��A���$�e�*�@��RMXz�I�qd�����FpcF��a&fI���o��h:,AR�(�z���#>-s5�;}��.��(J临���%���s՘�Ի�
�����B��wY��u -VN+A��q�1 ��k�\hF��~H�<�������i�-���x��$z��m�`��v�$�gd��	��L`�?��Jz�ӡ���8V �Q�s��z��� �8,C�X�ЍirQ�������<��+K[#"�*]S�@��fB��k�mrB2B2V�U��ݞv� ����*�B�JMH��q�E�����3��a���{`#n�f�[Ԟ4I@��嶸w�/E�>X��ރ�����y�x�\1[߷�Idߴ���enB���X�,�j2�x�֎���+��O]\-��������B�q�NS�E�f�ϱ������_�R�FqjJ5z�O(�M�')w""`�N{�ɎP~�&����h{���y�R(���sJ��/�p����a�n�jĚ
 �s�뷼@Z�2��
S.\y3V�%u ���~��؟n���t
o��U�٦h��d=�%�7#V�?ں쬃��`�E��3�L��7�	�;�t�a���笄y��j�q�s�e<����� 9o�=zƼ�5��Ҩ��OB���\�CQwT���pt�m �����l�vV�*Eh;Jtj�äZ"�?ù����N��u�;f�'ON��s>�'���'��9e�u@���Μ�E @G��뱓�\N{�!ԁ{n��aJ�ۊ[H��X^�s<�{��5�v���/ߦ?�Vz��3��o�ʹ�3K��Ĺz/�F��Z(����p��ϔI�W5\F\�pXV��Tw���<q������b�5Hȃ�9ҵ.g.�tpٌk���`�s@�R���j��P>0rP_q(IQ�kQ���ؠ/	k�׸16^\�F5�P���ٛ�s.�i�i���O��]C�p#�b�+`&C�]slsm1�'
�h�_���F��MΗL
�8}+$��x�WE0���33Z�Q�t�n
������z�7cI� 	�}����:|�'��}��xϊ�hJ
uW4G��T���F#��^�xB@��a��QC)�v�}}�eg΁v/�OGԌ6��0�m�y�Bv���<!]7wl�]�G��O�	��C�"o�6�ȰY����s�#��bd
��0��t\��'1T���ư�ũeXifPs{��0��{k8�����@�'T!�� %��O�+։�>Y�؞�_E/�u����f|_�r�`�T�G)w�<ZHQVD>18����c�����֫ߍ��e<��7�tE6W(!;d���<�9��V	9p�2���v T:�p�j'�8Yvi����<U*6��c�ǲ���Gu�@���Rz��jd��$�e��"%�U�|�2���}4�^���FO.R2uk�2�A��Xsr4*�4��� �ʧ"e�ZO��$�98*��Ѥ���B�1f�A'�S���<���7: ���|a�q�1�=�ޝ�%���:�{b����=�qw��$�>����>7Iwܒ8}�X�|;��m �6ܷ05����R�h^�ꡛOkkZo��1ԥ�����6�%9�G
�ѐ$��@��j�V7�?I���;	�\�BY���Fy�t�2"�1ڝ� ��d��9��Y�h���E������J��®��,3��ϖ!�~�j��Y�Yy�����X�Ljl���?Y:�t0L�J}ZhR�U-�����!� �eN������n�4��x!��{����Ni���\��8p�C���F��q�-B�>��w�2؈����(WL��.�KB}��o	E2��r��0��MmhI����0ȥbU
��i��y�/��~�)�b����e����~p��_��p��
}��ɹ�3�/�-���K�[p�\�1HH��F��Ѯ�j��4���=rHy��<�\'g�v����Q^��L�d�W�^�����^e���x�*^B��,�b-���J�.��7,$2� �kՒ��mѓ��>�P<���8���6��%V���ŕi|��Dc2���)˶͉��G�/����:����.�vfh�P���K��Ӡ��G�;�vP�	)�Z_~N%M�}|A[<ё����I8��5��Н`�kei�_��wi�;p}kns?7�3H�ξ��\;"F��Vܳ,X��m�_k06���u���ϛѨ�*��a23���K�at{�2�at�@�\9|U�I< �$�S~��NpZ�rh�n l������������)���T�\&0�~V�m�����(P֙�j�P�H���|q	�m��Ҥ���}_{?�2�����)�U%��\���p����YjWq��C?u�cz!�����,9$����T)��	�a�n_�����g%�#�쵑n0�\9���H=| A���{5���G.@$`8a��6s#�u������`�����-u}ӓ��ɭJ�n��L�:ّ�#��@As��Rɹ�-��)�=�^��eZRU|�`�xhf�h�@R���>k%�G0���G��`P
��xz;�ӎٺ�R��(j� ��*@�w#`~�s�#tۀ�|���r�^:o��O�G��edTbl�3
�d�`�!G�:񋉾�����E��J��n�.�}�f�_F�'�Q�W�B�����0~�8|Lᢄ,��l�+ (��σΚUF�Rx�H���N"`͇��h���624���GC��i��-�zfw���5F8/F�,��.����) ����v���ns����M�U�G��ǿ��⥰������ޝ�%�eP#nW��X��'4���H�${,d���:ѻ�q���>}���V4�"G����O�II!N�/}��ITY���O<�JF
ߒ_Q��ȣ��<	p'Y� ���L�{ղpn���d%p�
�_3�]����:�����V[���߳�7J��I�s:י]c�V����P�M�.�L�f`���)!,�2�q������u_����a�$�����v��kMA�3���h>{�����)�0�Φ�@s���
���7�B,�og�rX���$�Q�1��	��e���=�ڂ!�����������c����U��&ݓ1��E���XهF���6�yJ#����YpnZ�q0=0���ڧ����\�4t7�C�b�W��}
�9rHy�s%>xmȵ�2tČ�	�90��f���m,�Mj3{DR���ˇ��%(�즍�L�tI�Z(�ԉTxK����6��4��R;��a����|���9_���P*w�r��.R���`�͏"CJ�qj	u�t/�h��t��:��z�7�C�RC-�h`:���V��r�,V���j�S7,����{gr�=6�:-qb�f�V�E������N]�h4�ƻa�9��`�+�,Ϭ��F��u��;�	���J,��AQCe��\���,�?�@��Y��&F�6��|��y�r���jd_)!��3��}m�lV����چ��;d��p����±i�	'�꾯}V�o�8L�K��Y�u�_�v�К22�F�� m�q�zj�Y�/��_��5���m��(QA���;h��ϙ�y�Jj��fl%�]��a���ޞρ��Pɢasv����qi��K��q�����9��_��.�*�eب���"�mFF�uQb�E픪��ʼ8�8�r\�O�>�������C��#���7(/��[��r+cp���Q`�޼E)���s�sݫ���w'�aJ�L����ScIf�mK���S�;���������9X�8�|���k�#�/B����3g�f���P��و�!�&7�J�O��/��}�v�����5rr�(���yO���N!�E��B}\q��c�2��OWw���NF]s