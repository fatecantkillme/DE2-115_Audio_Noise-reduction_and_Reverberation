��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<�y'�I�z�OB�N�0����h�w��3�?��'�e5ML��u��4-g XM�������p۟����ĵ�����ɝ�s�VN���$	ځf���<-+��V!u���#�4`߈Ր��7����Zu(#����V�{j�d�ў�ф��f\�3��	�w_��H������&bSO�3Z��W:�T**���k�93\bOذ��;���+P0�}����ivz=��}2!��^k�e�1E�+�$��B�edEW"���J��
�\�;W�ԏH��-A0҅4kd�1k7�C�v��T��(Y��v�K]RA�P/�ê�0�����I�~ӗS��.���w2 ����2�pb�14����_�u��Ε��Mn3� (��EǗ,���H��o�>])Sfo%�!R>���μz��گ���H0?�����`Z	}��"�=��4�:��ż[/���4�z�*���Vl�xM�֙I��꺇���4��I(��G�����%Z9�p"X�qXZ�c�J�xJ�B����yr�)݈��,R�(�6"�U�]�[��W��tL�S�@�N	麧�lulplnX�dN�E̡�ޢ�@ ����� ���e� ��e8�z_W�V�{t��q�X�m�)z"�%YSt�!3��n1�*Z���%A#���؁�	7s�'����0��և4����95hS7��VMi�9	~[��un��q[}��v�9T!e�3	�.z�QSOĚ������LZ)���gAY�DTy6xO���l� b�Ԑ� �9���@S��̻��拟�5;A�u��s԰KYF��N�Q�:��6�
Dz0A�|����K�4�b�}]�X�p8,3~%���q����軈C�檕�fsg��ML��G{����*U�f�q ���	�|�yn��? _�e�I����|1��y�wAM���J�6��jg�F_a%�Y�%�����i�j�h�d����~��$�a�FC��B���l*f�|}i|<�t���o�u�ޘi��d2������F.��Yq^ӃE��A��4�悇ᗯ�d�1I܎�ӌqvf��]Y!񤹹�b P~g�%��P��7=���GPO��6�xb�[��X|�1��ֶC;Qb����=��c��fuXX�r�=������rI���������e���ہ{��:z-a׏/��_d��S�^8��U8���NYs3/�c�|��Lh�c��^a^W綒��@�dʄ���m���$̓,�?��s@j��&<�A�A_�'�Se��F���rO>)���q{.MW-�bط��<�8W��}��H_��c�y�&x��G�D �7�3�^�b9���R'v�&w�8�W8Eڶ]ܓJD�n�)&ar����`�4_��.���}��=a�'�_��נ}«ex�	|0��P�^|B?>�E#�-�:�n�U%(�)ЇnRh�NzW��]y���",�]�s����\��X�g*qNi�D�K�+�,\�W��NZ�o��cE��Mq�w�DZq�;��y��TG�]���[��q�j�G� ,���b������)��Œ'U �QZ�=_��/_%Ӽoe	���а��.�p�<d!�l.�����V])^���w[LB�Xj�ب�6#�����xz��\o��N>���� �F����x}����~sW9x���"�-N�Zp!���70�jr2��RKw�c���Y����iы'�~� =�����Ӳcx�Bn)����o��|�㎲�����l��mI�BE�V�wF.|�N_�ˇ
�H4Z ��3~A�e%�2.k����	�)���1-�H� �wb�F�!�}
;U��_����3��,Gc*���Bv.���\��$1�g+�����cvTU'��W���0�����FR�Xc�fD$�Y2[��l<G��.�Y\z褫L��F�������g�+� tQ��+���F�-��ƀܹI$��������7��(V'�wb� �����<��2�{��}�4�xnNn+dl@9ES���C����y�L~j$in	�ly%l$�f6?%A��)�����9�C#�e�����Z����+�]&��������W�lx�͜����y���W�p_���TYe!�ߕ������G37Zr �"������_�+���x�v�q&�i�b�I]���APݫ�y'�D�?�df�[��=Y�}HZ�{-ǛA`��ZB��]v;��B�VmM�n9M{�O�8��`:�}ᬟT�+�M�0k���<��0�`ۣ�k�9ZS����I�[�6Z>�î����)��t=tIЖ��)�:��f٤����o��l�mz���y�o������޼�t���(��^���ð?�����7��RA�D3/���g�2��7٢�l',${B�]Y�!�v>����!���걈�\i�#>jy�+�[L|�^��2�����.�<c��wNHT+a�ր�}SY�&�a�	'��k���8�t�rN�EI��0�85�6���T$dtx�0Y���4��*���N��7Z�G&�����H�����h�V��q͈�o����8iL#�w�{.�:�w�����߿H��_+��/��ّ e
����߶;�����������M*=���+0u?�r��߿oV|o1O34hwZ�8�qM8�P��������Z��9���r�$�3�����(o����W	�w��Y��Ǡ��M2����
�ُ ��zs�M�܃�LL����-���>��;�F�@\�i)р�veS^ֹΌ��u�5.�^���r@Vm��.ӥe\����Yҋ�)w� p�g���E�n0�*��P��~15���$f�죫:�q���Wfi~t�V��	:(f�$�**������w��mV!�;(��e�euE?[��Q�!I�(��&b�e�:I��T���Д�6��fg)��yd/�YdB�{(q;&�^ZXWǱ��N�iOMӈ
�Byg�p7���OO��R����z��p���FDlL� 8����v�CK����e��6n��E��/I)��4m�Eo����K���#�T��rQ	u��h�M�w�5��zbr4��0���nhB1ƞ�%�������O�j��Q�Jt�X%z�Y���ג�/�Y���tD�Լ$�w)�y���$���i~!��G�V0��C!!��}]@�.�I,�Џh&"<�����~7ᐖ倯�^��;��F6,j��{���Ȉ�X����(q(4E�6�n�v2s�)�H\���$�U+���V�b��j������r�S��3Y����_���<)�ެ���݃fN[IM�g*~���7zJ�Er��b)�3������L��X���N!�˥(� �4:�x]���K5)���ma� 
�<�yt��3][�@��Ɗ>�('xy��O`|��,�:"bA�R��:�4����~��z
65��P6�k�?=�H/�qw�CL:�-�dt�H���n�롬�bi/K\U,Qx�ਃ��/��tNfD����|�*?p���-@m[؋Ҳ�C���E�?�ʢ6��Z��T�JV�1���(ٵ�+��,,}�҂D���9��0ř-�Va�ľ��Y�{��hN9��q��8���a��CS�����du��/.�WC��c������v3�Ҕ���������Ŭ1I��_}f��C�"ʘ\�^��DWW&�r��͸]��u���}d`"{�	�p?��)�����II?��,e��|\)� ��.�����4�^0��%%^@�y�贅M�Ni��R:���e��J�����_�$���>�t(X#�[�38�iE��.�W�������肿N���xbB�½�d�-��7����oPC��\��I��W�J�s$4\Q=}b-�����1�w�m��3C�#ù�;m	�`ٖ��$44��/�?A�3a,4&X�.���
~:e�V|����I�<�7�7!;[�+�E`���[�'��$���=
���44��I�5����A��j��p[��Tȭ�8�]��8��sl�z� wnl��n`;������Y����J��^��g�-�h��|XM��$�r�n��e�'��B�|�#u-u9qqA�Ĳ���o��/��g����:pp�)�ɪ;��'ɜ�iw�;���6�R�e�������Ba��`��",������+k�p�#�!	���j�|%�Ҩ�؍�s+*�+��=�v�3a��N���-D˩��2�(Xi
}���m�{�!4qI��u�8��GR
����?�~p4VۇS#�Ef�ކ�ё���G�	�݋r��JD>&.���]g�V���@U���uv�'��)�y�F ��0��a��q[����h��&'?C����|��S�j*�7��8�s.��O�V��5�*A �~{!f�R��(e��#:�@��P���K��$�u�qh�t��7�V<�e��rP(zFI��LQ!}��A/�O�����;���t�
�Ek�r�J����A
 FB O���w5ݎ�U|y�l$�1>y����!�lA�J (���"W۟Z��-��
�+&�������eޒs��n,A�K̞�KI#}��X�o����Y���p
��Wg������Hk���hP��l?b�}!*�ѽ�Qjm��[�\�����+/���y�5f��?Ƴ'-�\�v�������ɢ�/_�{��w��~