��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>>�Htd�η��$Y��!��+��ɗ�����6����&bq��j�#�o���ٹ'މE���QD���0@���G�wAT�ܹ x�*�'afڱ�L��+�'5P�.?�JSb-+�D����Tls���(}���&���܈�̜~Sʚ��18]�故@����/.�#_�S&�[�FG��a�0����Q�o�h��T*��љ�v�lKn�)K$����.#%DȄ	�`O!H�c(_�}/��&@;�`v�Hf�F�����Z7�8��|dS�1q��Lvy� �4�rhșbr��J�V�Kd�:�1K�0�`Q�7�^B��#�'�9[���
���+H�1�zg���SC�9����a��)��C,ݼz)��D[��A�A^.��t�H~��4sh�-�w�p����9
�W�UF!�ZA�?����:���}�/	�R�<�x{��C����
K�V��r�4���cj�օ��Rk�T��g���V0���?��0�(t ��q��q�Ca6�P���EV�8����E�\N�Tθјu�Y�9ߊ��"Ge���5�uB(�c���Y�;T��wS�(i��2����\ì��QB�1!z/�� 7bZ���XYhRʦ�Ɯ��~)ӓd;%|x��N5h$��^@�u�#_����^��&6ǅ��qi`bS\��W�;\�O��S�Aq�1��������.��@�7��à�HwE��@N�A����>֤�8��m����8ݐ;оA�C�]��
:W��w������@���C����Q�(�⠴�x��Si���=mp��q�_E4Q�N����x|?���Er2�G�ɹ*KV
F�&׃�<�	rR�O�*�K%Q�tİ����BP�����T�v�z�Ò�����7S�:��u�I��?T���ݑ��n�bO:^g�?A+�c�j��[<#���ES��112��/�76)�F�~]��aq[WFM��f-���Kh�aEX_�V�� A���-��2)!tV_�Ȫ�����~5~�K?�S:t?'�(O��������c���Nf�H�Bz�WHa�c.��t�$��t4���|�D%|�:��S54�U�ުS���B��*;���؝V"ū���h��I	��	��K�q�Z����-�p��Ϝ����s��n�ƙu?�����&�/_%��j[W�lY.�z��c9�/H����x��E��y�k+��P���x���p���w��;h�#^7Q2"�4��j�`,B�~������e�3�r�����fw�^Dz��<��A=U�����͝���L?<s.�����jYzt������.b�����j�$�)S�s���Y�$}�����)QVɩtԶt;�j��aF�IGқ� �}�^�!a��i(_�36r5��G倄�?�tX�� h���8�v�d���&q�l;ܵY�|�~�
0|z)o�#�4$	��FأQ�'�d�	��!151�-f���Ƶ@�
� H�OB��+4��VMl����>��4��HTG{/�+��Ss!L<o!�M��.ff>�V��o�ޫ�� Z��w�?�>ܑp0����`���4�qÔ��S*��3���ğ��X�a!��P���]���	"t9<�糺]�`��/19ʃRN8�Ģ@Ƞ�H�W� ��E( �|	���\��dZR/+C�+�����vFܯ�ы���� ��t�Z����Z�δ����w���3	mg��*��n�H	����X����Y*�vC��a�1ؤI
�h�RU|V1�fo���$�j��/�oR���� g�S�E�0��>��o]���#�K�AD�0�k���0�#�%%��*$3�h�q�7_�Bn�WRSd�Lo���2I$�ԓ�u��+���2Vr~��[Ν��A���v��0�aR�Ӆ�
��w�B)P�yl㬑�x��F��	koL�Bj���n����4�b�pF��fz�!Cp�q�vl��� E��W�c��"ìHN�*��{�D_rڞ4�:d&�.�`֘��eb0O�o��+�)��Wb�7ѹ�,�L���/�_��(W�k|݉ȍ˦Qi�Su婺�@s��f�@��iȱ����&��Q�؜��Vh.�~�����������\��[�)V"�D�\�9�k���y�6�"}��������~�n_�+Η����ʜ��q�yz�ZI<"�T�AXoȐ8b�������I��Ҝ��<Y����b^��-����P���. ~K��s'&Y�v�F������jtI$:d���>-�J�mk ��_E.P>H��u��q�*N�<U}��G�������G���э�ϲx!�n�TJwE��ˎ����ߓU�G�7O��?v[�й��BxD2O2N�j�� �.�C�ί�վ�}k��
�',�R�� �nu]F���c	�xk֩���҅�9P�}�1�����,@��]-�7��MR�)�yo��-������ɜ )�r�W�B���U��F:�j(���L<A@~ELW�6��c
�q0@��-�JNJ�tb*�0�T\�H(�蓕�X�W���x�p=��X{r���ߍlg#�����q�Zoc3�l^OZLM*Q�]�3-+]�)d��Q���r�	|��3�#���g�.�@*=I$��S�&�(:&���u �����Կ��ETG����;�X$6&t��>;B/J�=J]��_u1��`���L�O7I��2�A�Ҙ�N1�*5�خ%m��y�yt0��س�����ý���o�&�d�(̪YqR��o\N ���K>9X
�7�k�4ɱQ�t���IƮ�@�QiL��'�V�]��֚G��T�.w��>fhj&А�<��
�1�m�{�n�A{�y(�06�g�?季���<���S��/�D����l��
��������s���ЈR��L\��.�r�;�8���A���B=�q����f�]΋��I��e����*�Ȯ^��r\k=:�jZU�T6���O�D�[��P�QS1$ b�	�i�)�%%,i1���R���T6��fo�]W����Jb���6�`[@��|D�aM�~����>�$�ds�7U4��F�6h5�7C��Me�gP�+�~3�0pv` �n�uV��c��G0eH���=�I����zY��m�4SJ')�p��q]2NlN�����ix�+�IQsM|Ü�W+�p�`I-d�����D�b�1p��u��R�L��$M��`��scĪ��Pǚ���47$�i� �&.�Y%�2��liX�����3�W��fe&�4sI�ϛb¡A�����}�H���t����,��