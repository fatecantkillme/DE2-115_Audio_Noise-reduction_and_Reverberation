��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<�\���:�[��5���zM�vd�G '�^e�6@�6��-=kv�����B��e-/b|o� f���N�	Y���+��PwEՃ�'����dB8�l[���fMYE�7���s���/��i�Ŷ��И�;CYap�1j'}�q�Eq{L�G����� �oJ���4�AL�2��źzL��XA����sƼ��(��|�.q>��V��$���!�����O����i?�LosCկd����p5y��V4�P�#��_���4���䰤�|Q�f��Q���Ъ�j'۬��$G����*���Xg��~�9��5��%N��'ĜԴ�"�_��|��WN2X���:�����,�	r��m
r�>F�����7�@TX`�л�*x)�jD�=����XS1!��ɴ�4܉m��v�j�Wy�:���F�69����%�.=��\�+w��͹�� b�� }��+��&����dx�$�[8-B���)+�*<j����T��u�&_�[%�>�1 	���2�,��B�O-V�E��<e�'���#��i4��w�b�{+�[&Q��N� �֬�Y5�&����I��|�k�N��
q��sO�`C�F��5̕,������j%(=*�AjMuF/e�o]�p9��	�\�p$��Hu�%W��`�kk�V�cyxv��|R�Ґp��e2��EJΓ#h���wá�@�����V�zl���hVl�/���'
���us����9��)��-2CJ,c�޿�ǘ=�2^^�P�f����\��	h	<KoTx�2�y�_��Z:!q^.��Y�4���o7�]<�)�.�������N*:t�|?�v���X/n������!��Ḇ��XB-�3_����D~m�8����6P=��f�W�����>lCʺ�AS6�+)��nu���V��l�W��c�O��b}�j�;���$�hL^�ǎuj,����*B����IѢ�p�qx9�+�"�$R��0�r��XV8�k0�K����@�Ȑ<�s���=���de��WҁW��ߤ��&��,,�^A�1Wロ�n�o���e��{G��NU:�ƕ��R5�'�J�Zb8aV+���F��!��$BzAK���7�<�ZH�&d9
,/�
3G���&���{����C��<e�����{��Z����ǣ�s�PuL��ݮBi���]�M-�B¹���c�~��^2Y�<���3�L�� sc���v���+�:�e=�ч��v"�SZ�)7�(7���9�'�!p���J�K�Q�Y���ӦF;`Gv���·��h��o�����@�O�h���u/O�I�j?P�pmKd
s� d#�x���Q��YMۤ_�2M�:؇Ղ8}�7�!?P�M�|�.f�?�uy|U��m@��C��Y�;,4	h�)p�f��~���x��?��z]}MA�A$���E��R؄�}gQ����О$�[C�{[�0����Ƒ�ƺ�dɜہi8�b�O�Lt~��;������� �iW�P�V��7U�*D�ۋ�Լ��^1tp�/�L���r��GK��#x���3��9JKQfzf�y�Y���n��cV`�a=�jH7�Y��Փ�@��ɣz"qγ)Q?4{$q0�����>��2.��F����h`
�:�p%�b�+:�<��6�y�!""(n��A�a�����SV�<���G�Nܷ�P��`�\E -�[۝lT#r���.�pa��#��g_�{1�W���M���dgK|��F�O��5�՝�{�g�u�,͓\KX�͑`���_���/��(�p�S!�-�C��N�ie<�o���(c�8���y��}�~5.<$`�B�+��B�e�VL8���+�xa��a�Z3��q呎�7��4_�vM��1?-]���4�>F"-��a�Bt��J�l�TF�=.�B>��~�[� S�g�����C��cb���#��QĹU�O�>��Iʑ�$
��PT��q����]+�G�=����8i��$1SS��-i'�����Ѻ��Ra	�hT�E1_�"�6u�:���3˙�v�'=�Q�7�ߋ�"��yv�q��i�z��FLn4��'a2�E��YFߗZ�-�GE@�P��n���~$����{�C ^!X#��0 �:9ث�v��X5�X��H�S���u�� ZΖ�OFK3�[�D���f�05gj���~&=�r�vBd$�Ӵr����"���5����T]����Y�� ����o�S�h��a�O�7r�"�p���M&]<ts���!��4�4��+d]\2�̈́�8{��S�?|ֳ)Es)�ƥ�0�6����o{�^�㨉r(���� �*sY�������<Ƥ�(�T�x4�sܼp�I��y#��_��\�z=�^���E7��Ǌ�J�T)��3hw�����0y4Z�@�f��g��@�R �a�"�Xh<a����t�U%F^
Ȇ�{����8�#��nʪ0C/(�%��9�\ۅ�q(#�����Lޗ�T�\������.s����N�����
�1m* 6^�Kw�p�k�2@8��D�?�Ť�띟�K�R�6�W�.�i,��]�&��:s҆����R�;�`ñ1����K�rb8�s��z�6��Hm񾷙m����L�|�g��Onqi��Q�E"$c|�q��F���1U�l����*�1It��ӻ�=h���U`t9h����CB!�9~*����ͱV��
�&؎�5o	��.��v��> uѪ��gnm@�a�m;7�������Q[��D�V  63�G�E���
6Q!���j)�3`��B����BX���H��d��<^O�� ���A�k���>4>J�|��yj���x�����;txH/_e͘
�����h��#CU͒��儎�� �������|�}�2�gʑ��V��-�3R*ܢ�����8`MW�?zףպ���L��'N&H���~@��.F7V���d��hxR���=�Bb��m����7y��'T6ߦD�x� I�=�>��_�ѣ�`��B����ð�V��+Y�\� ���忇��Ĝ��܂3��$�f��o�4��y�u�o=���*)�|���]�I
�N���\3�*�f�*��@8��@�z�f�$��yf��X�ВK�Ƶ���ג��W$�5�9Dd��^p��/=��}��4�g��E�}߬����U�X��	ڼz�<���\������� ĳ���@��wI�՝ϼ�'���-k~�h��;�&/@�g�7��-9��[Y����q�C)3�Gsq�2>��T�C�0�+���j����\�얔@��}��<殿o|�|<}���}acd�<��{纳�0M��A�>d���-"h�E�6�Jj#��S0g��}n"��Ҥ4��3'���Uz2�\7���^�������+���eo��I���j2i���#|��{o���x��E�{J���i�.Ƞ���­��^Us�KM��.ݦwq ++w_��w.��h�[��*$�&;)��f}{��q��+�����볧}��P��`��H*�q�r��5�Mh�-]Z�*���U[���$z��S��v��C4�Yh����uJ�U.41t$'۴a�'�eD��h��;^��d|;R8-*3�1�L����|�������BD�x%.B��wAQ#zR���Ď>�FF�'@^F���w%ڭ����}��jm;90�ѯ���`$�������:���T^��6�$ر���o _���J�f���Z� �0�:��A�p�2��T�����g������j%S��`�!߅s�ѿ�uz��<?8���E��僎�26�#�����Ҍ�o�v����f���������HX#l�g0ZHU�a�M��@<
�5��uy�Zڜ�jv��C�����p�ؔq�E���"`8E��� wdK�t��\���F��F��yz�L���k�?v$?���X�{뙚׼v>��F�+ܴnhhh�1Mw�]�Z�~�n~���
%�����ꍆ:1)��źw�9w�- {t莃ċ۰G{bSI�׳�ͷ�O�DZm�R{Mm�� ��hlb�N�4��rTN�d&dw����	��B����'��͙���\�Lyť�\W&����s��:
&]2��.H��p�ă���0a��-����]g(��'�,�����6�.�I�IU�&�䥂>j�_�$�R���I[���4�t*��͏ߟ�ߞ�c�����f�}��s̡,�ݤ�����Ӂ�}/<��Ҏ˒�t�҂�!�"��;ϰI	��`w1ISi�+��@�6������G�Q-����I{��:���2��� ���o������2J�4�,�Ii~�'nL���ڟ=y�ҵ�/�!��<�ܫ�"K3}f�4?��:���p�5,�%�#�%��Lދ�SM,���*��$�U��ޥ�o����ݲ��ƚ0Iz�N#h�#��7��U�֤X�M6N����F�l��q�p$�����Xi���f<�[E�����f����rPd����}�yA䨴�����<&%[Di�[��7D!�.نc��t�����u׆�T�K���I��hZ	&��f�ƒ�:��e��F��O��O�+�-�i�o�[���]z.#޼J��ff̪��EH��Ѻj1�v�9��FO�@g����<�[䫪����K^ ���9��0i-�nde��(Ġ���m#l	������ȿ�O^�F$M����B[���@A��Δ��krn�.�
6.���W�NC�Y(��<@��0PB�r�C.���H��o����а�ś���@�_���q3Η�:D)@�{sߟ��O������EF0��f0�o~QQ�;�g�{²�Oj��wC�n6��4�ҾPЁ�|9�p�a�Oh��q��,�&��2�����0j���=�Ǡ%�Y��0�d��}`�ۘ��o��{�cg7`|�����n��
9��UNJJ[4��6~��� C��Fs�?���� �YMM͍�%�ع��'�Ѷ�h�Q�XL0�K>�j���j��0?ɣ?���b2%2#8�I�7����wڤD�I�J<F���-۲���Q���a�`t-̆�mQ�Y�se������o/��]�G�i���kD=h��_A{~"ۯ�6unY`m��̘�s�	�N��ت%�y���V���K��C�>p�0�`Fx	�ҵ�����Lm�����,��㏆��U�k�>Pg��`~j���Y��U���u��3�����Gt�\Ʊ�W7z�y��RƞnkF�� Iu�kvnCV|��� \M]�fY9)��� �/���\[L�[�(G�ҵ2_s-�A8�!�rv���|������R(uDM���CkF={��?��'#)�
������qWj��)>wr�){d�aͳ��AfJo�iM+;i.r��1�~,����4���(.�e�u�b�\�9��������T|�DL��1����g
h�]9���8y-�X�ImK�YOu�oȦF� t��V��FO��7�;^ؓ�	?K��T����.n�x��c����0�.*�V���f�jt�8�0r��^w�~����E������, ���B���R���饚�5Ȉ���?��n�,���lew���-�Ui���֋Q����>t&��E���
(pK��&1�{K�3��1���c���p�dp-¾d���{�#�	I>ӂ(c�q���cy�	'�po� �D����9������Wm�Y������q/���J3�%9�I09�]����!Q�b3�I;��50UZT�I��e?�,�=��"5L(
�(�wS�22/x���k�Ypf�
�cNVʭ)7X�O{���t�B5C[%x5t�b�+������^�[c�h�U7���k�:��
e޻!jNz�Vʭ^�wi�����{*)*��|a���-D|�v���H�ڹ��H k�Ǻn\8��rԃc�"�mG�<j�c;�F�?�J�;1���?�Gdny��]5�����-�������},TL�^JL�w��S7"~k�aa~E��ȯ2yg�A�g ���aj�js���!�M��0K���G�SH�'�WőO�uy�
}�C�}�/�գ3��4���<�"5�B�$�t�XCDB���a׷
?�XF�'W�?3`l"��NDjU.^�œR�A�mY�ڼx�?�s*= !�OҌU_�>�y�6$Yj�H�ך���`�
PMw��E��*D7Y��	$d��@A��M=�ʫ���7�Jf�LG��H��WօO^��nVf?-[�3D���M�=S �`}��[IC$�sNz?��[K��9Z�H
����VT]�N�Q>��R�7���-	UmlS�,���]�,mvb�4%��Nr|��o��;ա�������cW:R�W�� ��H�C�GdM���W~�e.�;�� F�V��耋g#��l���4=�� �e�����=���[���E��ڕhU�{�F\S ��d4kl�Y9Z��A.^ǎ�It��2T�F�gu�7�m����)�_��ΖK��[~��+:N.��4w2��I`�0�r<�P�]��`�kJ0��G�d����K n%q�C��6���f�h�Z���\"6i��o"�vN�E�@��41�b*��B{T�6�;��8,`6�׹�N�Aif�DZΚ��w�H(�Y�X`Tst���$+�Ƭ:?��R\��4�5��۞�J��1>w ����)7|f��⦋��C��
=[�r�م��z1�s���]y�-�xX��-��	vھF�}9J�y�&��mYo�s����^�B2;%e�٪K�1Ӕw���ny_� ���ˉ)^el��ф����"�"���sG�iĂd�h�A�&}d��(�0�W��h-N�)�\m�a܆ج}����J���N�$T����7H/�(�o<�]�$*��VK��	AlZ�湥�]��Q���?��v��˧H��0^�ohsB�2���j�9K;�%��]�[<��0Sҽ�ݧePx��#bF��3�,��kSd� �,��]т������#�R$`,�̿�s�z�.Ǵ2��}\:b�k5����V�x~�bxZw�P�n7C/,��o�B9��`ef );�D��b��D~k
;vaLr1C"��z'��O��TF_e���tK�Ћ7���RU�]��qu�]9CM�bj��H q��{����l�*2�}��Z^�?�+A���t�H�QD��bh�;2S��;��_�|��� u}(������ꓢ�lOE��Sl�E�B�O���pI��K�a�%��G���2���d��_��F������ڽ,�e��@�c�a�K�0/1��
��x���2���EIzgi����'��+��(�ņ�U͝�YO�Q��.xl�I���,���j�k8�9�T��l����a�AƊW��K��<k�ڬख़�؛ Z�r3eȡ<&��J�Li������u��=���}��|��ܫT�i�������pW~1��q��?�?jy����9�+�zԅ:��2d����%MR����Y�Vp�N�Qx�?����KX�V��!WD�|�A�\�C�V�f�X.8��?ύ�l^O1ͩy��p�
P�yi�y�F�C�0��,�N..���1�@�G�	������	��á�u{�>��L�H.x�Bcː��FA3e���{tә;2/_X������!�r�zi"/O�!�XV)�72��e�g%�XߚSG�N(;56�7~�iP��E-�B(�Gs�8]�6F�Z%f.f�;f��=y�0�»�I�_���Y'%�˿bO�<HTL�H������]v��.y=�48�v��/|�Ph<W�K�gb$�?0h�w��+���Ї�7ż�&������!���r���\=hi7�A�q��M��k�I2o �DKQt�(���P\AF}�@0(����|�Azg`�%Jɧ�[��%��)�ML���M�+�<�K	0lߒ���y<�*���>�*�1U%27vQ�i�]�𕨢m�ŽGX���	B�tj� k*c��f�YgBԧ�oq�2�E{��,�&���$@��02Tȴ��@1�d��C�_�ǵ��`�ܻ*��+���!�M�[|w�T