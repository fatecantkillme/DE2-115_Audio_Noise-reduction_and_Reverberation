��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<��h����B%����!�VpMaI�n�7�ˏB�O��'1à�[�-
�3o�+�|�G�s�ۿ�����yh�yЍ֮E��FdsVn�Ӿ
j�T�a[l4�n����a�$������َ}$Op�]�T��J!Q�D��-�πy���so
��N�����؁o�%��A�RC��o/f�0}��/d��p�&H�`;��#VP���y���e���/�"�#1�;�G�cv�uM�Z�����pDs܊������Fe�z���kÖw�/&
,��Ġ�|��񗴳�	J��p�5<��"�:E�ݰq����G>�wd�KH�3������'W'/x�����<���o���6j��Q�v����X�I�A`}�1��9R5��,���tQk�\	Ȅ�mI5<��h��(�ؿ� dB5B4�MM\HW��F%��}�˖{Dґ|4��V1w���d�&�!O/����S�Ĵ$3��M��/Q6���f[����Z���$�O�>S�����3r�E�P��l9���H�6�P�r��@D�~�:=��*u�,���Xb���i����A�%�7�ʬ@�����qr�be�f�,�S~��K&�'�ܴ��v�l�}E)1N�a@m�#����m1�oN5p��Ƿ�0hYg;�o�^`����jدS�f���^�ED��&g��2+�e�u�gv��/9Z�F�#h�@+<��IӧyC2����.�3w:�\��ubE�ldw�Tb�P_�8X�C�9y,����R��|�$%e�Ј^.����� ���MM�ӗ:�h�dI��Ǣ��9[M��*�ݑ��������;��`@��!����7±vO�h��S��M8m5b�vjv,�v�u��T�Eu�������7vW�P��8�!/Yy��J�st�7
�fTw������L،X��}�}��1͈Iw��[��>V�T]Æp�\��U�.4m�7�￣Z�9ͧ1KRK� �w�A!*Űⳗ)`�2�(ݖ��b,ӟ�-�>b�W�+^+/2zFhg�kt�J1n��� M��WM�) �o^9��h$�Ne�"p/�}#t�S�w!?V[�8KK�2�r���m3J�Md��ej�ݣr���II���#y�![=��fu	�zN�K����		���%���ᣌU_�W��T�'Еs��k/2�c*�ƌ$��_i��;)����H�'���&��� z�կg�:A�l��x|3*�3��&)kM��s�e1C���A��1єZ�{��4Bkg��s�S�Q���
�n�n�X�F��F^=x-�S�tw2BoG�Ӂ`<����k�s�g���6ۡ�+D~���ňD0�����Z���1��Y��#�%�"]<�X��������w�$\���-e����rQ$�a\VĽ��h#�.�ץ�7n,�܍H%`����Z��7(��Q_}��6@�2h��@&�ydI)}�n}Dio^~�g�W�x��nK��:G�X�࣑4�.͹��`,c���mh>��q��tg[m����D_d��T�D�օ�JQW��V�zt/<�|�#�Q���'�{��lg�j� P.7KM���,ς�}R�)����oa��{�En�m7��Pl�i�(�P�%Dg�XY�C62 :�ڑ���,wU7�9��#�� �ٿS�m��^�6gy�!;�4¸E�L�.�BaFއ�YNS�s�+�zf�	P[9KK%�%�g�bP���7�����B�o���������7f��huߎ�H���$n�b������Fk��t��J"���d~{I��8�,�hLF���ç#��]9H,�ZW��$��a�M	�^������/%kaKc��J��t�L;�KH�~��K�xc��U�=�!-��<i'���{m�`s����.I�'��0_#%/���:�D�hh�Y�3(��LF=4Gα�^���V�C�&�!��TF'|���*8XO"0�v�,9!B�^�@x�L�ϱ����H�Zv� ��`�����'c�b �����ھ���h߱�����!e���F����	w?���옰{��G.�U�f*�b�ޛ���2����j9���>�c[�'P�Ǧ���KU_�F���S��*��0�������B̃�g7���0�|�u��
؜��i�����As���Ѐ츏��Yt����S���h�+З�,�� �X`�
�c$l!��T9�[�&�r��v*faT���tf���U��]�t����z���O�3����'Ǧ�2h��m��@(h��pni@�5�r� :u3�[�ᘗ5Z�pn�B�|��6&��9�=�� �dH����r�Ѐ5�j����1�^~0��[�!�|�M1��y�5�!�;�lg �Ȼ��f�2^�w&��60��2�n���^d��С��;>'hl�����^�ǐ��w �p�/(���C��菥j`~X?��y���Չ9�Q ��(�B2�b����֑�[)70��r��O\���<V�:L����EIi�h/QM���V�ë�*��s��eQ@x=s�V{�]U^B�Q�6� �� ���Z)6$�1L`d2��W+H�<����G����J�x%� 'D熟K.�C��W�ð]pRc9Y����@�Q�\�\t��Xf���!_�|��l*Db�:y�M�ܱ���|0����%��x"��[����8��'zcM�v�?��(� ���J�F��u��*�K0�����R)/(H��H"BöP]=�&7%Fƛ/!�J�f��������(p�
z��.�Ț����lU�`��K:��ry�9�R�
��'�x�z���9�?�+��eK��XKҺ?�GF,�Q����	Ih��dk�\C��!�M�a	����Wi
��}�:`_��I�}J�[�-���d�7�ѭJ)�W�=àd�\\DԜ�R�lW�p��*��a-��t��4�&�m�Es�T���?��N�ؔd��{����DoN���e��TWD���͞���hQ�6x{��2P"?�����op���.�����r������o��ep�"$��1���C�ɀg{���Q���~�� y�R��ĺ�E�v6%E2�'���m��-�v�F���Y��u7^u%�A��G�dY��,����J#�}�����O3M꠼d�1쬙3�ʼl7� )�kF,��P
�/���j�_���:��5�$���[�� �R(5�rqf��Y��d�&]��qv��y�����g�3���J\ot�J�؜�p�0��8:�b��;��Zڎ�X�� Z��o�@BFe�%\$ž�0�Ib:�28����݈�c$c#'�3yp�#��nw��K�}v C>4�ko��Ы�X�"�BʿV�!�9��9�A ���&��{����3^��ر��(��� ��6����^<W���N�ĭ<n�Ў�q0M�Q�9Y#����񻱿�� ��OkT�An!�w�����_�{��Uݹ9w�A[[	Dɨ�^g�>�1����<z��)-��-aţE^���N��z��A��Vi�63
Ӎ�=7��_���Ū�2�ҳkw#�1�I�6�o�ɉ��}F�N��������r��|��m 'i�p#+�z?�<�DӭU���Vu��(�P�?�S^���o��h"�
��Ny��]��q��R�=2K�>�[�(%v\� �q���<�a�=3�)��ȹ	ݢ���4�(W��n�Er�+) 8�F=u;���.c��i��O<�DR��� ���,�@+hŒ�>�y@� -���Ţ�.��i�o�9�ݼ�b�G��!���p��p�a)�F0ԗN�߇2~�}��y>�s�VIP ��w�#Eg�ŴjU��'�Dy�a�C*��L[�%�q8��dFd/�&�mm�A�|l��[��=�m\@3<�z�U	h�Mn�63�ˋJk���1�׸a���Sb�z��v�]��F	�y[�����Ѐ t�l��Gq�<�����)�>�'
b2ɧr�f�I ʎ�4�N��]#���>`h�h�,��9��D~�5e�>i&cI��!찯.���~-b��Ʊs�n��~P@����8�i�ڊ-���J1Pp^w$=�T�[��{����区�:V�Ķ��[N<�
)I��<HB�O�'(�~� Ȃ_�1+F*W�$�fhd����<��(���]�r{]lvz�� �F7+r�o�
[E������t������a��n��p��<o�'}�뼘�f�F_��n��.����X����₺�˨�?��jǴ�*�Q�����������r�5�P"�x�B�P�������o��c7������>��F0E���ɓ:�\�Z�>�~�����Rm9=����˘�Z�5UƱj�&w�����Ii4���C�ݢ�h���?��B�J�t��R����e�_&��p���G������<m-�e�p3=i�"��[�%��;��~)�����1��Ѵl�Ģ&ж$B(�t}�ZP�`}�Ƽ��ΓQn��/��א��P�3��5'��>͌hV�\�u��`рn��<Τ�0�|a�Xt+{y:x��M�2�B��`P��5�T��`m\���Z3^�ʨ"{dG��CsF�GS�|K.]#��rލ2�'�d�,��=R���x )$ylnU��D�f����;��+_j������� �.�\9u��U��0�����Ј4��0~\��E~�1�FmI"!0q�q�v�2g�s����Ҳ9�����;I�������'Ɂ��:6��_+�y[��b�Ծ@xc[5���vL��F4끬E���oh'UC�@�ґ}����	Ju.wq�Zl�:x��2����"�r��ec�])P�P��2�{#��n̺w��ST�}&��AbL{�W�Rρ����x(OB����>��<���YB}v_��	���&�]5�|(^�l;yK
x���U�_'3Iz����J����^BH�~h����(�`Z�6�X=UJ`;H�Gy�gMXtƥ� ����	�_n��\;��MX��z3��g�-��	����/��(�}�ɋ�Q|4����l�֤������'��k��A�幠4N���g�ҀX+כ���R ���+������z�^�*�{r�|)5��C6�g{�8N��O
$�6����BM8e	�6�A�܆{��@	����!�GD/�	_?�8nTϯe��s���ݻ]��~�0{�#��V�1���H��#�� MS>Ż������w���u9'�T�q�����Q��}4��{��	
�zۧ�Bi;q��`]vZ|��Z#`����Q�2Ha"B{�|��(K4���7إ�G�*[�9�����M�s��	2�bHA�%xQp#��#,U���ܫ̀���%]�i�4���,�NpNt?Lc�m(��<!���a��R�~�J�s?�O+�L+�E`(ܞ�{��I3O��Ƞd�q�h����H��eF��=u?�n���O������K	�=�f|&I엃?��eE ����;)`cS+�lLr�_��3�竏+���t�e��	XT�w�!���8��:��#��d	烆���I͆Z�7���*W�Ȉ}� ��fP��(}6�1����g+�۞;��q�=���^�g�F�6z���k�28װd,�Ʒ��%^� ]�/ϓ?��o�{�����_n��AfB#�+����?���e�kW��_�Zѻ���XK7�R������F������m�kՄ�Q��g��0�']������hO�a�$��ja��'�{���Z���}D���J�d�j_�͟����f��p�)://b�o:�o��?��
�h�_���$Mef�P[���ʍӟp���w���<�lD��t�(�-%W���Z\�P��(��g׫`2�mf�@���F���a��i��S�@�����'urZ�u�n�ԅ��H���R����ֺ^֋
t�m|�.-�=�9�\?4J�m�w��;w6��g�38ny�M%��N1����4ˡ�E�#�V�yDȥ��K�.H�C�p��0Xl` �X����I�f������`?��m|�\�`��Qt�����<��FV|�t�+͜�h�ݚ�D��Hgg�s|&"ű���>G7Ʋ�CĒ�V��Ybf���=\��w
F)�?��G$/����jT�HZi���'��9��1�x�s-u��c�`\q�~LC ��1���'��(Ȍ�9]\C�C��8ն�ڰ'[Q��Z�� wI:F'�hp�`{T�����}���9ݶ�P�DD�	��V�A9����E�R~�R�4�-�L+�6��@)�&�ʧ*-��A���]���V��y(�؎��2=r�k�Lσɥ!�����-��;.~2��'Enpq1�y����E��/!3��Ŭ�cj�|���&M.�!R�h�̃�R����]�ٌX�Æ��~e�a���B�S��O�B	k����z9"�r�"i۲�t.!V5ܜ�
�Y�X��	Y>�
\E�\��QaZF�
�Vr���-M�M2.D���w�D*���b}�֜�G��O�"9L�(��1���؃ʜ��[B��v�*��@��"y�AϽԇp5��}�b?�\�2��g�'+�����W�*t�����	ǟ_K��w���>�1���Ny�K��eb(��L�_�?�!�&�T��&2
��
�جx�q�
kb�?��I�Lo۠�aߢ;Q��)V�0	��� B��c���� Ӭ�o�VSVӴ[@D�(%��!�ڻ��,���2�L	��m�������Y.| �Ӥy�0�D�����+W�B
�c�w�|����+~Yk+�N�	�ϝN��{�j)��C�J9a:)�F�bW@+C�����N�[ƲF'�6���Vp�4P�vҧ������[��ZK�W"7v=Zp�R�D�W�y��%�ąo�N��V�ǆ�7� 4�+�,�eG�:7bKJ��>��{���P!�ΐM� $�!��� �|�V�w�W)��o�Z��1��fx?\�P�U~�"�E�ɀ����>��{��z�9�� �Z�#��V�J:��)������tӄ�Rh��e�e�Fc�)��7�*����_�˂&<K.6�(�L�ب��W�֮~f�8U�ti�c�.Ą�&���B�)���v[��m�����F��ݠ�iךtH�ǆ�3��׉��ӎ�="�O�	U���qtJ����a� ��
�/{Vq7���:��^0��:-�����Q�H�*	
Q]ם���@L���]�cx{��w8���=8��[��[|�n5tŮ����TY�H)H�z�)������mK� ��5�pƗ�����Mx�-�ډ��9�X�0���Q�O���r�;@g��]2�ع�{R����@�.X�M͉^��v���q�!
@7XE��vF�ޜ����Q�$NtFWX�UyJԜ1ҫ�c���hM���jEo�N[��e~:?�������zd����hoK�:�WW�r��߸O��f��;~�zA�{�H�̒�G�%l�/+�t��^�8�)���Ɛύ�8}%�S�ub	]���F�k�����(zH��4��!�V�;�5�_��Q��w���93�XT����7�0c��9@�j=�U�� �g���?�GF0-��H��D���x8zC��gj���.���8�;��� ��Ԣ�O���L)�L-Q}6��4�%~�d- ���t�4o=�}x�|r�Pds>Z8��<!5�8����.�>�J��)����.M>d(Y�?�����t\�w
༙����=b���xԦ�j�SB�J/�;?�e�4[h�W��\���Dr7.]��s����Rg��݇Y�-���
}� ��MG�]%MV���cป�JmO���~��C`~ŀ&,�D#�nv�T�;�D�C���f��C!	<���U]�=3����L�%��f�ʨ�.�$l\4KYt>1O	��*ڈL7l�ʻ*x��͂*Z��r��`[���@/�+����q��	w̻[�w
i�̳�X��3Pd�p��	���
�oz������d�S\�+��b�1��x6`�ML�C�lp�F�AC�qx]x��.��S�{�����}q������ߡ3��j���䟷&V�p:'�$��>H?UR܈ɶ��=:t�l%��_��=���"��#tm��X�siFʉ�m2��#e���uu[�L{Eك&��>��:%��.(w��0'V�*\�KBH}/�V�_I%G��W	�e{�4�i9�wJQ��#���S�۝�T���>>�ƴ{�Oy��W���	#����9n�Y^��`�,+�*U�G>���*a<���"�r'��ړa��0ₛ)煘/U||�ǚ��*�.�EQ�d�!=�~��ꖐ�#3�.{����#wl��U�ǢR��(s�v{~Et�%
},��C����KMy�o�a���a*�l��9D�r��T׿-qeG�L%�a��9�;�F��"��R��)9�|�jwsHlя�g���Ѡ���W�N��>ه�C�M���{����v�(��q�#3{���u��Ci	�wu��$�I-;E�#�&�gDڂ��L�gQ�?������@��s�;'g��zF$���Й`�J��[agC�(wʈJ��fd �K��0&7Q ���C�!�8�ƴy�Ϸ0��#��E�p))O�iz������Ė����?��p�g���M{�3�`�7U�1��Q�Z����x�2?v�S���*��wm�sq&	�<T#�ޝ��u���n�:�q�������&HlJ�U���
z�x;id�_ke"�K�T�{A �#8�Q��\7�[T�y�(�޺o�����H�]��C���$D�x>���)�����/�m�g�Zr��a�g��{��,���u�r��P��(��Y�κW�#��*8oE��E1-�����GJ��e1�Ju�����$1�Լ�9�#ol���W
�v���̖␦�.2�Z���n�n��]�ޙ�3��6�((_��~�� n
�36���k(w�L��� Q3����c�����_�[�0��&w�Ƶ�yd>��裐|�C�9z��i%HK@�{G$P9y';��]5�D`ݲXS�s�FI���m�66���z�8OQ�ʘy�aw���4�OQ:�5�%��V��y��bn���>͡�	�˟F�f ��I]���D��#���×��|�Y��҈4�y4�2r����K�c.�e'h;��{ۙ^nx��T�ކ��7Pr��zj���fR���M���K2����J�Iݢk��h>�փF4���Ls���*J1��배��xS�άf��h��r� sj]�.��kX��n��3oWl�u�.t!p�v���R�o�F�ࣟOj$�^�~#�A�HŇ9$�Rm��ђv�)���X�>���[Y����N�/��6M�M��'aDFaY�@�ey3��B�)�;?�[�+'DK6���F���:0���NfĄA]v��f���a�U�W���e�"�0���DXB�_go��nS�C���Y,f��і쓅|�\Laͼy?�H1b��sڋ�W>D6Ռ_��<���p5�4��,9�{>���̸�&�Q<��rs��k�ck,gv��P�Ϝ8��5W�HiK,p��	M�ʦ�[-��ЃP�x=���-����l����0��ʄ��D�H�4�,m���V�ǲ��F#�J�#2z��!#'<۪�5�gc{1��*�$�IG�.���yrڻ¸r�ϒZ�P�Z��PH
��3ʲ&\鈄觔|a�2��Yv#-ҌN�,XN�D�h�IjŖ�̔h������Q0#��9��w"��[{5�����)�HWK#�����{|��R��5}(���?%o8��TwwL�p���{��2��3Zi)���&݊�&�(d��M`m<�{���wz�᪫GAʽ��>]�s�{�z,�h>�Ěh*Ъ�#��mWEٵ{ʒ}��2��� O����%h/$X)w��p�!�G�)\��}`��x|m \�(�SO�P�#.T��	'���oIs��>�a8ȯ%Y˴��E��? %�-�̢��]����jP��:�C~�5	C�TEO㠸�}��:a����	m��ĽF$��.;�>d4��b? ;5O��F�'QU���C��ޥԞF[]y[w��@rм3iK�s���i�Oc������=���ב�6���&m�Gq�Gf�\�c�S	�(�$XzcP!���q0f�u��
���p�#�.x�u?�q����8x'��C�DMQ&�uF�������t</�&��{/3'ow�H��@ܑ�����#]�*kٲp���CRme�1��K�� C�h�c�T�i ���:�M}h@�2�0��a���IV���;H��@����y��׋^���@��Tyg�� �̜c���.LlO�0Y"�"��_'`:AG�	Ff�X	+(s����$�/8O;��t%�
�6){�:Ai"����Q&s��oAՋD���6�<��R-�y>l�R]�_�*�x6��D�<Y�!&��擊�1`�q��F��#0V�Q��O��JGY�5���l)RM�c��g0/��R�>��{j�E�?h��@;B�<�G\��b<Q�3~BK�(��V�̰8G�]b
W�|*^p�x�����4b�l�)ۼ|jE��S�w鉀��-�D7���!`g�o0OW� ��N�0�2��#$�ؽ:��P�����r�{�S�P��_��?�k��d�A*��B�o�:A	`?Q�P�Иڙ��A����F~�wf'~
,�M]�细�T]x�pP�Lc���ҵn��ұ���^�C���v�2�>���� 9��1(�j�T��~�������
Z��c_C�Z�c�#��rO�LLV4J��ؔ�_:�g��?�mU��ph~�S&Q��eEg��"%?��k���ÜVkh���3�I�d��ŉ���/�'fO���h��{����x�`m`��=��T/�I�i(�K�0�䯨�-W"QN�rn�h8��[�+�:c�2�te6��Kl����]����������.4L^�Fa��]P+��u^�v��OMdt{%�s��ܼfn���xi S���e�?f��W�e!ы4ϭ%g�
�I�O ������-���ҝ�D���5�&~� p����ǌ�g�=�;5�|7�o	�K���#gP=}-�4����'��}3�m�b�L���u�XIYP�zR�o$��e7�{����t�>���U�\Q�c��6�<��Xz*��_J�[��U!�Њ�Θ6Y�Fm��ȔϠ���yg�	\����5x�H�1�K�R����W���:�a�C��*�c��9 ,*f$a
i�������q	h��=�^P���E��<]s�Dq%Ho~\�6�5ދd֡51W�R�b?�����´EE�+���.�D��j:��[�;zp`\�nu�L�v�{�� /-�k�z�h��N�Gm�7ISpNi�� {ITc�
��I2~'/;1�U�ʢ�2ˣ�kC�6��n��6�X��:
,ߎ�~���9�/��[W���,�̚��;J��n0�<T� �_0�ݣ�z����%���^Y�H��|E龇�U�m��x�d��w�*�hbs�mq��V�����ل$V�|�O#z+Q����[类{��	���'hs	�i�v�x�U�D��p|EL�:�͑��͖B�B�n�9}悂�'dB�O�P��vѤ�h���@yg�
W��zm[o5`�?�op?ęzn���L���*"�Ă�WQt�����'���ȉ1���}7'�(��(���u���\���:��H���w&^�p���/2���:����p�_kۚe��!��œ9�6�׻=6e� G��:C/p�8���3w�N'Ic-�Nuֈ䈻T����sT�P/I�v���G�a^��~ʻ���b����Y<�f�����Pe�:����,�J�O 1��$^"��m���S���d�E�X�l#H�7���q�J��{'|�=M*�t�cG�	Ƴ;R!!��ܩ�X5L�B �~`���2n��Z���|d�6CD�]��PV�X^�o�k�(�o	AӑCpX�e��PR�е�#���eE�,I3"-P��5���];��|�o�B5�A����Եo~�1���2���[�u@���]?8���8�t/L���΃ �]�`;ѰE��(�n��+|#Wi���$�+�����ڙ!�оO-��UK]~��� ��-)@������@�<b�B�$<XI��
�k=�j@�aHL@��D�ͼez�m�����W��>�JW�y�ML��W���J����P�Q�hI�������|W&�t��	/��qU�ɐs}�x�?A�u:^/����|ڛ_� ?m�
�_^%@=�q#7���*��3�[�B�r)��ڙ��22�M�-���x�2DJ]zI�w���͜P
��V���;|��x��#W��h���7��X�'�#������Nnn��57POG+������&�0-������^��&�r憌
��b�h���[7#5��cV�VC!	nO�fe�]"⪼�ol$��g���<߇���U����K/3�#onڥ��$N��oo�byȚ�\L`miP'�ͼ��N+U��>�3"C�6���J�d#T��������ܤ�	ۍ0d� sg��\�;v�@�q�I߷�mL8��:��'�2��_Y�F���^��kO1�� ���F�����a�Y�/�W�~[�z����%��@�%�U��hy�wk�KIbOq��)swE�e�I���q�Z'V��ߏ��B��F�S~�Ɇ�c]n��Hfnc)��`���B��p���4�Cz��4�&9�߳�M)zK#y����BH����������L\}�lj��""�B�x�_5^S���ˆ��d���1�=u��ֶ�H#���I�����P��w\E	/�q�K<I�X9�OF,vZUoϒO�Ί�7ǌo�� ���&|�y'x����H�eCu]��2A���1-3[8�+A�;~���(@�W6�g"o��u�L5<��▩��)p������~��=�;��<�Gd��dCZ��������<��:�^�6��NK���Js�;^ a�͈�b2�B�o�Z\V���E
�KH'?~�%3M�f�C,և��
�J�t���t�q7��[��h\W�-?�L���6ίs��ǁ	�VWѯ��rӑ>�"��� >�P$�8g���f�Cv�������t0n^��Q��C}Vvǿ�>��ei�ddtw���rG�@Z�YfsA|}�P%�`S��T�#�l��(�Z���!�T��̙	FǙ�����a��4���aE�$=ٵ$�[����,�������B:rh!�B�B)U1e��怈�w2*�C2�y��/���_û�JLP���8�y�8~^���j`���ka8k옸��e��0���,;EC�2>��)�0S�MP���p_����r�)Pd]�(��/�%�[�7��|r�X���	��M��dpo9Hi�B2NZake�N�$��T�(��~(`Te���]	&��k��^���68c&T@e�k�u/#�~��{�L%�'B\�$f5�|�����͛J��X�% ���<��q��Z�6Gi^E	��)��I^}����	�?@b�t��'��Wm����P9�d��;�,�Z��m��U,l�7RQ"��Z�)c�"&~̲�U긣h|�gН���6�Xۨ"<�6Nn6?R}.��í��ͯ�3�Y�TA�����`�b�+�P�*�b2��1�˟�ch�nt\0�zk�fY�T��5f��P*��AUO͡&i���Ja�q�9��w��o+�����q3GWXRx��I�m3S[�K�(�?z�D��=J��j�����B��N�-=$1���ܘ?����4�����^����zTɡ�~�'���F�X�6�p3�d�Q���z�Z������ކn�*0=pa-yoI�,vE��q���8�p�p١|9Y�w����E�d:���´�eޓk�=��z㬃G�_w��Nl呴�y����8�Y�&�(��H�G�:@����C�9�\�CK���s.P2�8�.U�+'a�Ղ?$��+���	�����d_qQ�vj@L��B��X���O�"��E�9#ou���J�on��LҶ��~�r۷�r?niq��UKZ�3�g	/�����ď�w�}7�<�لvW�=l��HXZ�Ɵ�e�ڃ�S1��<!nq�/���3���z�B�)����u7�{�� �2��{���C�1�-�\ҜY"��B�/�j��"����t����erl9�xVp3��@�k�Y;��N!�,.G�*�R�w�
R����wa��ݗ�1?z�l_�[�X���!Cap��Kp�D֎�Rȟ������n��I֞�c,2J㿫�V����_��t=�~h�]��}z�Z�W��ywSXWu/0�|#`�e��L�Ã�u���r)Wl�g��6�t��V�{�@�	�h��%�K��cZ2����|�nUf�ݼ3#``�d	�$�*z[X^�t%�T}�a��3Q���4x��jkf�8��p���5�h6힂��y����;�Ԯ<��a���g��H7>毴�Ȯ�4 ���'�mh�N$3��a�>���"���p��H�͉͢Xל�`�ҴO�m��	$D-�d��\~��w��A�l|J�������P�t ��$���͜��K)�X-�ji��E���8�<Ѝ�q��"�î�l�݊ݺa���x΂߯��.!��򳜿�����+n$���X[��OE!K�7�[��#:b6W��"R��l
��o����}��d��=k-:�zo�r��k�K����H���V�lV�k�r�M˜����-�tHy�ܱp�}���)w�4>�W���Kh"���Jb��#A�p�d9��gox�s�ɳa��}�b�bNF�!�S���0�XD
|��]qǑ0=���`�M Ae=ԙP�%�]DC!�o��Sb�
_�M���u96�C��il��kd�M-��Zt��=c�س(�y��7>^	%l���u��-��Zh\��OġB�Jpi
�̹�>�4�M�>w^�RK� ��)8"�����B�c+���.�b��b?SC�*���X*�����c�ѽ/����jl�B������ھ�̱R�����!՞Q���Y�2�E�±����ծʐ{?��A}��~֋̂w��un���5����� �a�ࢳ�͈H:}�z���ݓ�:!]���H�'��j�~XM���y[ ϸ���s�(�ɛ��Y�(��lI�*~���{��"��^��d��ë_A�����$�@��$+�½م�ΰ�"۷�t0���_mlV ;SS^*���I�Y#U�����[1��!��ozD!]�+��� ��W�����f�l\�F���.������dB`޼R��U��[���λ�Tܣ�EE�Ƽ���g��΅����oQ���� y��T7���\O���������0\R���J�)�P�������&x����i�v���hB�X��%u�������W����:�՚gPhr���� �?�[{ě���7���Z!��{�įW�22le��K9�z ���'k�3.;�P_y?�ޥ��6Ի�8}j�g���d��<1�J^Ց���:%c]�<f����(0��֍-v_�̍I]Ν���c��t�F�KU��Lz��}��`-��� �v�W/�
���SI��+g��z�҇O�`*�%?��6h�H���54���	g m�j��sZ�HJK�mŸ�֡p��s"%b򛧎0�.����Y|-Q/�w	v\�O�.�	g�g>��<�͉�$V��x��h��jnh�h��R�e��}y!_ڞ�D�_uB	������P�jG����!5��Ѫ*��
1_����\��߁(��%��1�N~���ےR��}7&��4۷^�>*n
�	j�����'��&��ܲL$t�=i���/|�&H��HE?�����:9Mi��h��>@�;�jT���z������iy��P�3�"nM�(�Dˏl�S��ݹ��d� ��܅���4����Ճz�c��YM"{��
;����e�VB�J�*�'�+��@�G��b�B�%�L:lI�b#��5HL��,��WS}���y�:�7-�����a��e��\|�m�i�K�@�aJ�n�Op�U$�X���6q*���#d'��*n�5tyvb���[i�%�����N5w%��%�z�����Ow+=���I�hC�6� ���1&��	<q
#�m��tj�o����m���7�#w��!Pt|W�6��f�Id�cf�v����8qɥ�f�"��d�K��=ҏ�b��/�l���4ľl+Nn0�25}䇠�3���ҩ������Ê���ج׆�����l�,�/U�+�*n�WG��1h<]!��)�8�&-.z�g�ӚW��M������c��P����C���Eñ�M> R�O�6G,*���3!&mH��h�qN��X�$�`'��2��0:�Ń��+���)��WS��\p��Qá�X��F'�/w*�H��Zn��(��o�(S�vDs$Ɏ��)���7J7;�_��|D���%��+�t5P������u}�&J>0�*S�U�뽛��p���~L�l��|]2�UK
�L�S�� ��7���f!�^����1�ƣ�r���-n�%0��ڈ�fX ���$V�����.�Kۋ39)�"�������e#��D�z�dfI���qjV3y�>��@:y�d��J"g�m�Q�n�TĳV���Ԧ�=�9uV�-�c*q�
��e1���ukk�J���20�iV+�W���W�w���V&��S)I��f�� �^k�
D'ʪr�V3EQ{��)�����*t�$�%�]C�ME�E9��<o��$��E66��y�Q�%Q�C�:a��o�z�]F�Q_��d��1������F�y�)i���Ϫ��sGC�<�'U�6��������Մ`zp�nZ`h�`� �r�Z��"�܂4t��o-T�P���[Y&B@)4P#�pb1��FI����"��W���t�b̑����郄�4�� Hݡ�}�z�Y;Ȩ�6��uJ�a��Py+E^�˴᜕�:���ԭ��̄+
MH!:���F�*tCB2Ǩg��斒�P��ۜW2b!mX붫1]�.i�왺�r��d[xE��p��7�m��c���AH�A���Jt;W�w��������k?�1�-��Q��R�%Z��&�,�����t�t^,�0�����uWN��]���0P�s�l�ak����w���js<&�Va��Ix^�'ć��p@�k�R{����Q����g=�c��z�^�:��q���7���S�'�#���64�wx��V~�!���ؗ��S��aZ���:(?���ޭQ+?��ÞlT䗷/�W��}7<i"����/S�x@C߃!��7���҉2��4#jZ�l��K��h{�Kؠ�=[u���p5(�ٳHb�RPKp��$�B��,n�P�a$)^�Wà��To@�M���#�%$a��Bʢ,|��l{Zܬk1p�}�zz-�c�T NN�|Y;t��jc�W��Vn�h �
���å��.:]E\�	��[�ޒ�e��#k9+!#�'�Y�0�j�3��@b�<�;3�zju���d��dcqx�:C�}ٍ�l~J0��Hހ�m#8⧳�9d���k5C�I�!�J�ߌכO��ʋ�Ó=wIF�u&��'����>W���+É� �!���Nt+D��+R&����|C^�8V� 	�#�"y�G�0�lK!�nfp�����P�g�UX��5g�' 7p��|cFo�?���+tX(ۖ�g�V�r�#U*��g���'yK���Ӯ��u	��Z�Ub�oʛ�c�N��L�E%"�}�D�{�#��1�-�����Q�������w>�Rmu�x�+�d7��#6������Z��УtE+�O��k��kVQ=<2�]�')I}=%K�U�x��go�&%�_,$� t��s��'��2�L��Y`�E97v�FS�8JK�D@9!B�GB��^#ި��L��gw��KSq�|��$�ベ��A\+>��k�MG� �Ó�(���XDvq�]� ��!׼"HI�e�2� ��0۾�yM	�A��7�FCT����,�f�(k&!go���Ӌ��cÁ�ɢ�iWpgؕ�SO��S�yU�:E�5�ǔ��EfO]�l&�� j+ʊ�l���X�O�т��&�f��I�FDv���SK��e�֤�������dRNa-�#�w᫣��ƺ)q,
��dօ�ZFZ%�S��
�)6���g�'��7h�7��L½-��Y���E���O3NM�2r��<�HTq)�$0�u濻١�s4���hQ���x�3�������]���a�,t	K�鱽��,�p|�r9L`�i�wj��e� ����@m)0'�8��crp)��s+>�y6�[�ͨ�{�����J���]�Zj��.���G��?'8�ǂ,b_G�#q�2�mt�e���i� rNM��3;�+�&27ۢ����g�M��L�j�\F&��p2=��a�t�%�%��Q��yd��cp��}�s��s����L�!���Gy�/����/],�[��.%_�7�*1U��-�&R����Z�`�6ȡ�4ܼ�z^�0~d'���XhU��;�a�F���8�N�~H/8��yeZ�L��������C�8��Ȫ���(�5����C���\+��������Ӏ�����h㫟.���p����n<�\s�K	��F
E���e']DԨ����b�8�/'�<���YF���\��$\���7 ��5�[s�:B�l��\�D�����y��x��^���~rw@�	��5�hT����xve}��D��o�����*��b�!�I!�C�y�F�>��|�pT�@���� E]�J�iL���A�udo�BI�e����M8u�{���m�Z9B�O<�ߖ2��J>J�5�����r,"��QV�5����1ԫQ������҂�;�H�%��yI
z�d;s�L,"���b_��E��aAj�1&4���-��!�v��0�X�(���΍�[FVw	<�i�*���������������ͻ~]z�d���ٌ��F=Ť/;vL��z8���`Kf@�s�-np�7.������9�n����k��������D�V^5���,R�I�a$豕f�nYKf����X[%9���Y߶�(����Ka]9."r�w�L��ᶣ�t�q��	Et>aIU
��f�{7l�4.G��C� �����ג���+�4�Z�ck�������$)�ls�"�C}q�?b���|��0�-_��]wq��8�{]��Aw";���)2�7�TMV�yg��ĝ~�&�Ǿ��b\OS��'�m�#+����$9�a�Ψ!.�$)�s��xMO!����3C\.⡑<��=�.�QV�0_�w�S�@����pc?-�޷�j#sd�|%��&�G��#��Ǻ�.�	O�"�ᬬ~��R��$� ;}�;$:v��rǿy�����-��~�
Y~D��D2�k�hH���� �Q��9[�0��H��D�f��1�P���%�cC"4^�� ��V$J���<�˗
�]�P�f��D=Z���l�,�oRs4��CԊ���dw���irl�&�ʷ����?"���U�Mœ ��9T��J��:��� ���
�=�Ȗ�*z�+�d"�Ox>�����燅�sh")���Z�iB$LU#'4���Gz�_�R������s�ͬ�W���	 ���\����|�F��3Wl	q�D�]�LFr�51���C)�ܜŽ�t���$>��I};lU�J�0������놥i����h��n/���a>}>MIK�
�q����K� S� ��@�>���⁋\�����q~�Sj4Ȧ����\�&���ٯy�2��ܐ�l��Y���g�b���¢>~� ;�Q	��Q��g�5�����gyT^ ϝ�;�v��pǛ�F��I%�,<ߺ��΄�/��<�F�784:}Q��k�D0rr��/�����G3��_�Egrƒ�.�l:�Ș����!�J=]�H+� -��AX�tҀ( �a���C�@6&����_��P�6��y���{�����_�Tk�?X�pf��0.����o 	hbXv9�_Nvo*.��������MK���΁׮2At�b��Y�5��~�0A؅ѷ��ZАQ)oșWJܪ'���S\�=�4�D�>���Hw{:�A�$:�L�_7L�v��2kM�_Z�N��. 8��+ȃ�3�i+��1}alᐷ��6Cq_6(��{}�"��n$ST# �ZB�C��q����ͷ�t�m��=?��(0PF�,��&ΞM�Y���gV���IxNǁ�f��,@������F�&���9��- 2��==�3Eu��X�m~w���B{;hTR�G���Y\5��o�t���,�eV����Jـ�y`+���Sⅵ�q2zgn��JB��T�rt8�_�q�m���Bj��j�7���!V�ĳy��2��sN����^�3��-��O���r�l�DA9xgL��"d(����F�q�}T�4��0�/hlj5~�����_�͡3Ԟ�q�d޲��nb۫�	���p�tΡ�%�5x'�Q5 uH��hSn�����ex5#2�[/�����D�0'&^O�S/�����E�C�GMy_���ԏ�߯"��oWw�L�Q-�� ���C��S�F�{�D.����Jfܥ-/A��&�B�-���5r�CƐ5���� �%_���o���O��6�T�R���+'~g�B	P��R?F�Zn0�QdȿO�'�F�ihl�Dl,OZ�ydU��G�I7�nIۦ��U�OP1�tń��.�����w�z�8!�[�3<���i���u}��ac���t�|�8�`cqj���d}9�o�e�H��{2��3\�������?ӣ�d@U?�@W_���eC�s����wt�
��'��YD��[��b7���P��{�]��6/���������W7Z����q���;�5� ��ٜ��R��Q��x��ު�V�+��7�\�)Y��֓M�UU1h����V�i:Sӳ�[�$%�:Q�#�*��@�յ��o
��,�@���jSRS8�
 7����ū�$=�2�;�v��m�z�5B��y�7k��]�%��6#�f��V��2���ۖۯ^e4W�8�w�U���j�69�(����6��j%e���p�Za�y�`N����ʱ��D{bt�x���5�:�b�s�����~5��Y�0�q��g�dI�[Ƴ�;ᕉƌ�RK}R'��.h�m��������2�Й�LT��$�y��L);�g��;��{�޷`���g`����]~���oY��/�k�Uk��=n���˹K�5ۧ���=�A��.�u���X����)���,�I�\p��9E? )W�c ���l}Ё���<�>��������^�]��22�!|�T���`;ʈ�q>I�����ƣ!DXq����Mά����J���;,�l ����L�9?��BF(��1��m��פ�H����!�^#�����.p�T�{α��L?׀c�����;BL)��Y�p+��ˋ* ���<� ���12I]���@0�a����N{���V�B`� J�S�<8��+��9p���S{�߭_0��>�C]��Z�TA����eo�m,�?��v���1��!� |�	�pxG{�""��z>ɍr��^�u��_=���ʸ��0�xy�dAK}V#;��fU�1#�Y߆�<�N�Y����$�j���}���/�+:�0��,��{A��T�C�0]�K��I���{����8��l?x��`qa��A�JcΉ�Qt��[�`ǲ�x���ѮMſ�q4и�8��G%��nf��;��B-��J��oZ|K���E�m������~���+
�F���ʏ����[t̲��(��cץ�5��qz��@�����~g!Y/��^�KB?@Citd9����썑��#�x��mڴ�;(��e��cr����%��u�R�c	�'�^�z����c?|L�v��gr,D�Ęz��<�vU�QU#S.��oL�<����q�gp���-��t6[�e��6hL;�-uB6�4
%���n
��S�Q�M�8!�K�CFM����}*x�ㄹz� O�cY�t�ɇ�#a4�C����鮘���!�[�F7l*�e�Ȓ�u�&Vm)p8,�D+�3��a�ђ��	g��h�'�����m�J��������,@�����VVl"2z��>�#��7�A'�J#�)��$˜C�'�Ss�x�l)�I���yw��$;���G}G@3���Z]t��Tmd�E�o�ȽJ�;��9�7WY�[����A�z@W��ګz��J����,�Xzp����oFn����@��~�7Ś�>e�����̹gg�\���nL:��]n��>!ky�K����~��'hDDd�����_�`Y�a���D�G@a�ܴ�������:�jd�Gl]�<Q概i5Ώ�ؒ����B��@^�j~'2&5}
f�E9gU��$7A�Ц,<�A���Ʀ(43���.�����q�֡�+�;�&�,
K/���3�p�(� �	+e�+�y�5-��d�����-_�#J�^�2�-�88`�u���A�M��L�.<�ۗS�+a
�W���[�%��e���e�
-[�Ħ�{(�K�H4���g��|�66{	n�h�U[졶G�/-��X�B	8x�m�\>�K�Ol�[yq�uX��#��v Gk��_j�1���^h1ټ�XB0�J01�r��9b��h��Ac��[-�Uק9B#��|����^�f���=��M#	(��t���8�
��� o8��gޞ�Z	�>�rԹb���Fj�
��?�Z*��ϐɭ�&����r;�wS�W��B>A�K���G^��J>��<��F�B�����-R��l_�Fs1�T�&�I�Jm$jU��y�$���0P�����(�2���v���Q��RQt����X>��� ��y�K;\�!��l|:^�W*Y���	)���xJ)Ь�C"�u�C�ȃ}��t�V"rޙ�~ZY�4���54~���^tB;8 `'N��6}/QgC-+��s�q�}����Z��:#�3�r����ٯ��s��zڻsN5OJ['��#l��aT��BN0y*�D��bfg���l�s��\ܣ�o�<�Ь�K�X�\�ԟ ��2:͐ż�V�"1�j�(�L�y4�Ů��:4����~d!�ռ8S˸i�bת��Pz冇�saAO���3�e���"�E�y^d]��f����^�u��ү'u���M%E�3�3�8� 8V��d�@����g^��+b����r��Q��2G�	���B��<��lR�Ԏp:jHo�!�>��+�9_���wI��^��F3��C��5ڒL��ན�&VT���K�K\9�T ���/$�[���C�d��0Ua�z�t�:[-��/5ӽ���Z·Jׂ��{�k2l����Y~�_�v\*=�٥J��B�Mi�ݒ1J�p=ev�7��"iBB2�5���%7`��@	�	Sl���Bl��Ԑq�u[~:�?���Ȯr���'��\y�O��b��3N���0� G� pX� �%zw�v��z���|�m�4SL����!�6�M�6���Vi����Q�����0�S,�q�}LkD����U5���_��u��Jk���.�+��w�p�x�C��a$<,}m~fep�8<�%4oo"�HA�6-�����)���#�	5� 1�u���D�S*9F7�j�y�}�cXP����o;��^�gC2U�B� ���|�f�������(�A���3��ޠ	kZO�xY��lY�܍4���
���$�����XC�S�;<������Yǀa>��}_g�4#�&ۃ�l#��P?9��vhY���bS���B��]��B�D������B�{��C�������m����lۙ�EL�ž��j�A����K��um(�8s��b5h�ē:�.���tb�����j�Hh!Y:X��ze{��W���x�F>geT�	q%�
&�D4��������n6N�7р5����c�Ŀ��O|�����t̔A}w��H�1ꄫ�����f'T)_.H��d����|��cV�� �1��EX������Dl��M�b|���;n�Q�'&6W������Uc��}=�[$��������tlY�~�D�-��B�p�pK[�,� (����o�^���YXIt������P,C�r���=�Q���܅��N"��eRnuatd�lx�zW��>�FnDH�k
l�l��u�E��:�9��{f�*��Pҵ���$7^F�j��+�AHZr�T%^�<�اܖ���>�ؖZ/E�y�nbC�x{?%E|�k�1��d@��X��,�=��v���'?������64�Eݖxz�hF�$��3�zn�`2��j(�X��)�!�;��ٓ=Z#��@��?B;%0���䩺)�@�����4c0��l��g��}�-}J-�<��$k��Yk�����<�v�ͦ�B��k���'��Vk��`��o9��u���5o�!��.�Ύ�*��Si�2�o�M}�~j�<������J*um*f���zS{�E��%s�G1�yx���xY?����Gʴ���{�\*��Z����0������(d{�զJ��ռ3O�,�n��0
�^[Q�	��0\}'���W��A�~�n��!>�_}�1u�{I
�Q��r��<����5a�}��g���w�Gxl��|�4Q�L%���_׏�)eӛ��g�;3�q���#�`_/��\��v0�V�	��=i�lڲ�_���֘)!,�|3Ѐ�I�p�wO!N���jZ��y���Zc�U��o�O���1C��H'�P�����hfnu���5����V��N�N�k��W,�Sz
F�L����x6,�����ݚT]sA�o��%I�L|ՙ�rX�C���6�����	��6§���� �q+���l>d$Z��a�M[��}�,������ⲡ�P(�-4~I���c�G����f�"0/&�FF�Boa~y�V7q@$-�6�?U�p�����̜F�fL"�[#)f���pQ�k~[`��<pd�Kџ7_[��f?�����J&C��CD�x����r�o�l  ��Y��u��Z�)?ǐ�	ϖ�C�ѵo��c�U�|�_OR�!�l�?�ܚ���?Sì22��޸�y���&3���l�6�ْTڢ˦[=��'%��@0O�\�/F��(⁮jEm��7�\K�fM�3��Kr��q�n�[4�Ħ�PEA8�MJGz"��7�^G~=�桑8�[�i��n����.�db��GU��`�%�?�mjo,�/��)��"�ڢM'o��'��;�����7�h�[�6I֣vɼ �(�nݩ��~��ZP�k�7�qB�/#�eO��&#O����9JT}���]C0d��>e�������	M󠴂O$K&�Ȋ�{-�wBŌK!���w�׉�b�r����xĜ�i������r_�~�8�����Vb~T+�ˢ�����B��خ� �0�(TP�jT��Y�RǄjM궔��i"
1{NQs�X��} @f�݀�	)��K&�~���5U9܍W�u�h�i��.�O	����"��0�G!��D�C������M�l`���l> �	����������tmuɗQl�����6�B��X�&����.<#7ȱ�~ �~���jї����u��{9�JD�h1 �="'Ы�җ�������t�x�n̗�Aˁ�c1�8�	~h�*���9A])s¨B/���!;��q��p�~�
Q��ު��!!G<Gl�Z͒P������ +�]q���pd~�Wa#_�j����R���vz�ص�����N�!1���W��b�]9y��ܮ�ޓ����_��N`õ��Ӝ���]�mw]�vC&�t�I'�"�!�K?���*�'��T.���\'A�C��~��!Y-�J�04�0��H� "�.~�#c��1g��C:s����F)a ���qS_,����{{f�꽡_����,`��u��||�eoB�S&�U��	�hdS������B)bq�Κ^ͭ���S�$9�X)A�Ψ�Nm�@�b9f��_�e.����x�Y?�m����㭍�v���ҿ�0xgIyO(�pɳ�A��[}��	GQCc�Y9�g���ր�9 WMD~��9�nAk\�󻉨�ugm��`M� ��������h�ٿ}�|�!3�*��� 6��?��|T�y��:���|!��\���о!:�a�+�^�v�Kfb�q)�C-f�Y3� �~A���8�	�xq�lW|�
&�8䕛Cۗ8Y3���w�t^�4E���N�䱇��Jӊ)��ϙiԨ�U2荜���1x��)v�AN��ę�7V��Ki~��$r�Hӈr����0�Lh�p�.�
�{:k~M7\P<�e�y�7�.z6@����2�HM|ѣN����6�L����n��xi�Χ���4��[Ac�-�ip���s���A�t�4/�?kF`❧;����.,Z�kT�9��F����z�%�����1���c[�H�C4$�a���u�6 R�H��mĚ�I&�Ȥ�)�by	�d��Pq�;�$�����-u�����L�9>+�xQ��`:r�4ꖟc?R�g�7
2������`�%1�Nu+E2xT�ꪢ�����|q����~�AW'��-o�?�u��	�9���L�Q*�L�g/`ܤ�՞ ;Ez�*�_����� ��/��<�
�#��t�i���'4P��Km�5���w�.k�,�\�N�0�����a$�7�-�3���s�m)̡6)me���d=��&[[N��Rղя��{e"Xفd�S�^,OZ�w�0R�Ǳ3��\��ތ���n��a�o-��~���v��qV9b]��s^���u��B��#��eb~ ��j�w*͝6ظXڙ�R^���N��|Ogt�V~u��������%S]ɨ2�X+�� � �t�R܂��&�b�%���ԇҍ瑇|�j�A�c�E`�iZ���o������]mђ�>������+��Uy��=�e������<��˼�������T��\�3�g?������)��ݩ>,T���4�t����PS *P�X�	sgVMG�Is�D�V��(��?HgxtQߘ�H���q�V�B[��,��<�9�bC���Ih���$�����;U�݁:��.s=�`>�\�A-))��^"�7��
Ex��w�C)<��( ø@��LW:��>)x�;H�HF��O�`����H�FO��x�R��I�� �-�����C������ϒ܍K��֥k�m(8�(Li�]�R���3���K�kкBH(	�dwy�&{������7 y�i�H<�xT��7��X�z�(D�*�Lz5��i�W��b:6Y���4��d|��l�϶�l6��m��T; ���I�oC�x��;JҐ2F���.a�/��0�!�2e�qO�X%�oS�Y��].함�~�Y��e�N��Had��th�S|��Y�!���_�e��pX~2��֜�K\ط⟕E>;��͛$��'R�>#ʛ�K#�s �󃾁��M�a ��"��	��*L�H�Nf!`���z@�?td�xɏp�h3-��@��d�\q7�������,2"�~�hmT4K��mu�ӫ0zz#un\-P�QU��7z�L�є��L���Z�w�b��B� �L^o[ܝp!$7�%�\?�$���ģS�P�O\4sZ����`bK����^��h����v��@�����Y�wZ O�z�uы|��;�鬭ק1���0�j����M.�u��߆�O���
%��&v'p�$9M��TQqA��������n�v���o�9KF�ZWGG�nS������F�	G�r͎�t;>������#j����d�j9�/Z)��:�̎?;�4#��8>#C��1q�Pc�0ᆉi��4��S�G�-�ϰ��"�>P��L�i��JSP*��&bR�]�ߍn`"�ԛ*�
 دN��K�Ѧ5��c��p�5Ҕ�a�L��8�c�c��o�'��Ձ�@�:�E�����+�lH*
����,�D�F365�9SB�d-�aŷ��c���KK	��%��t+�i�3��I�$;�
�&vܙ��0�\�q
}��V��Z	g��D�+,+�A�8{ՙdf�9Ŗ�"�sj˿ɿ�'m������qB]A��`�!�)͞~Q�d?k��k�B�����VUx^䘸H@�M"��Lot����=��z
AoM���W5�%?lEl���1-��8V�k�� ��#�qg}uP���w��i������ S��D��^n�P�0`��]m�74��$�UY�H�S������Y��Q`[��]�]f{У��s���:>�#�!�aB��H�̩V&-�>x9�����0��o��g]�Ŕ�ٷu�܊�v����@Y� MZ�$1Q�nK�X?��2Re�$]8�%_��<���2D��� rԉ��r��CX��b^����b�%���$��k����Ү欦a�8�$�w�ԯ���'B/��[������uiq�;С�M[��ز����]��k�7_�����*�dY�Iښf&\$��r�oD.
�C�I�IN��41�-�r�*1����c���bI�v�J{V���:�M2ua9J�,�-���G�d����E��s}~������^p5C�:�˫�{8�u�G H���Q�4�������PWr�u1�O��|�1�*8^��!2���B��̖&�0ϛ���S�m�le��`|�[�/+�-�\P���ɰ����'��g�>QMMaő"�&J����ծ��t�tQx7��F��TI�og��*��z�|z{������j��x�,	�ǖeݼ���,�I	����m��H�x>���[��`�#|:0���3�%�Ƽ�!ڟ �G˨GX�,ڸ�E�B0��+� �.�}b@�u�@�a�O�wM�%��h�E/Y&��z�q�f��?9�j�h�͇�����-7%��ɀ)�Iz���<�Ɗ�B���E�mE�O�%����v�*��s���!tM��Af\�0�uK$�ux�|�����'ţٙ��͌��2�������
�5�u0y�r���x����ڌ��|z�6	�������LH�$�C�����4��<�|��4��Rs�ȹ�DYb,��fϻwUO�$�X^����7a-�6P�.�[UȻ��k ��V�~�_-Q��c9JITdW��
�F	o5r�)�Q��n+���vL!�O�J���Sxf��E�Ϝ�N�0!��ztr��9h޿�2�X��wp�v-�C�|)7K�*VV�h�S��CBH�1�@������M´�u��.�S�s�"p��_JϮc��V�$��_����~l��6dJ�N����R*�L�.[B*��g�!ѐR 4��`�����bO
H�����2������ 1@��kE�L�a+����V#�ʷ��t&�9���8���ct�@���|\��Шq�ۿDl��} DJ,U�m���Q��6�Z?�����`A,��N��S�����لUo+�!�IK(����A�I��ز�W��ᗪ� YD������j� V��"Q�A�}"!WI�Q�/Npw��Y[7�5�U-����)`�P A�?��ԻW�ݮF{�E���&�����w��r�McjO!`�#0ٛ�5�ng28��:v����M4 r`ƿ��� �V���2úmo>3�P5��<������� 2M���lJ�ߡ�+YՄ�PI��(5�d��?O��M%�:����%H���/]ȅT�Cy�0�zi_RV��G�����}&�s��]]Ϡ�n�K7$�4vat�~tg+������A��~�W���o���������;z��[p��=�[}�C��$�w���_�ǞK��G��}���2�g*�W%�ϋՂ���j�7��⪩u�ɍʍ�3~m+�K���]�+��]�-�������㲱ҙ���a[��<�^i3�l��j�`�����'ٷȇF`���G���²�����l�F���Z���MDɄ����6�����N���8�h0:#ǩ�P��w.u�at;5t7�������.�J���տ���C V�"t1��֚��7�/�w<�4�����d9�'���3I��`�r��b�6{\��q�-wD�V;��<JȯOR�EV������r��ɨ.�O��*�Q?��qHNJ��!G�ﺭɶƎ�-<��;V�M�"�����C�i�2&�6��m����x4�'��y[��Bp����gFX�$������G�kQ0���Ғ+��E}���5U��5if�]p�D��7�Ҳbm>t�B���Yz���q�ڱ��w�Z�}����뙠��Y�hZ,	!(W�?�wƚ�,��茦>e�����G�ا��?��_t�%�A}����7��`ۛ�yr�c�����UP��m p� MS��.�3���~�]�8��g�ܟ������(��F�1c���tyK�$� �9d�j��BZ�V���QP���l�Z�*෹:�yY��&������[�w��v�.!�!�(+*�tr,l[ը�p�?\jT�&��9Ϣ�O�1�h��,ͪ˻sqU���8H�fPᚊ�Ol�B"(֬�f�(��`'r-G
�����z����-@��c	c��GlN�؆���@1%�#"�����ާ}�: �h��z��E�&�W�������aD�Vd�d���&�~�"�yЊu��s^AI���nޅ���$��f�'y�;ں7sv�<=6�� ��S���\���0|�~�F7cR49@J	��8�L����%� �H���d'�2�������a��vqP1�{�E7W{����R�J�/q Q�oQs�#e�J�R)B���TJg�H�=�*��H���)a4*Gܠ<X$2ls7�;���7Q9]��K��!�`���̴Y�읯�ԲD�'$QGBeKѺ�(�\�+:��W�?�O{-�K��|�
���;d�/*�.�}��E�2�\���I_�R���>M��G�%��	s�EM\��8D�'�k����;H�(]�NHJld��q������?%d��i��&dx����~#���D����>��Ѽ��S16��L��1o�>q=�]���Q���p�0�;YOO��B��Z�B۽�)���u�����<�cRh�/1@�����M&����'XM:1���`�H8�fHC��C�pMp�T�&N°`03�c��a���h�:��L~�"�w LP8�A~3͔�~�V���i�e�]-��¯{Ԛ{��.0E�K�1��L�(���h�D��9��4J�+x����T�߭��J���^�z���#i�,V��0����	�(E��6l
Ǩrk( ��1d�"u8z��!�^�5B'@��՞��a��@"�{�x�����Bu�����s��>���s�G<����B�uȑͮ��W-AR�]�N��cY�E�_�>��h^�!6KƷ��]jQ�g��լl�>���J`"�`( ͽ���3�������vȣ���t�*W����h�ֆ�X߶z�ED�n<�^,�b��BÜ�F��K`ZwBV};�8E6u#A�7\�5QVl	i�����0�+0�r-4'�z�!A]�iM�3a��ɽ�}$ٞ�s%`\<�-�/N+Ampw<�;!8B�RHFu�V��o�ˈ�ɞy�k�s��	P�`gp�����R��+��p* ����������9C\��T<J���]o��~�t<��W�������u��)/i�B{w�;��p[��L�Κ=�a,� c�)���Y�諼'�8-&���1�Q��RZ^�ON�"k��F+��X�����#��:���m_���h�؟1��־�����L�Sީ"���6F�������<[�j����
��<M����%�*�+YӢ���3�ŎC_�ɯ�vI>�}�L}`C9���ڂ�{];j��E^���>��K�{h�ZsV����}��&E�U�60F��y���n���.X!�F�ri�T��N��1)�>+'xMe0	�t ��M'K9 ��*����^���iduϻ����[�ra�H�R���fDWT�iͽq����d;Kd)�FHk��v�ٓ����Q�_ߺ��9�6�TM���,H�0��R���]׋Z]r�6H��]��B�����JZ��iI�;��""֦�~@��ưJ,(u��8�F\��eT�����߲9!���Rt]�y`�Q�F���4QM�;�� arա�gO�Q��R�19�\5�ni�����\�/#\�:|m�p��" 1�k��й��7���]����)�;�*�[��LI��[����q�M���� 󂕧�}Z��p��6;4V��ܘD	�ߤ�������L�Ů!�d��5�4s���ɰWD*��eͺqJ=�1yS�l��*>�����3�G�b��hT����]�:��uǂub*;5D�msc���,f[A 
Vw�����`��r&����O^[K�]	��>-$;�<1%�
�Z�q.�!��%nʘ��=ݥ��6�
���._��Ӏgs ���m!<_���&�O�� h�y�,�/Ϫ����%2�c�k�7�Km�������Yw���6�rOW�	�P\��x$��������2|�6�Ae��\z�*����22L�M�I�N�������z59�W��i%��ǵ�����W�
��^b����n�M�W�C5;��/l�~בU~�f���H���)g*�@�dSK���6��	�{���Vz�m�@\V{H���g�1S����rK�����}��ωy�:��FΟ�XBE�Y�1��Z�/�-� �x�ǀ]o�F�!k�
!#�HY� �K�c�b��vdU�M���#)����~�پ�4kS�'�#�5�-�j�C@UXs��(��ɊL2"4�S2\��'0�G�y���c_P�MZ��EXΌ���0p!V7[��^�泷T�u���ƴ0j���-r�����T��,�i4�|U �c�@*����=]b���~���	} �����@��X�*����oiU>�M�_���T7���+l�o�3���V��:�H��� L�H௡��Ǭ��̟�ҫ譔��8}lg\�k��ω�����3�I���~�K�N�g��$�ܳ+�ge�,n��@��]�f/Lh�I95���B[i��Z�Zܝ��49Ծ`/��([ҩ/b�\�Cy����3�ǲNL�IQ�O�+� p	N��8`�\��V��eF����R��|�q7z�-ð��͕����9i
� �[�2��������2΂�|���^��5�sl�@��d5a>)ى����`b����N�
sH2$���;��4��s��yB%��n������
p3�����Q�����ޛ~ZI��/�;DM<؁y(�rжA试�Wń,b���j��_�L��t��.��jO����:W)\�l�Bj,���0�5C���|�hI�	�]�"Ӧe�W�� �?yc3s>���0}d; 8�*���V�Gm\w���_�8F�W�Z��Ud-D`���|����ji*�j��lU˄N4�(tdq�Xn�l B7�A,p;�:��b(+aY���f$&���Q*�F����J�F��ѥ���̐��I0���<Ǿ���Tw�#�%��\�Y���ۑ�ۢ��¥z���a�bf�v8�;�vY��$w9zj�ⳗ�����lO���ڇ`Ġ�5T�z��e,���.6(�X+=��4h�߷ۂj6��0LC�	�iY]�pє`f�|���կ�"i #��Bɠ?%���	}�U��.��RN���@ԏ9�W[4-M�
6����r�Y�w^�Wt0��´�ђ���IIr&��)3�/|�fY(��=3��0��� ��~gc�o�:p�=1|s4������|�L,��Rq\G�̴�'f	ͳ�XJ��F�:�
�ۺ�oZ}�"�H�/��Pï�K)��7e�k4�.�G����7��U�j������Z�&U��.���I��It���{�j�J�`��h'�p� `��<�+� _�wy-�}�#�>�$q~ʯ�3ՂI,��Z��;� ��S����[Gd�����)e��k�aY4�hxp3Y�}�u��'Xv���3�cpg��i-N�I	�GΡ��Q�����g�Q��	�Zݾ�57+[�.ni�U~�ݽ��^��Ƶ`�iß4M1��uN
T�4oH�w�d��L��t��J� ��$!e�XF�����Y�[xS���s;�~1�EYf���ڞz�S���H�,�;�9�d �a�p��N��E��������oM3g�<�O�A�ޡ|*�K�\JB�F&LRh]ڛ����hR

ƶ�P+�6 �������7H�ҳ֭�)8�=�%��%Bz^w��R�W��n�����d�����{~�� Xߊ˝��W'�2Z�:�lǜ��:��<�H�ns�s��~r���ݓHJ�>22L�bUl�1Qh�꽝AlP��Aim��hӊI(S"Ŷ�g��0	���K�NŦ�|��æ���tG�~t���&�����E�#iI�p��1&�';���>x���1���v�$�#�dg��p�5tp�h����"�|$�|��:��j;f��IB��w��x���;N=+�.�y��g�^y�G�>����9��ۃ�; �ƷCJQ ���؋#zɈ����r�C+���l�f�)��s�R	�Sv�<��:δ0ض"���k+,�N�N�h�ƾjoT�-:��k��[�q H���ۊ���!����gH�W�$�K[a�
)
V���u��b��#}�޽i������^T��K�y�=1�'���$6Ȩ�3qY�T���3�ϻb�j)�8F�w�E�I�����h�F3��-V��t~����\�_�Y����[n�n��"�Z���\���'c��#�6p���hȯ2<F?y�[�iF���1>�de'~b��? �7�=5NNl�4��~+�r���UGwfLA�����U�Q�ԅQQ#�F��q?ZD�o� �b0W��'9i�}��X��Nľ�%���ɉ��~���NX����i��l�/m1.�Ǘt��@�.6���R�8��}��Q����m������Fu�F�������Pc�T�|�aj.<�G����v�Ig�߶
�J믧&ݦ8��&�$Ă�qV��vЭ}>���\K���`Ȫ�Ԉ@b�3�� DҼP5�=љ&Sy�hpx۞3U��>Bʏ�~js�+o� #��Z��<��"|w��1A���7޷��5r����j �j�i,�1彪ʤ�Y>�B��c����_F&�-�K�0���{&�I0��?��yq�6�F���RA���S����N����8�/Z��Z?mܱ������˨i����rՇp �����|�jӄ)��3����~�(��jñ�"B}ߥ��m�z��f��z�vz���-��{���U"pp�ҩS1��j\/*i��(�}u��"�$ǥ�r;��?'ӴxW��� �c\{�wz}�����.��.�r.̣�4�-�s#J��__
��^�$>|,#�pD���8�LYJ�]u-�*qjV<��հԆD�/d�;��M���`��>K%Y�F[��s0���� �{��� �R��y�)�`��<~ s<��3X8�te�L_�%�>	Q}�*xK5?j��N�Ʌ�0"IY�PBt���*v�O�A�.�<z�5N��>����A���;���:c����8E�%�o�I����Ϊ��ʛ�(��O��@�i�&���d�%[�ֻ	=��Õ�3uS�L
Y	j��%Θ���o�;�u�K}����D���Ke�ˬ���W9�G��v$g�h��)0t$�0���L����u�l7�V�}��T�WZ��G�H_�=�~�ih������L���S��CE�8�0\`��&�|R9
��ʛCؙ���o,؇�o����֑����/[��Ց��4�R�]�H��vvL`F�dt\RҘ�/�r�A��;��c�X�����ᒧq^Q���a��ڇ�/VQĥr�N�.h�\1�%1e��w����3}�o��W�˪�?W#�W8
Wӳxj���I ���=��Zÿ����uz�"���l4�}.�z��h^"�y@�����𥽅ӄ�c������"�x2�&X�����E��q�A�<�wW4�������-t�i��0���<�����)�-hN�>M�>�?�F�%�R	a�I�1&~�f(3pW�;؍��?c��@�Ia��%E�I�xjӢmK����qo���?<YS��Y@��j�Ƥ�Ý��Y��g-{ji�_��#�"8���`C�"](J�aA��áO|�v�9H@��Q0�,����K�����澛�J$	�o~jB��I��4(3U�������k�h�&(\}:���i���Q��s�����`� �^Q#e��t����?n����9���c��a�y�f�0I���?p7.<�1����ޢ�J*{%�$��^ث�͈#��#=2�I���n~�i�m#�ؚ��{�������!z�PP�桷�Q� �z�KL&nH|]*�1��r�3>N��|���~b�����m0�e�����L��+Ɲ0S�}��v���y]�u�|�@B�k�]��k��\3�O
��ˑ7���!;�'�wf1?�eK�\�������^r]g)�b�'d+^�mz�{021��"4ĥ�C=XЁ�Ze��~K�.;���|VՏƈ���)}���IB��H�n,u����It������n|�V�X���j}M���ϱ��b�fk+d��"�D#+J�g O�"����kV��|�`�z���������d���c��Bb���xηuĿ���P�	Q���=�A#�jHD�E��,����n���ERO���F�ԨE�F���7	,j�p֚�3�/�nY5���e�S�Y�w/tLZ��L���B��8Ё�O�!fP����k��o�ҽ���b�c�b��e � �F��/������f�+���\��*�Aq�:��Z�s���ͼ��p�'��ϗ��(AA������wB"kL�v&t��6]9���kt*��􍋧�����尊�A3�jV�<>R��E�J�)N�&�!���[z�
8�B9k�Q_|ٔpo�:@6X�U�i�niQ��D�HV.O�!�!z�'��������p���-�rg�C|���G����`�N	W��E���R���Y��U{|�S�ŗ*�yF姶qu�ÿ7�6�9�k���oh�(��nur��(W=������7G ��X!]��.���� K�A�����O`�[���&�7�����̎�=l�8=��P�-�s9�ȼ�(�)2�E��S�_����H�Y���]���<ĩ���W��VlDد�ض^_?�!�	��֐3@#H{G�@9���(���t�1�ڟ1ٱ��kJn!\k��A�h��ϗ�xj�,-+�^�8�=��%Z��_#WB��v�c�?8�L�UﳐyLج���\&Bٖr��1f�Ի:Ix���������s��%b������r	l���8����ݨ	'v#-�Z�0����;Db3���Ѥ ��^��\+4��<���'�.2m��7�;�t�1���M|GM��l[��J��+E�:r����)���m�[���ss#xB���ˉ�	��V�>�eڀ��&{G��m�s�E�A���EA���k�_��-):+��n��j��(�x0���*����3����V1�_^/q3�
��1�K�Z5�ܔ>$@�?�Ëo%��p��9�����	����dpG{�?�1R��C�3���b�����>�C��(Н�����b�R�?���x�W�bd!�⫦�Ja������(kv�V� ��궗��B�9sM����p��\5�6t��nU(�V�)[4�D�;T�rRM��a(^Œ���ݩB.}I`�2�g����M��J�H��@f����-�l�#6�1�E�<� 
�,b�ͭu���^b��M;򇝋I��Ԉ9����!!�R�]V
H#�[KVH��%�2���N������\���q4>!��i7"$4(����|�c�rm�2�����fJ�kY�2��m��rc�KG�	�VQ~T���9�]�~��5��b������!���;J���� -eH)ھ����Y�7�-s�`Z�H��tOx���cV�$d�z�ak$a�$HUd��>$㺂�4��`dC�r��%W���G���8Y+�Ggk#��a��=�}3=�O�)�g�T�V����0L^]V�R�4@�A�H� M�F�A����Ii�]�aR(u���o�u���N�V��9Q堫�8�ԗ>�p�z�)]���]�3d!�c5��s��S��7dn��������g��U|[�Z��z�I�� 3Ԍ�T?s_4~L��\J��,���8-�i�����)����&��s�j���BV�˨:��V���/
�(wr�d�0:Lp&�����~ZT�N7����t���B7��o������^\��_��m0C������Z�U��tV�����Wq��G��tb�p{^cO�&~��ىe�1�}�q'���3��h6p7�/����.sx��ҷ��\W<��}n�K��']ڮ�Ｋdw��.@u�KR�Z��kA�6_\��D�:�Lp�^�ufkfϽ�'g�B������[�l�+�!���L`Q5&�JhM��澉�1�!��E
��򏼫���>	IJP�޷ıIml���u��Oӹ:ܴ?K8��$K��n+��w�L�T5d��S4�`w�1��D&�;�=�Xt.�Qw�B�~gS�,�nہ��?�Jq�t_
�:#ٿՍ�#8Z�/����Qߋ:r��}��_uC]H�C�ǭY�(�.�!��X8-���ap�����'�s}�2�$�-k��.��\���ؖ�*��4׮�oU�\jW	����zϼ7\r>G�M���(��k��b���|{�JN��"A=@K�&
{2s��4d:<�1�_�F'&�2/*:���|�{9vHQ�J("�L�UB%.���Ne���WC�k�M����_�m����\n���aH�ڄ�9)���Ú0��=�Dp�B�Ⱦ�jb���;�����~՟�����1�_�x<)�D�%*qXU�Տ�B�Uvډ�+޺O�ܜ���"��-��z&���5�҆;��Iz"A�K1�N�*k�T\C�`ʬ
:x��<�1i����u�*�p���e�`s��뾇a�_��y�f??
a����f�r�&�`=�߼���ɍd(����^�����T�]D