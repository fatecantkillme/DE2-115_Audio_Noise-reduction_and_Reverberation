��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,��.��̡�+P�FuX��d-��N��$%�I߽7>wN����u�]��j��ܹ�Ucל�|�=í[~��k�5�P�ؐ��T�5�����#�p"&�l�z�Fr&b6��,���Fԟ�Z�_�X�;���93	�����Ǘ�M�~���٘�2�c�D��������f� 3łߥ:ա�;kv��ތ(�}��r�{|�Z�LP�����!�Y{������I��܊7Է^f�L5�:�	�͎������W&��b��wD���Jݎ�IK��et��1���Lt�:��6�Ui�;F�o��!b��\#�Z��k!�Y�#Ao��U.H����Ƈ'U������0JN�]�[�萙��5��!M���@gb�t2�-�!�&���%9$K��:��\\_4y���I��^Y��za��jLE���Kԗ��i�h�	��E�3`���1�!?��rh���-C8q5u�:�Ng� ����l��uwY�����	 �ѕyO�6蔋 '�^8W9A��}�VR汷�8L�LM��0,ǌ�Nb��'��5�.Ր�������}"iGI��M�~�ί�w��A�w���!������
I}yh���DB��h���Q�����/���d�Tj`E���Ĝ+����S}��"sbw�[b�p�16E2�Z��-�3��9����������Ѥȣ�_�5�88��H|�BI�:�Z���ae^�(�H�gdT=1��t�+��XI��#�Yo�vr���pW+{��z�����S�/�F�hY�Ӌf�W愡��|��.��$��]C7E���J�H`ͨ�p�9eS��Y�66ǡ軩p ���.��'Q�x꿹�?3§�	��!�vֳq���{�:�&�$��Q�rH���ܢغ�o#A&�;r��;�;�^�\\�Z'��xv)W6��DaP�{��s�ˮ(<�D�Ns7��ؕ�wA�s ��Y��/[Z��i�#�x&�=�0Ki�O3�;a���&"�G0��.eꖱ�*�^��.�cF�����Y��sw�i�6�s��\��mU>(	��0r_u��yX���a\S(}��9T��Ac�,��r"�U��)�����~!۟O�ɧFXS�; �_�vr���ۈr0*�,��f2iK�W����$� =���ihJ��5�ҋo�O?8��b��H�G�/�݂���h8�;�m.N�O��l��m���~�($XL��tp6�1ݶ�����B���*����f�5�mJV�KW��K��3�RÛ��K��S�!C��U��Q?b�^�C�����A\�Q�/�PaM�Yw��g�2�K/���bč���Ǡ�@�Ӆ���);!�����)��7:$O�+ȋ��D<+�1{K���4�j z+ 	+?t�"��h��Pf�Z����/�k����Qn�fecs�������f��}��.�|,��;�1A*�-`�ʍ������g��C<gql�Ĉ�__��%��.�[vY%kyd-��~?F��g��}��ٳ�0������9e��	}[��rv��1N�SH��6�!��:k�����lƽm�y�S��UA%��}�	�<I\�^g6oc��Bf7� Lj�Y"S�S�i���j�{	��*��B���xi|Ngٓl���h��D�%M��9Ĩ���x�0gh�/���~Er(bi�y�I��ݠq�*�j��P�٩&���!l}pR�
�Nd"m���`�u��q�z����	#ft�`�j�e�1�彘B�a�����f4��"�FhH�&�(ٷ���+o0��f�:9��y�y�@� lII�ߣ��H���"�Ꮰ=���H_��%;�\_x�LY;���D�f� �To���T�^�l�af��q�D���,G?��h�ʳE_�*"u���Eթ�/����po�_�x&�d��0K���j��G��['5�0F�����Hz�续�1�W�/��՗.ʑ��dOq��DH2��z�]�X;�k��=�����ōs�.�μ�l����<�57�O ^�e�l��UF>,I�X�FU���A�RM�p'9��3'���6B7��R:6c������z�X�B]�%e�h�����	ۨ�Q�vdT+Q�$8@#��������_t�A��`P���S\Gq(y�
<�^��֩����P��_��B�Q`Pܮߡ��m��miq��dX�?�֟`G��@s|�G`���`�����Z=A��ڲz�h�9v6Įi���DLM��I����e~�\��<���	��(*�Jp�� R�N����y��TQ)�wf���������"u ����M���b��0ڭ �
�����^�}��e�#~�=�����W��O���	G@f�P���p�L�^X^�Y����a�QӐ����TY��u�)��y-�!Tc~�钚��o��L�o����$���b�A���B���g�Q��؏R�s{C#gV�̖��7#���k]�B�$���t�i��Y�_��<��Ο��bXO