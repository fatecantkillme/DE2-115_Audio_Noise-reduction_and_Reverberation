��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>hs�*�U��Q�����vXH���p�+ׁ4/3��T�?#�ھ�ь�RT����u�Y�����/�Ti�歀R�O��5��s��
�rOK%t�R�QT�� �>���Pr�
������:h�����"��I���*�P�ne��M�O�	r@�/0�,/���/�NcaʘՄ-�a
�lm`��ܟ+T׎�+���Y4��`�����8[�R���A�V8gQ�����@�!]ch�C>s*�v�&.�?��6�=@���I=���hs a����b��%U���,&�U��s�y�ʦv>MF�*V9�:�n#�#����� ��TPN�,7���������Ա�Ћ��)����x#��.�jp)=Z���5�v)�����j��{ܣ��e6�6�9���j�43�%ƪ�����vش��+�V��R�֎*wmP�K�p�r���b������%#N�(O�j�Bl��tWD�e�uw;�s�/w�d"���&*��~��q�"�����z٭'�fp�߸�x6���S<���(p������֣ ���{DN�p=By�;%:<j��K�;oϿ`�k�����F��aV��n��(���ԠL6�	u�pN"J�n|��:g��?�\h�B:��8óڨf�{d%�� ��դ),�m*I�����[r:$�X
`��N�.'fue�]�g}�~�8́C���D{_�$��CG�����v����"�I�Ogy�km� &�:�^��![?�g�M�m��2��A�|���6��vGS5���Q�f[]���2|BH��q���ux�D��{cj��%�G*���ϊ�%ݠ����y7�������e�:C�N�gY᦯m���'V�@�sޠ�tP�̈�g, �6 �Ά��D�?b�>��������ʅ�s�~&|ü:���6gӎ�!�k��Y�@-��)$M�q0�aAK���+��ޫ,�E����Y/KL���c����;0\$��9��(ݣцj�"!N)nV�3pH�(e������H�D?�}Jh�B�a']�`lFæWy��ȅ��)hꡊ̔�KVOp~֎_��
�ʴ��߷��չW���^t��)\�{h�@c����k`�.�Lfԯ�?�����^p��My�Xw�囩Y}����?���c��WδN���-�.�W���H�cr]��R�$��'� �i��v2��6ٵoA���`�@[�qFa��d���B+����^/����Z'�r$P����ݰ�#�?>}��D��ƅ�G���� 4�����"�C��Lߣ��HDs�u���Ias/
��i��uD���kbi���J݋W�ڐ���ߘ�)��ǔ��OB����Ge��T��y���`dw擤Fx��Qܘ-���i��sD���A��L�q�N��Z�ϪUC���۹�^9�� N�v͏Nj�*a�R�{̯p�6�R*�WN���x�`�x���:�E�j_h|�׭���\���vSdx�/�����+@�8�d���������g���Wΐ���⚪������O����ޞ�.0)�~m��x9����xb#��tG�3������+|�I(-:��;ܥX'�p�]WA���IZY�~]�"�����ݲx?����|`��]���*8�k���z�=�y8	!Y<��J�.������P!M�����)i"�?6��U\j���ߏ�2p��]L��<JC�1?��;��֡Q��fRƉ�lD#.m����S_�b��>���j��x���R� '�H+'��V��� =H;4]	��g�W���D��n1�N�U����4	��
bXMQ	��Fĭ�]��X jlο��P�	����,Ն]9G�{���h	|"��8?!P{GF����ըt�pἱ���,>/�YLb)��ب��h*6�je�]�k�zǲ�������Ҋ~�7=zI�@=P��J��{�꣔aS"џ#�%�����c�$4`�q	!'� ���?��94;�_���s,=U��̺y%{�X�ǟ�I6�a�\mπ{:�x�梧�ӯ^�|�^~v6������73O�o/�'��î� ����@�~p*��h�ML�X�oU����>��*i�t��3=Ǧ����^
^�]ͪ��m���ݢ�9 l}�ٖ��R>�W�r���h�1�x!(��1#���\1z�����*�V-�Hm��f~��U[�����,��ca��W��$���< ��q�@U��X0^��ޞ{zV�p5��Y�4X�8��g�	�$��>J��W��V9�x;��7;�]OcA�nR>}e����������}s�+���"(ucH,����|%����Չ�H������Tڄ�0ؒ	��>��Xzs���-u�ȷ�.�����t�v5<R(��dN���#�;�R�ϙS�F�+��E�f���G?u�@C+������z��q�D��y�-�.B���&�Nо#��b��x�D��J�顿����H�G+��C��!)仵6�~�Q�`���b���ɳ�J��R���qLM��Y.ט�?������'�ڂ�y�?ߖ������-�Y��!��{�����wU�K�LO�*P�gZ�����z�Y:��,e�C�!��X�Ċ���_���"���������;U��e2��&�-��W��۔S�k�"�ԷG����_�D�π�'�q1���˝�LT�����lA��3_-���U����29ʡ����i�Iyٳ�������TTC۾Kb#(/vط�IH�������s�%��s���f<K����N0_�좨$TY[�몯t��ATv}�%����y`�^֫T�2?T��̶-U�>LC�Q�oW����*���5M����#x�� �'�#�}��~NB�x���}[�'ah�dc?k^R7k�P|L"Ҡ�cG8���.
�F��\{�D�>U�V��}rE\���2�%+�%��5t��ZN����Ӹ��v�Ks3]�xYM᫭xZaJ��px[�(udh�q���a���ܧ0&Ȭks/!s�4B�Og�~�[^~j3���i*�6e��;���Y���{/�m��V�i�Y�R��T9d~�G>д��9� N�Ӆ�D
�����j5˳;z��jC"�����k]a1܀�9i|�ۙX��K^���ӻ�O��w.t�져>'����>�z߮�`��nI�ɝ��A�9 �^;A�-�a�O1�ޗs3h:|}~�Oa��	!�+�Vҝ�P�Ec�̝wܼ��sv�__���O-]�A����،�$�c����g�ߠ׉EZ�'+�3@5W���ʼ�M<�H���_�þȋ�[��e��Qd�C���g�w��#s�Jk_�oW֕��޸
(������a��:շ¶D�=	L��rB>�+`���{�G��M;�eh�[S�p��_�*��F��������s!=��uc#'�@#f��FU��h�(;&`R��n��
�42��ʆJ��l���FL��_�,|N��f�r2�d���~t?���g���%ߏo��Fy[�x\4
���\�d4��駵Q�pK�1jp���J�����3w(�5���g����c��ǔ�<��Ag"<=���ܔd/{a+�(N��Ē�x\٤��=��ܡ���)�rLu&)��b���s��RF�>�:�B>d[�t$=�䊐�݌�7���J�x��� �R^�V�!6�u��+f��B��� B�Я��艼�שe�L�g���M�^���[�]ȿ�����
�(��E�N�����Q����bm�3>F�ٶ3�{�; �T�%���h�?�d�n']�i�'�Ls2����ߝ�s�C54�"��Bk毀���J21��R�o�G���D*˜R"��F�C]3G4 2*��7>(�M�����3}��d��i�&4�%Ǉ
�$���9�v�urj��^��1Q��b�[W}��C�I�,څ��-d1;i\#�fW:�����9�<I���4}�vb�?o�� w���;��V��m"Q8NwI�o纆F�ϖ�����9[�PV�B<�Y�	 ���ps-�^z}�cW�o��-�bO<�<B-Ox�Zm��U �%�،4щ7심[L����S,�C�k�A�:���8.�@��W���MV��r��t�a�c��dSej���jt#&�;���C��}� ּh�m&Ebf��u�g��Ҍ�,�[�*��͈�ܵ����%}����ǀ��������xE_�)6����{T5�!���b��q҅.J�_]����V�_��f�nd��s4Ф�w�+a�H^�����b���7n⒂%$�\�yI��}���G��M��
�b�?��NVJ#_�˻u��l��.(�� ���(v{�t$S�Y)�☻�&�E4C�˼6�1T���T�WOhA�M`�ο�>h�4n��fY����u�z�� H�Z��������m�޻���>���^�Ꮜ�TM�1�4���K�Tl�v01�&���^_�$$j����@0���z`����]e)�w*�)
�ǮgǿAU�5��'��99��jzṯ�<C��޲���(�y����{�5�)� ���M�hI��C��ka���GL��瘶Y^#�T� oiP�b���Z58���O(7�`��V�x#/‸����vh�q�_"����inʛ�����)"/�d0!�	L�H�J�H ���qmc`|�C��R0��L����J �q�Cߪ<eC96��x��d.Αl~��1"�-��2(0kR{��l|�ߋ��+���3={r 3�K��W�<�]�;l�?7�Q�ǚ#���oM�t��+���E���/ۙ,��Z���?BPQ��@�����8I��^1Y��lp4o�u�Uu��.yh��r�h_L�;�Ջҏl��-!J����Q���7�C�d�s�AX��[�����Z�Fm'��8��V���F��Z���#Z�[{-*Is�z6u 9kh����^<8��	s��%[!^7���o��ᦀ�z��#
�� ���3X�[�=h�$5H�W^p�U�S�k�/�� ��s��Pڧ��p��ҷ=(~>���t��MV1Ͷ��v�7f�sٿ0u�V��h��N�iC��^��z���`���CS��X
���rSS�E�y�ۙR��˼�-�PɶYuv7��Mu���Yir�Źi?a0���N7	���J��SOz�����Ka����~�a�	����[�?,���)��,��������2���V;��*t*V��Oz �}��iB�[���,�nX��/DK-\���3D�����!W�'7�J�@Tt3^q�0z�xP��-�Z�v0��ЍAK���̉�/J~�>c�X������<"�r�0�TQ�oC������k���?1Ad�@��
��1����+?�8G���>� aW�֐�l�R�2[n=�f4I�m�x Mk���|7oP�D]�a�!i��o�m�~�}��~�iSzftoME5Y��$
���
 ��3Z��fh[�)�FN�J4Y�y'��)�k�-�X}e����a���"�F?"|���# A�l�̳J�/ҿ]FU�ZQF��6��ְ��\�2���Ͽײ�@�13&8b(�-a٬�g�dH��8X��#��@N1�<�g��k�)��*�a,'�~KQ!�j�Q<w����ؗ��IG+� �R�/w-�O9��J��3i�ҽcy�A@���}����pU��j�4�2"���@��(H����O�*��A��{�v�O�ٙt���o�}�M
y{�$z{� ZG�G��S�[���7�a�N��\S�.��8��������2MJ4�K� ����}���_4$r�Ad�ٚ1�r��*�g��N���'$ԫgc��z��ȹ�R����+�go��bָ�ʭ��?�
��1���bTt���l~�X�����Nu�fgT�����7$-����A�́�ˊ�J���Q����.h��骷:�}�{��W��웢�Q�T�x�ƙ2�<v�t;�Fx�s������*ђ���K�-�ؾ���f[[�}YQ=�4��H�sQ���;	��,8{���O���+�i�I��k�҈Q���M��{+0K�)���~tb��pyn4� �DF�m�]��`�S��N�i�s�5�����j����&;�5�Kb��Z���������GhƄ|O�̍[aV2��@ӆ��6��tR�ۇ˳��d����tB<
3ں���V�c g�%2����7G�*W�����+ruc��Y���+<�H��oy�!?�T{ZKk�3��Z�����I�;=I�x�gs���Ƅ1N��w��O�d�hx��2�o��S�o�T(͡~s�y&��
h��Plp����N)l��|�� 8OڝZA�˒�n�Sd*z�{[-�EK�8œ��H,O�l� Nvfh��Q����~��;��iWBS�sT0�ix�%���>3�ƚ�L�Gg[*����F�Yʴ��}�ۄ⃀��c�J�Qh��lP�����K���<�y�J\��X s�#uE���F!@|k+�𳃍�p�j}����7Aq�|t ߑ���W^Y��$��=�b���*���[�Sn\I
��6���|$`[\��b��"�?�:�}>�Q;�6vsс�E�vέKŠ���fa�t�~���Ho	���\R�q2Nb�AWbt�6tI��&j��{|{�I+�}�	��"�����lK� �U-���K�|��f_~c���ɉ$9Q�2P^�p���n���RQ�k2]G(/je��^F����&��V>�]x`�Q�@0�k�1�ɲ�t8�k�^9�5�A����(�q'4�Msؐ��m9l�{s�2���_�r ʡL`�����`��cZ(�6'I�~��o"��C�ͭ���ZuK�Z��'�
5����K�(�����e��5(�H�>��"p��e��2SUy`?�ʞ�#���u��/O�%�z��z|�1P���+����T�jxo���&FFTG\�NN4�ߏ��8�y�������8kC�ҍ�GB�O>�ꏪݳu����k��DC�΢����P*�-䭃n��M��F�_.u�e���i�a-�T�uU��H�� ��%NJ�C�M�S�>����,?1��Xf�v��N~cG��;�a>���)RY�O��&�y�Z&�p�����Jړ��!Vd�d��SHڔFI�%�*,�`�p�̷WhŽ^��'��}���^|d��Y>���ק7�-����8�C���}���X~`���]^r;��a=w6m�G�R��\�<�������L`��K�bu,I1���**vo����I؝�@p��vC���(���!�O{� �T����^䚑�_�R�jW�[EI���L��Κs3C��m�tH��Bo�V,��Q�b�a�3��1�A&�ˑ1���mH9�n�}@KL^W2K
����#�9�C��T���v!��.�i
_o
��fi(!֦���E$���;
�$���������1��M�Q��~��$�s�
��d� <হ0G��t��R3&��*�%Ieh���Ef=>�\�����9tt�ZO���`^���N��mP�~\����P���J�R]XDl�x3��H�
ْ�f�@���䞣����