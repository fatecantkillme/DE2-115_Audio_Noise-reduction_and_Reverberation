��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>�m��`K����٥J��5ƨ"���Ur�
x����.6P��E¡���Y��ا�o�j�T����� 7%�gE�V�}�eZB@�'��ӹ`��˟���aO�EѸ��^��PMR$�?�QH{�o���KW.��0n2	BE�\5�J��K�8В����N����?�-��zs�����Q0�7u���c��j*(l�Ej�ܪ�v�:N��])��O�jk����^˔���)b��*L�$G3�"�+�i��̏S�����Z����_bn͕u �?��^���a��T�|�Ӻ׍�Q�P2��=r�e����;B���XF��/k
IeC��![L�D�hKM��Eǘ� ��hP��SL|���Zl��z���m�E�Z�����a�t&	�ܫ��M�+��9�.�������s,a�7�g{E�Q~`�u��P��ѝ�M
�W&.h�1G���zS����	���x���g��j ���/�1J�H�to�����8䧓&�[v�և�#:Ig��E���^�Q鈥����}�N#z�'5b�W���Ʊ�h �t ��(�*��zʰ㱲"�a�����6Yb&�i�7���"�&�5y�ف��zl�s��)F��O@�?R�`�FA�f&�{���,^���`�ܙt ��="�O�93k?�e�`�ƝʡaH����[0����ǣg(FJE�f1��\��DD���#P��2��՚��vK���������j߾�`R��۰�%�$O�����E���vU�-Rk��8I/�,^�=�#�^���}p��<q�������UdݥV�4���g��57�f��� �*�"��N%b�YdP�x�bw���m]}p�{rD�T�l�)=�I�fWĠ�{vb��V����rǱ��7���W�UP#�,,�����[� ����̘�ͬ�@E$�����G����W8�>?���OҺ���
FrnVK�\X�q�wD��{�5?�Q����]�J�� �v'�JO��Ae���\�Y��������W�7J�Z�.OE��: ����W����5M9���>'��q�d3�������<��o�%p��嗀��M�&�$�Q���~�_�����1R�Tb����[	,�g��H�}G��b��[�����$?m����P�.��Ip����+5��6�!��S� ��yl��J��������'�XY�Ig-6:�+Lr���6[�X5>��2��ų�|��K��������Z]�\1��\��^�q&�%����bX>�m3D��+q�v�+�A ��,Y� �a�z�a��+�u�����R���P�!�r<˰o5��}�u	�Ҋ�U�L{<L�d���\Q�jG��zn�F'���-��*�gd��pe���j�c7�N�ìwŝp���E��1B�yЂ�`�}|�V���x�|��WS��!A�z����!R�7Z�j����'T�3jǑ�v���� p����M��ܰ1�:�~*���E�ۏ�?�Y�f_��˸&J��n�/q��u���15�%K��ZJ�s@�� �L>;�b~�џ��0��m�:�#Mi�eQ/Vm/�X먐����U���~��5@U����=�������^�ֱ�^��{o���;㻟jN3��G���3u�+f�q|f9Ӄ��<�_N�6MoQ�!?�.-OZ50n�RI4L����8b����V�>{���_����ϰmz�;��/�c\�/l��ANUK/�%ڒD��r$= ���?3�X&ڠ�;�aw��A`|8�
�"�a���q_����>��*��r���ެ��MOr�� g�v5$�U_\���Xж\"�H��"���_� ��o�jk(�<۔op4w:��D�4�E�ܠg�x�x!q:_'"u���/�!��Ar��p�JNk�C\:d�Ľ~�k�u�Ƚ���/Ii̽y��Bw�W<}8��v҈P�}` +�q�/���K�Sh�������{̩�+e����A;�p�2��z�!'�[�1Mf�v��/揾׆��Lm�"l�8�sІ�2��@�i�-�Xq�y�m��ku��D����젠4܎�Dl��K^%*M���x�'%�vW&q:c���u�Z��{`������+� m::���'���\��%M�̹�O��|�� p��<0SR�0K�W&l��0	�ܻ��L�S�O֞���Fg:,�I�=�SY�����D��t����9��t���I��@�S,�!���1���O��is 2X�S`�pmA��,��-�&����)�0��U�@�/۱���x�oҮںӽe��h�X�'E�J�;�6uр��o�'9/5�Jmw��U�
��C��(�G�&�v�o�0 f��.�ysU@��,ukd��I:*$sŇ�8��/ouq��9,S'
��a����^ܪU��C�w-?l�˪�j2�7g�m	|���G��2b��A� ���\���T��p~��	�?}���in��H%� ��ҳ�uT=�w�r�d�3�}n�I/?2l:[HP���A��T_����tZ�,�?�}w��F�{kY��st\����_��K�B��b��~��qc˷-��V�,�0�����TKW�n�a4;�=��u���_�©����w��"3W���.��S[`r%xn�[�'��p/0X/�13��(zk}��7����5M�v�$uBH�������qD�g����n��(i. R�2J��+��&� �!"[E)ǙP�it~����q��o����q�9ϑ�Eʶ���Jo*��< `���:P�����5�a��ɭ@ds�Yy7/�n�Ƹ���%����9z�����V�^K<�.\럴��)�0�_�!m6������ޝkj�}��M��Gnㆿ�]��JԬnu�B�|�i�g��1��Ҁ��mF�/��bKPA�l'�X=����NC\�y�"�>�����P��.�1���������?�>�,Ħ��;��Gr���3��앺[���6����s�#}��Mv�5�zbB��p��`�H��Ca�����d���b��-�l����꟢�Q� i�kujQ�~>å�g�Y�6��H�ߊ�������SJ�ވ�dh��#g�ʭ��X�`�n�#o�"24lNWß��W+��ٞ��U�/�;�'����'��{��e�";KUrP�(Xb��*Kw�#)��lX���`�L�+t���W�^olt'�[B����f�h� ����,��Tҏjx�FMY|u�U6R`s	e�%��=2Ѿ� }�_$�^�e�!�cS�̚/2ԟ~�I��Zh�ŉ��b�MX�����;�<��,�
�}�����l�.u�T�����w�O��sk���jc��s|A�V�@&��G�g4�������ﺹJ�σ�ؑ�?�qf�/����