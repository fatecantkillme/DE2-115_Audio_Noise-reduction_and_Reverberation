��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv �|�
����Tӂ���^�2����+t2v�g�VU�r�H$�\%8/�!8�1���1,c���'���c l	�� ʁ����h���z%����\�?�;�=�6����w͸>/Q'\p�~����|��k﯃�`d�C\br��a��D�z)*�&fV��X�v��H�F���i$�MJDK6$�����a����S���ŋ<jN�q��r	-��?��4��✑�j9č�O�r�_���4�l��`���l�M@7���Xf0�����5�㼬��[f>�Zu�*"C���Q-�`��d��E����Pk���Bb�3B_�����PV���f���l��4?U[D07G^�������7v�2qZE4��R�g�3\ĺ2�H��h=q�2*��*K��1�ԗM�=��JZ��cрw�du�)K<*�ٛf+}<����Tkf��!}�ߙ�"���#q'6�KT�r�%�~��}�`"	�q�'���~4�:Sk�c��,>�{P�w�@�PG��aK��0b�����7g���h ���ˑ�W�U���a������������v�>��\��'�Y�D��u�P@��A�uw��
�b�+�?��*�܅Y�~��;� �ԅ�����:{Շ6j�P	������À�w9G�HY�	��x�޿��72�f�m�,���P#�{4(FJ��Ә���f�M��㛗�?�-7p��,���`��ɽ�GQ�ؖ0�V�й�`��؜��_)a[�)��+r��Mr�ܐ��K~�B�N���j�*|�CS����.��'�KY8J�u�,���/�Pa��n��M��λ��
��!?4*��T!4�2�&G�t����|;.���Yt���2}�k����s����"z��9vTd5"��3#��������uf�y���a��F]��|%z!�7/�'���l4���מN�������ǘ0v��c6���0����n9��-GpC!<�m��5�	��MqXV��a���,�
���w��N�#��rN~߆��!�[n�>��R´������)��9��k�L\ƜC�aj�,<�����2#�]Be�
��y�z�37=(�zI����'ݖn����a*�xp�o���G�Pz:J�l�! ����质]w�}�e\��H%�����Kx¼��ћ|Lq�ӽ�6��1�T���DK��k1�JP>�Za��z@cK���\�I��5UX
�Ze��%K���06E1�'[Vi]WU �j͐~�;0P�l7��	-"7��S.e�2"��c���iLilċ1�C:��i��ހx��t\^�[���2Ш�	6J����c(+:̞��� C%�0͘yuOR��V�5]<�*4��Y����r��I��!��lx��Uԝ3��ޓ�I9|�؆H��+ʘ8��6А`�߸U�6|싘���Y��_ty�K�qdE��	�������}�X�f�<�ǯ<c~���5�y덣����ob˗:�B��
X��P�SOh�b:P���(���QH�}e�k�@�Gs�Nt��a�K&a3�k[�v<�pI9���J�}.4X������y�l�^��EJң���x9�s�����.譝X�6��]q���4�����e �� <{����P#�D�*.��2>�bdI�� yr��m]��� �&�����c^�oZzmw�%���J��
M�s�ڕ6^9��;�� H�a;��	��?'�U�rf������b�\a �3�u|�O�&F�d�58ҁ}�{��͐�{u�dĽ����[�>c���3E��Ŗ��͚w�\_Y&s���gLi昇CI�x!����g���'^RbJpO[�k��欺uz9���mx�zzG�4���m�u������5�C��@��;a�"[�&O��	ūP5�cW	�\����� &�;�%<�bB�,)#�� �!p�~����}d�"k8�:sa���i�}�H���Z���^�������5@�(H6���RS 	�K�>n�N��(�u׊(���TL�� j���3�_���Cy��h#q-��96#R=��4V����O6t�4M�Y�]ĎVQb�����.
u�5��Mt��ϭ�p3.�ư��� ����懀ء� ��F�&2u�h�0�K���Q��v���f�A!��?�uyhC����F���߫�F�"�AM�A�0�H�HU J�glx���sth��NvC�ܑ�?G���mqSJR�3�j���3sj����u��i��ש�}�.-�lZ��h��"�
>l��O�0!@o�t)�\��R"C��<�㹴�������1���T4�^>w����,o�*!W���DċT;B}��%SmK(mr��6M�m��{f�"���O�!���h)�c��[Ж��4���|彞Ț�^T���T�?�l�y�������)F%�cGȸ�ް���Z���i뱏H��1���D�<���]�M-S���1�����{1ђ������/0+�)����}_:�7%�RȢƾ��MB?��Ļ[�16R��P]��"^w<��@B��M��6�������v���C�ݯ�i�KIھ���R?������b�ry�h��T���F-%�Aw�����[+�ohF�ܨ3��Ok�Co5�[�S�90�+���"܊hݾ�=ט^�&�^\��3�`-��zbQz\|��C7J�e	qd�!�����q��*�VՈ�T��S���߇�U��q[�m���/�	C���*M����A0x�������8�ʃ������Y�\�qZd��Q�3d�S�Bx�ܥ�����0Y�W��RlJc�2�����O�a{8�(�$�_o�@�N�T�;D�,�^]��"��1�V�:�er��ǜ���M��M�:��GT��.;���$Zc��'�%I\l��k�@Sd��d,�%گAݱ.�q�~��]�4}�U:�
�YM��
�B0�/�pR�� �Q��:�@�J@��{���Z<E�8��xS.�1�4D�Պ��VR޺J>�P�"��Z#�p2H���9a|��aG%�k;e����f�q���E�-^��B��y�03i���a8����x��2拖J�f��:!��G.����z:�����7̘4�ח&��^��q��B:*h�7���b��&H�1��'�b2%��	��*W�w2~��*L���T=�-{�ud��1����=�q��`5��س��y#0;��P������%�ϵX�>H�k�$�SB�o�V�5{�)�Jhh�VV��
�Q�(�g������5 ���Ppч���ŷ�����j/;�U�n����ѫ�P��*�V�?̐�_�9w�P#jr|ҙYl(�~�H{��#H5iѫh4h�PVR�*��{�ʮ�D�c~<�o����crtN{�UnI��D#��)j�4�#HOV��w����r������I�Bk�4����6��7a���#��qZ?}�"4e�>��؇�ה�죱Ru@>�����W�K������N�eu�ܧ���<qT��]L�i�~�@ �z/TD�$���@W�)WPA�!��r�5�|�q��,D���C���)�,�����:���,�y�K���v@BƟr��جkdY%}[��1F�MB��ow�'iY�y���]HE�dlb�'X.5l*.�A�:���YDct?$"��&X��ӅH�0CFj�Ю~�.H���z�CtE�r1�)yН� D�~���w�&�<�t�:��FuE���y�4�bHx7$+b����a��1�7��V��wC����kB���nu\��1.q��LpK��*]_�Ԟ�mvu�2�%����D-��`a@i��柹A1j"ɺ�6�Ҵ9xϲ�)�e4	���*��C��G�'��c����DTK)ߓ���[�ڧ G@$�_�N����ͭU�1�� ��9"E)�6y��z�2hG_��ɡ�`�@W�Q�}�W8gd��	������=٘�Jg��R�
j>�**O�/uq��ݫ��]3m~M���1xEfS��fԁ�}aSf:i]Jw�8����[�#�`���\��b!t��7��ī�b���)1[����V�u]6?ɞsN�d��@,�vh �!g��/��ҶN��D��&���u���^�[R�H�������j�a�}��=�F�N�[hˏ�#X5��s;y:!��r��T8 =��"A�pU�ZhRU�p�.��I�Ҽ�-kճ(n��v�E��ɗ@ t �����Ha=�3{��`�㛆h��%�L8� m?����ܿ��(�K�������[���~_ƃ`�v�?����+%!)�R���@��d?r~�MJ�Ѿ�^w2�&�K����D�<�b'����^�[w}P�A�������8��hȆ��S$��׿|����Z�0�h�&��������z�왧~���
	%�Ý�v���\'1]GdcBG��2L��Őd��?Lm���bPVCmMwu&�g�HI"G�Ɓq6�C�W<���H]���S�l����0����<k�%��\�i�j�����ur`T�f���1�@*\��,]!�,�GA�*}�A�Kv�h!*�6	���9�I��}kaj�ޱ6�SZ�Lj����]��A�k��;d���1rM�XK�g�ڳ���O��O�4�I��@زm��h��a9�e�K���<ɛ���ۣ�o?p�Q�7m��� vj�}�����G<���;�,Sc���VA/��^�S:\G�W~o>�}<TE�0N�-C���Fg"f�9�;�*ϫ="�䑈�|t{��K� Ĕ;!�r�K�� �TI�#rK�r1
9�ᴕlC�GWrD����k#�����̊"QL.f����P��a�\LY4�h��C~ݡ��Pe�L�H\ͅ�!r\Ɛ�΀$��>{[��E��y=�A!zߴ��"�#���E[:�K���s�6���*���Pc���D�jăڟ�K}m�K�a�
�0ȞV<�9$~YM&9oɟzN�^���%ұkT�B'�-��n9"	v��̔Ο��ȍ�H�a��*����Zq�M+�'�AC�^+���2FƠ�~\���Ob�T�i�	����5���+���֚?�y
;��'���<ݧdt�`l���U �b����Z��4 ~����ٜj�uh�O��d�	DVJ��� F��e*P���!��Z� ��s���@��AYA�-~7��:���[�BY\*���"r<H� ��"y�5�H�x�u�N�Ju٦�q~����eC��Oa�1��o�_џ��G�M	��\�����u9�A��ho)�V��cϷ��]x��@qS-С��"&��|E[`�b=':l����Ku�ީ��j��֚f"9a��@�}��Vg�����j�T"��]� /�mD[M�v]��*��.?6�J ?�#�w��F,b�\��"鵲\L���Pvs���7�.��O+�վt_�柗�/5�^�h�	m�>d=hd#�g5��l!��o�߼@ �%�9� Z�*$�(1GˣBwއԍ-�%moNQ2�+-t�����L�v���h�MI22�ɔ(X,�$��hlz�
�c�=X�	�/W�����'B��U��]5Z!��ӫ���/%�Y�t'��6����h�{��h9H��E��040�>�{P>��|��he�.K��|)���� o� �Z��j�!T��92t�%k��c�oF.���+5̓1�J�|X���m�����p�u��X���TQ#��C��g:�<�,�>&���Z�=V*X�b�,�؆?�"�Yӓ<������"\z|�����l���K�LdѼ��ۂM9ﳂ��.��g��Z^	gG?iA��(�n�a�*��{�~�>���W�R�
3��P����Q��;#&Vc�F��kO�%F���}��	Ƿ#Ǧ^� 5�F���j�?�}	i_�Y�Ę��a���@���P�GvI�~�؏�@r��PmZ��K �Ng|�$%W�T�n��C�#��e%���۰aV�BCk�T�+���@��B�@��"9!��%ך��6!�9�v�7��@�2XLAȜ� ��N��衝=͗�Gz��&nd,r��_D�%劌l , {b ��f���=����?�o��x'*̹<�V��tm�%`L�X���}�H��=�s�U�������3s;�r�����)�y�ȍ���Ѯ
=~�i<o	�����#��F
`����+��2`|hkFX�>����E�Bd�|72�2S�Y7tߵD�{8��:k���{MOJhZ��p����ˣ�Emd<Z��9�� �0�R��#F�\R)�ݖ������%�	�?'R���+��,��*�F���ca\�+r�����NEQEi�����C��у���^�=�ȿ����Α��ÿT�e���ًcGj*u>t9�T-��$�C��v�0=��h#��֙� ��ڛCJ�Y%s��[琟�꙽��q�&�<w����#�����/ne�a��w��ZL���(g���2��������*O���=����$>ӯy���H��/o��0�k	<9�/�����:F�ǒ='wW&1�NmǘX��P�ܶ��A�9���Q2�����; A�ߥ?���ҿHj�%+G!��>����A���� é�܏ƥ"����i��)SX��ג�)3��{�/��ۢn�37D�6qt�v�?��6�W.��T��p���Bx�%`�^9�7Ҝ��[�Ûz2v�8f/E6��-������s�~�5�������w�Z*�aO>��|����j�N����G�z�=n��׷��-M,�M�ٔ��;�3�P�݄����Y	�旍��#Q��5�s���u!�e0�-ح���B}���e|�;���d��8�����e�.���VvX:Ja)f��e� �%��P����3��~���jbh6Rb-
%qL�vծ	f-+ @@rE#D���+f��#�B����`O���c ���0ڀ �n�ͅ@��/�ߔU`��E���e�iI����ʿ$�R�L6������z�C'�W�{ Ň�}L��/����먟	;�DDi����\�� ��sþ�޻����\N�X0K.?%���W�L�q���H<N,�J
�����T�'ν�*{�d�U����"�1N�k@�*ɾ��	�x��i�O��+��ˆ��X�<�ڑ0�etZ�l�5�tV%�9$|���]Q�L�D��wK�I�\�-ZWl���h�~����wXo��B�� 9�U�ʾ����v�$�;�fh��(��)�\.���-Q�)�`=�.�b�ny%��l�
�Mޖ�g|�a�����N��O�����'���Y�8,�����`��Bh��z�T�(AF�i���פh��h����L�ƹ?�.Yj��b��[�/��рM��?���͙�d�4�v�����5��0���[�((�^4�Kz�B��K�������;��)7>�{Դ9�*e{��/A�@�^(���ݛ�"��Ç)��!�;f1:��
��LQ�̘�Yf��G=�ƙ��CNn��E��r�J7Qɹ	⋘�u��	|�9=�e���@��k� �A�H�� ������p�G��˸
��1o|�������1�f����N>P!|p�A7�91E��K*���f'gvyu�nluS��*���dn����-�q��mH�)Lc.蘞�t�f��c�%4�+G�º�s�(q:j��u�,}�j��E�R��(�c��B5����/s��g+�cq�ť�b�PI%���TfTNW�v�3���xƁ�z��o5�J�K�-���'*�٬��k˻��z}��	�u���yBg��DEy�6��p�
�N$��adX�X�zX:m�Y�2`J���>�3?���D���%��|�� �?2-'��s�,�=�t���޷�S�m���9��`�E9��W��W�$v�a�U�]��ߐE���ըl�.nf�}�J��l��XT7���<�sײ���:]�7�<��-��EG��\Ch۫ԍ}�;5�*�W����%A)i�/�L�'�%�:��WW"\�$
��{�6���D�|>8��D82�&���"zE6�Z;�XY��.�lC�<6y?G�ma�](��\)�7
&0�pQo�ht�Á�|��5]� r�D���yPL�� �U�ۑl�f�s�r�&��;��>Pˈ����@�8ZL\��rW
K�����뷐TSk�lE��&tvs�|V�w�cfƇ"^mA��۟KѧN�  ����U�.�+Ǎ�}<Y�'�����t�l��$m��}���:���rN2H!���x�uV>�>��Mu:�0�I�9��5=�;;w��::��l�sA�@�Dw��X!h�5�-6�Z�PwD(5%�	z��6�����R�d�PQ��0���v�
S��{�V.��>�� �8<�A�l�0aO�m	�\�0r�!&��h�����$ �/3��ld�o@к:�8���t����%������a+V�� a�Q===��:EZpTBa!��u�\�����4�������2��P����]ݫnŹ��Y/���^�Fm��IW���C�����"u\����}Z�d��8]��o
E��}DR�p#2��{vޢ(�n6��m���T�+[=� <��QS�������D�D�4!ij��Lm��Q�K�8�/�����`hr㞆��!]Dh��&!j�
���B��=�0����&�X���YBS��8��L������_��KWe7��8��;~1d���c��2\�6�!jQ�-1.^bg��ē�Ռ�6��`�Y�s�A�gt�@�@oԡH�U��X�S$�^Y�%0_|j��I�v4�"��7M�t���ϖ�\+� ^q�g�|U�!��$Ʒ^�ɇ2�kA[w�E{=	I�����~4_~���̴)_̃N+�Kr`��#����dyQJ��uHqUT�E�{cmp��ӹ�3Z��c�/dpp��%��n�|{i�y�2Ej��X"�I(j��Ι���A�!5-��k���}%5ZN7A��q%U�0`�b�s9q=�*1��ڵ� j�(��;$�j���1��nL�$�k����z!#���v�E�F�wϿ#*|N*�$zs�^}.ʱ�[�&8�.e+{�¬p�B\��9�.�5�J��_�Շ����g�o}��rj�����_���䍬�}�G���]#��B�*��f�`r(Ϧa7�YsM���I���������u��m���Z�	��7P,oJ�V%��H�ܥt���}����jq'S���nZ��*D�wǇ�)�=�51�Sx; ��k��ac'�ˉ{�����)�Pb���酐E�Q��'���6-Pk�9��"4�<چ�[�N��@}����ǿ\0C�땾��(��{���K���c�5~wn���$��0��y��0�m���L��Ǩ�'P)��CDQG�;��۸�L\�[A��Riq�4��n���)@��n�\G6���Py8� �ۓ[:�%�{�����k����uδ�2z���`�=�BH�?���et��ݥ��ڧ��"��e��j[t�x��9(x���-�}�i��=�̏��^\�sSe�����΀����?��l~Nv^����>�>O�X���������gpؖ�S�m���x�OU��{]"�������l�����Ņ��z����N&ڧĎ�>j9	�(@9Ҳ��}�G����}�	KM<�*��myci!W��ߣ9�W�h^�*�JCA_�|㒻��Bq�c�F���7�`=̱ކ�����4�-",C�D���]�\������6���n��ˆ/��z�P���f�g������63��c��t���q�^��M�����^J�N���b�5#K�H��4_���g����[�F\H/ϰ?b��C�/�g����`k3�����.�B����}��g�s�m�1�jF�;��V)�.u!3G� �~��AF� ����Ѯ��6'��Z���6g��\ݣ��`�/�����?�B��\	j��D�sv��u�F���/*���u$���[�TP~��5�·A!����� �$�:&����)yڭ�B<v�L*�c2��u3h#����:�}��n�B��X�[	G.+�7������x�@��F�5��Ul�k�객:ځo�@�M�����-Y��E!���u��x�"M%әzz
�Υ_�Lƾ@��j��������)Gfm�7�2�Ila����f�܅i��V1Q:*g����cV�,���4�����[_�u�hK���Ż�����nf��0�w�X��м��܀/<e�o�/p�"�~�>]��d�k(u��O(8�� ��$d�QIR�	��S����e�M��k�'�P�aŏcW�6�`�4+��ؕ{�[{���'"��9;��r�AD,�����Z�<�vK�.�6V��ynb�:!�l�uJR�59��ɵ@�]�r7�e�<�j��f��%h����\?f��YP��l9�a���U����?ר�B6Z�qb+���1ow�ª�O���#�r}��V�p,h��
jŮg�U F�w�h*^�h�\��ϔ���k�\&##皛.�S��4��Z�*3���R��&$��#�/�;n��+?�21����O ��=c[w��g��lv��M��>hQ�b�8��?�ƅ� q�L+����t�yCsS�?����E�:���1�-����p�aA?�_��Q�>wЌ�I��mp�����ǣ�+�v��T#q���[b�\u�+.]�g���ݖ�d�hzY^� �y3H��4��f��ǧ�P�~Nz�tw����8?���YOh7,#~�f�<|^�ie���Q�C�VT!F� 7��B�a�x���IH_�'X���D��K�>8�Z������CΌ����|T�c��o�Y�y�g�h�����S|���=�<AM�K�6]�	4���:�q��׬��l������ՙau�e��C�￙Qݚg��jG:� m�=�g��W7�c����fZ�mR��q��@�D�4��`��e�����qX���.�Mƛ��0j��t�jR����@�S�f�bs!3%�u�1^r�zF�NA-��471�`��0����3�h�_$�~��bD�����Jt���|����[���^ϫ���s����)^e9;��Q��r$�k0hf���2��q��46)i�Wc��	�7`K���i4�+hVP-r*�?�ȝj�T}]�J
�� X*])ǷLOܕq�w;v�H��v�_ɓf ��@��x��m�P�mc#�+W��f���#�<
 �	��K6�������)��8Ɔ�SQV®�ٞ���fR�_�F���b���ժ��w��0��Α%��`T�Q��P���~����L���O���V�w?�(��<@�u`���=�1�W��~�o6�T��ۉ��7�$���od2�>%~Ⱥ��l"K�����J.��}�(�3Y��c
5�f�k�fߓ7��[�L�Z�] �4�C�6'v��O����ѳk�OX ��RC��/~O�P�$�<�ЮÞzbzb'ܕ����7�)�c��!��2(��3����7�η\4+;+fH,��b�8�`�g7�#��3գ������N�N�'��Yt2 yej�ߌw$y��G��:�n�8�����^|�?�ئ�T���(9C��!�1��ߟ�/�K瀥��5�`@B����X�h�D#��ݤ���ZN��&�6*R���=G]|Νg��Rc%ūA��Cڹ��Lh�7�Kp;�{���ܗ1�7��P)\��1�ƞ�����1S��j8D��1�p��a$|h!�76|��̼H���Jܘ�g]�O��6�G֗NW��1��'{���v0ᝍIp�M>�7�n4ϊl�	-�����]�9������xG�L� ���cpi櫶d��?Ǐ_�Q��\m�Z\��ؼ"�zI&fޓ��3�;��:'���q,�_�7�JN�����I6w���<WƓ�/���pq�APM�axd�{~3�!f�\����7J�8Z��<����Tl j�[�A�s2���qm���Iرa^��Hhpk�ПC~��/�Q 9"�t��c>�U0��Ap��U-���Ԛ�f݅��H��=�\�^d�د�1A��`���w�VE>*J.=[Ɨ����.JZW4��m��0��adxa�D�~�D��4���q���A"��
W�,N�z"T�/�J���9�?~�ʌ����/Io㦆1V_!]A�ߋ��?���A�Nh�����A��1��x�c��;`%�����aq��u-g�$)�}�G�7�,O�d�!WK�7O@���/�.;�UsW�R�id�Fd��k�L�B�x�wv@&ykw1����a��Ee$�o��{@_�tׅf�>�u?�£)H/������h�*����&3��xDk�N�E+�c N!������7cz:�2���?J|���!K�����<�0�w�M�q˚P��%Y��-�`_c�ۉ�Y�S����ˮk+T�ī���?�����j�L�FMFW{3J@�L2�x~�e�����}J�Xz�=3��#���H�0s%�ů�n!(��[8��Ex�*��:�Tww�<Toɟ��l���X�M����'���4l�`@�1�\�5����ZB#�n�hoCׅ>y�yoO�g8�*����	���@Sc��"��*h���;�7�Ŋz���9/��5�R�b�A��Dhr�5UnT���YtD����Y'Ы ��8�M�W�^p ��#��׸�:��+�c��H2�V�2�/~~m~ǘ���8Hq�Ｒ4����v�����O��o�H�W���#�WN`I��W����"�g���bE������%�T�4���z/*�v��/@��|�/��Kl���H��Wns�^�pZֻa]�#�"���L��F�g��Ä�;�7�k�J�i��(��7��E����CM�H�`��(ס�ױ#'#m����\��>6�[����ib��L�{��e�T��$ipK��B`��<qv3���d��Wt;�(��A��P���{��\f�A����ň2ts�;
�c��Ԝ�E�Ϲ�� ҳk��J�:�G)c�+r���4߁������R��t;�:;T[����F+����|��`<�[�6��=US��P��)����#;���<x*���p=�8�����u���O��gS�v���c��x��i*��i��2q:����&o����j���vG��Jyw<�*��"_E`+�_j�8�0����r�W�*q��3��O C��Gn>�r���!7�"�xf-(������0hQ��%����"���#��N�ժ�g�;��b�򍔛n�r���Z`�#Ȫ⚫����[0�x҃
���BV<l���%�c�N�Rtԍl���s_�U�@ v[������3J�ɓ0�i����l�J�C|+b��O
.$q�K9��C�=x0�YdQ��!��*��o�a^-~��~�"(���;���yDiK/��F�Ho�ܞs�����XU�.��v���Eh u�!Y��������,g���<����%��������p/���?�BWi%���l�d�Z��[��^"@�Bz�	� Oy��ń�������K4���r^�T�3i۟9	��y\����<L��^[_T�u���8�+�$����m������1�t����s�u���D_吭�����o-=ci�U���J
�"Ks����U�o�#��&k8u�O۶R�,�8j�}q���o�o���%vNN�i/���.ת\`�Y���5y~����,��+����P_Q���'�/���7����
�_�1�B@^]���"�P�Bݪ~�^����hs�?Qi�8�nO62��q06]�7���LLs�%l���� b8e�M�(�^�)ZDt��Q�b7�řZ:���zb������Hw<�YS[����]Q\j�~��Z8H|z�PFY��y�#������W�,�Ɠ:o�~��F��3��m�?0�~ւT���Fv�f�-�RxH�<����۩���P�װ�_��o(�	�A>��Ϋ|�Y&xo$�:��AV��tkD�\�YN�w3�dco\Z��Z�짰��b��O�H.���Q8���o,�+V]a�����Ͻ�������>#jo��c���"��8>��M�(Q*Տ��$��q���U����>�Ť#��N]~1�R8�WF�c�����<(KZ�_��VV1ƹ�	w���Z�N�-�[PmC��g�Otx�k4�}�Y�1y0⁜�e�/j��f���ܽy=�����NI�֩>����'��O�*�]#E��\�W��)�j��˜�0�PQS�~�x��+2��}f��7��=��ij+����*��j��P�9�X[( X<���PV�u��U'��1��΂N2uT
�F�[�{a�\�2u'��W!���(����kf���3��@�,���u���[OTLhH#�l����]˃~�S�0�}C�Ϳ�Vz칸�L��VRJ�O1��Ӿ:��&��1�$췧�B�7�
~�t�vM��?��~H}����$6t�R���?�+!�z�?�c���D�;η���ʯ��B���Z$�g�h����[)��Z��bQo��w$-�PJ�\�S���=�Mi���6LUȊ��{s5c܊�gD�B��8r�?:��.�cʖBid���W�"��q��X|
p�B��Scr.��Z���CQܷ�\�$DxO�6�W��De����fw�_-�����F�$�V�x�������)/[>���b��IaV�⧿z��D'�
��m��Νl�����d�6�(���o|�U�zQ����lh��N��'�k-M�0�ߓ��w`��Xs)r)��[���P��f��״~=)�O��՘N�8E�L���T.�4�WL(�b�W��w:�wtG�T��h^{ �B�x���s�1���\0��
��k}5�fwx��(S���ZRS�)�5yb)��k�,��p��^��'y����Z����䭡O���J�j��u�l��`�����Ǜ�;)��{�uc��*���z���Z�����" 5<^�v��@�#�R��n
�������.�TD�<�JD�����-�l~龍!I�S}SN��tB�%��?@&�����)���uz�5fC^��N� ���{�Ęx�Y��A%�H�����/;��F����Ô#/ZY���.���p���7��Q�f��5r�"�~B����>��Lﬁr(�Z� ���by�-z.?5/,�T@Ɖp�`�n����;�+Quj��"UކX�'���OB������FI6i���ΘD��C��fӌAC�}~���QW���v�]_��pYIb��)@bX<u��,nNKn6�R$� ۅ2.N�Zx�`��bS�M������3�mrmK�j�o�Ir(x�&74��F��N:��댼�nI�5xN��ݫH��`+�b-�*>]�|�hv&hK������%4�%�"�F��;�C��|=4,'��xI~��N�Eg[v'c㍛�Kb�~�o���|�q�*L��,�'l�"�64-����׿jk�t�
�O�:zv��[`I�0�l>~��7�Wew*Œֵ�?�V�����>ye_�L`�F��H0��X��U��e��CV7F��&��&�u��&�����	��?b��"��W��2
o����r���t�!��@|�d��le!��8��>��p$��?5O���|͍���;Y~�Yr��+>G�`v�c��f�
/�_�JYr��l��
��2��D��{�dԌ�U�����������4rl>_�Rr����u�w4Sf�\7+���R��5����b�h��(���oqh�>W�@����Xo�1�;����=ND�@A-����O�@kG���S$J�jL���^q׃�V��Oĉu�j��di ��wO &+��X��g"��D.�$l�5X�&N��L�͢�d�Z*m��q�5�8�3\�Z��@Ǫ(������Cw`%W��%r�)4����/ZH������Ϫm��I�ϟ �o5{*�u�s9X�:�:����qS'��p���]�g�#���t%`�{�U�iHz���rs���*�O�f��N����0�w��m�ڿ@���^�X)V��A���D5�Tu�C�4������}V	�/���SP�i�,�襗WĄ}UD�۲�9GS�4�L��E^�����y�@dX� ���V���Q�@(��[k�7Y[ufqnc�G��#LP%q�:B�����v}�ʖ��	~��F�GPn=���;����V�7�y��ܹa�=��>���1�>eO��뺡��ӷ�x�����k��M�^�*Ŗ�J����=v5�R���D�@K<��P{�[ň��q�}"'E��d�>�"�����,��E5t�/b�`�v�U zH�c�2h����,N.��g�4���`�˸�=c'�s&6Hak̀�5O�9�_"msƳQ�����|�a�ؾⅽ���?a��̝�"�Q�,b�L�*�Y*4��P�o�H����
��-��sC��զ�t�iC)���K�I�{��ۋ�'����	n���j��=��3��k��+<a{�������A��&�4A|D�������C�EnZz�cU3�Pc^;hة���2ר}���`��l�e�H�u�G5r�QZ5�H��>�
M�Ăَ2�������a����X�~Zѐ1�ܗ���@8��kt�鋉�s�R��S���̃ �_ @8a��y�T���.�Z-Ē��kL��2��#l�u���u�>3����l�,������vJKC�x��2
���8�����蠕JkXhO^^P���|��h	�&2�[�M҄�a�/K�\��	��}��T3z�}OR���t3����Q�fx	<6�-Q�9z����7��3aHUG�=G.�=IL��3Y�qp�z��i�B۱���W��B�3J#�|f�ww��h��#$�������l,���K9�HG���w$�|:��(�t���L��3X�s���g$a��L���>�<W���mB�6��<�
����j�rw�2��!(f'�hQ@��h<�������*)�R���}��b)t`U�'�iA�\�����@�2rf	Ke*�o�]]s)l�\Zt��%oJ��.w�ں�͈h�pR������lN�=�rgY$�V�˱ aG1b�ζ��Ɍ��S�~�З�0B�Z�@�D�-K�n�p�ɫY��EC�����b�q���Vs�?��䩋X.�n�y�$w+��D^�М�30`��L/D^��x}ʶ�c���X��PQ_H��9���ӗ��+؈��8���v���m|.~'�W0���:�!3�� S�>	&���#�}0��~����b�$u��ms�%�R¥39��d����A�y�P`���j#T'd���S~�6pý̝X��PN�$�(�ª2��Y�5�S�z�O�1w��!d��[��mXr`��)=�~`Q��򢤂�݈�j8�	����E��ѐK@R]�� �����Ƀ\��<7
%<`�T���D��3O�ڎ��[/�=��lD��v���'|���G�:y�[���W�lL�W�R�э��)�5�����_D�"�q*Iц����3֓w�]���'����|["h�7�Գ2�h�hk�%�����F�a�U,��ݸ��m��:�1��s������B���e��/-@Mm�9��W������aU�
���Y�T�rK�`b��Z�P+b��FQ����XВ+A��m�尶�R�>񦟇������1NDr|rʻ0V_@�-�p�J#���Lh�����yAf�m3�0x�GfvԇswC[:6�[�I_,P�JœW.~���aoTA��X�D��EH�	��R�k��V�ݸg(��5�Ƙg5뙟�9-��|,BX6���܋R`���dRv������Y-�YF���@ �!u�o�
^��c3�R^>X������s�z��3���ݯ��+a�M�rW�T7m(xj�L��S�E	m$f��1�icMlC�!}=�zӰGq�����@ț6C�:KԤ�|��p���A=���}��G���SШCs?ə?��6����1�{��Û��E�iVɝB�R����\,s��#H�����:�c],��fp@��u��Q�ȟ��Pg=
���iv
�1�ɹ������P���$(`��N���A¯�$�jp�e�x�4D<�B�&��>�����F	�<�3���W?eH��8�՜Z�VQ᯲y���9T�D�O��=�$��$L���A���+���L�`��tЩI�����˼ǯ�8�3V<���J�8QSǜ�5����ҥ���U���-fTT�y��ϯ�7�p�i-�Xu8 ?I^���sw�M��C�u���5��s��������i@Bs�{�I@�Z�d�C�4�!�/�$P Y�Ե"V�7u'��u	�����37�p e�/�z���.�V�>HE���h.ZD��&r�,⾭6��L�'�|ؗZ�3EN��n/we�,ge������mփ�Ӓ!xu��F�A)w�b�|)-o<Ũ`]CYkjo~X4>�\R7�V'�8\N����vh����)���ҷ��o��3}s�����y����"��ݷ]F��*��1���	��z9Ԏ��|�E�,�I�ЉdD���)�N���CĜ]�1�,�T��S�|%e���ݖ��XmD���Y�d���h\��]��MA=Y�@��UIP�դ�j���O⛓��Н�:GЩ�@l�����_7�F��|Y��(����me�ٌJ5�a���e�C�`*��k�p;��on{�,����y�-���l�7?�C_ ;�N�:�Ŵ��PT��G��n�/$@�Ƈ��gX�W��L$�A�3�Ő��������#���z��q�tۧ�h�d���U���&�o�6��}t>�^{'�"��3^� ����Y���)h km`.�}�T�JցN���}���o�C�w��;�ڜ�V�bշ��Bw�7�M��[�%(�Ц�p���ud��ز�6m�N7�@g�<Mv�+�9�^J��Z���/:�����o�]�x@�֘��Oj�����i�6��2vj%��M���ŕp�ٓ�� ��>�Ri��c���:ܡ	�;QX}⒦�����|f���_hJz���܌.��}-<�j�h�6<�89�1h�� �1��t��D����iy���2K�1չ/m���p�גF�'D�h뽡P���f��]F�P�	5��X�Tk���y�4��Ȓ!�	L��_N� 2N,fu�{Q��A���
:n�A@P>�h͙�;�E��E���x�q�9��F��;����Ķ�u��]x��So[����4F�T���ʩ#��@kң���˦�3��u��!�(Q��s'e�=� ʉv�r�G�`�F���ѐ2|�p��t�~%mk��u�DH�/y&~�����:ӭޅm>#����%an3�V�\*���w��d�)��d��������I%��_�g>�btL����(�v˙���]r�|$h��/�m�e2����� ���j����,�W�*Ȓc�
����q.O�Ċ��Iw��]*�X/>�Ɯ�� ��J�%A0�9�@��9CA%���Ǿ�R:��k��7��G��w�Fla���0��@��1ݬ�'zY���1���\l%��ͣ�\&{�B���s4�L�R��W�x�w�2��Jv*�O�����P>s?�^�ț%Vs��f}Z������F��/.��W��@�Ҭ��>5�1_��t�����F���*��gj�@3� �0WĽ���-^�;��H�gW��}E���߱��r���!x�߷��R|�3���û_�}-�-�z@�Vw]�)���)��4Mc�TvT/"V֧u$���_G��≾:Tk�\Y X��m��e�j�t�ޕuA�ҹT��eۈܐ ��Y�1�yC�d�;�W&s���f3!%����ūh�q���&�.�$.�n���W~�
 g����j18|�Pi���W?>_�v�"y�fL�{�
6t�aT]c�?t��8M
����LשE����؅¢�����n�[���*�#[O