��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|۶��-�E�8@|Jq�^����`څ)h�(��Թ`�4!�s̆d���GR`���"b#	�ޯ�2�������_'/|~� ��� ���^����{h/f��Z0#��G�=Ǹ�k���M:��i��a������bH�C��q}f��Q�*c$��g"�o����O��(|Y�3�b�4�F+�\��K�P�&HU��+4�`n��~̕Q=�uJؖ��(�9Z,Ua�����7��l$L�S)���ڮ�ȱ�s��*~v�a{�[�Ɇ�m��z��K��-����0Ë���,8���a��a$s]!��2,ڥ8i"n�C�]��<�9�!VX{m �z�+�HkK���s^��:P�D]J�WY�3���Gå������տS]+��m�/ݯ�Z։�v1�����5Y� �����팱s�}�Y�,&�1_[�EA��+̈���5;s���� .�F*���?t�^d�/�����Ƕp)�$�\&to����,_&(M��cO"��߽��ET	v�awz�|*q>rD0����Lٕ�5�m�5� wՊobb$����ӫ�{�a7>�!�6f�m�;�#4�S+n1m��`~�H���$�F-:�	YѪ�LW��j"� W�ǊQ��$�mN���>�nƺ��,R+�y[����ו��/!�!L~�ju�t� ��ep(K������"^�.6<���却�3�1lI�;����r�y�=�&t�7���P�b�də�gâ���#�rږ+5�J�>oX8��K�G޽Nsr 	+�+�;*DLL��/j�\x
0�*���4YX��x�^tqXY$!S�r�`K~�7�}anJ�-M`.�u�VAB�\F��M��s�:+R���0�ƻ~���⥸�EO� 2Z��~�ɀ�K��I���K2B��<&�|"_�2!n�S�?������C���Yr��"�0!·*��}T�j']��x��P��Z' E�C��]�|X�u�4C%r1Mf �����>唯~�[ٞ<�ҘN�<�+w]_�� Q�t���PY	�T�E�\�dP�cj�_>���#��m@��'�,�]El�$�����������b���ɱlsԟ�^	/���x���a*�F`�B|,��e�X���xh��\���3z��_P/E��l�E�?�M��j��O�P��ƨ�H���F���>i\(��n���]ń��W��I�0�L��]Tɔ�(�HI�'��A��y�܉ NδHg��3�Z�̀�J }�JV�`�6����Q?�{���&��A��$-��G��z�=�w�@R �j�{��U��{W6�Y���Y
29v�O;���b������o�X�6"2��G� �\�h�D���r�nd��s�A�W�ě.�3_��PxvC���+�~�� ��clS�Kt+�$}���)��)C��,-����щm/P
��;�� �' �_���[~];H���S�P/YԌ�&�?(cXv�@`$�;�¡��=�n��Y�}b9��!�R�����@���p�CrDO�4���Ɗ�x,DObU�P�c�1Em4�U�2<f�}�;�*��K��rՌކS���4(�1�ǈL�g��d��br��)�?4r�Hϡ;c��&�Z�����f/d���!��b��d�/}h�n��3�[�z_�B$)���ѕ|�m�'��"C�fnMݞ)~!��Q�Ar���0�h�F|m/�N(_��/ -����)����1�'C����׊/�4��o� >qy(��>����d�e��'8��?qC���?<P)1��?�z?R�\�:�\{���K�w��m�+g+��d	��<uP�'B�,3��P��O��	�@�6�{��زn{�]xI�2Gm>�ʱ m3�0. �[-��;��HK���d�.)pD|�e�O��H;�}ܪ�uJ��E��'OP��"������s%{R8�<���!j1��3{�]Њ9[�]�&<�ȸ��mi�O�.�G�c�V�7�@�l�K���񌇺��PV��yeK�ߕ�΍o�ȶfO����?��ֻx�𦳪iC�6�}䐾8Б�G�E��`a�����p���J�����"�^�5P`�ݞM\�:����9'YzB�5τ�q"z�� ch��2�֡#��,���� �������0�j��`O��XR�y�I���ɀ��%��(ד���\w�#y��λ��Sӑ�t�l�P�$�Y���A�3�j���zA�������.��ͪ@pr���6EjL]>�2�����T�oț���j����h_5��S����\N6B�6��]*%������vPp��)�t���V>��bךq��-F%�%�G\{ ^t�9�V-^E�14��6�$8�9x~M*� ��Ba�J�G�-�F�s/x-S<�ɐ����T_)���1� �@ {|��䞣l���� �E]l?I���9N�����	��b#���M��R�8α�Q>a!�O���>T�/���8	7�@)���jC��BΎ1�lLL�%�9(�.t�0>A��Au�I�͸GV����Xl��#C)��U_2�q � �D�Њ��o�F���Wi�0�/:��hiYS���2nʃ���7��l�L6~��J�����!��庒K�c�-l���:�[��b6Q�w�
˔A��إi^���`hH��va�4��S�e	�t��Nf�����qP@.�Ϣӷyڔg��p�]/�O%���m·���z�6O�����K(H�,���iwCf���T���+��$!v�u	!%�� .�����}��SnH���s-�"�v�~bYN�!~ګ�Ȋ�6 x`����Hق����H~zF=��G����,A���E}�����M�ܧwZ�6���׺�ے���%�ǁC0�͋T������s�w(�.a���Y��)�z�V�ވ��J����J�-[�)EO��c����)����	����#JtFO�󬀡P��!ۖ���xT��3��}�"�#�'�=��1�8D���c6�
��"�[4t�:4���Κqrd���ǔc��!nmG+�J�ګl���2��$��<7&r��h'����!I���c�.�/?���ue�5_�M)�����V�o2�y4f�,Z56�h�`����p�|��W�g:p�G�.�^K >_&���=��;�&�[��Q�g�t)F6�D�� }g&�愭[l� �D���[��Y �k���� CH�q#&}�p�Ԉ�� lod�"��(�gh�w�CX��N��:�u4�{�������Bi&�YOSF������?�� ���f�l��\�>����a�`�&�TaF��
�`'(D!>����D]����D]��cQL�O���F�
����CS��.l������Y��g��D����N�|���h�7l���Nx��mkB��߁��g)���|ۖ!V���Rc�N�F[=�y�b���i�3"�t2\�}Fp|Y��Uj���Nu�]E�'i��(Q�'���Hs[d %3�ޘ�b��u��zl&���	f��L���(�V�����r���A'��������.�+�wΓ����d�2�mOh�zFk�REuC 9LP���lW��	X�(a)���=H���C��Z�ڪ�N���k��س>2;�p�%�Y~�)�^_igMH&d����F��"��ݵ|<��71�H:M��l���G-����nN��a��,ú���xY�J�sAR���Ap;�w,Y�
��k�E��&�RЧ��H��/1���:=80Õ��U�-k�x��h�HI�r���~.W��f���!7���=���o�Sʰ�����<�b�a31>���e��v��@��y�7eo��P^��� B����8l�	{#u���FY~����֏3�SG�(���6
�ڧ.OX��d{����J%w�x�2)��l2�A�[H՛���x���*�qоRA�R�H��emz�c P3J�Ol��L���r��H#�maYt,7 ���N>ΌMZ�w���OdP����K�Yk]q�4� �ATv�g�,��J�0u���%뜦d4�֭N5�u�>+s}؛�"P�2{6��8/?I�[�N��l�ľ��R�����4J��ں�-�X��<�����|h�����O0�;YMa��ӭ�#��K��c�J�awR�o=�[������j�9�<�#p�ݏ1� ��v��a��	.��.�S�����BO�+���:.�-m�kJ +����==���<�����-K}6'Q�R_��X�{#�iT.�j�YW�o��.`�e�h��T�o��}��?����r��	��BP��j!�5�~Ս�p�2���I���b`3uy�����@�8䭨t�lY�q��7^��Kb�@�Ae��mw��Qֵ2�Q��7G�87���-EG�-!���01�.QF�$���pɫ�v�"% ���ro:�%@�����hKL��]jщ#9f(e9�
����U9�:|�]!8���*ӛ�n����A���`��%E1p !Ի��$q���J�4�#��ח�$��RG�K�����o��P�����;��i�E@�_�������kr�7��ee:ΌO�;j���N^�T6�xyՒ��֮uZ�~�;l؈b���r�����Ћ�	3h��Q��Z�J0]���F����������H�'D5*k}Q��w�.B��/�9A�����f���>Z�6�H���&�/4���d7X� ��(�#Ra����j_$1�
�kDϦ�=R���4`t�d����,Xʶ�q��&��Cu'��|�H�:���]�,�7<�ǉ�C��p�/N���*B9�4��E>�HZۣ����X����%����D��
���iTk��>����m	�g?�tۊ�⭉*�׍��x�8z�H�;yb��m�WYU�ɯ�K�F�-����co��Q��
M��B99]����ҏTx#ϔ�ێ��w;]�����h���o�{��mO+�z=�A��D���d�����Y7���L�K����^W;�U���_vhZ�z��R��]�y����Y�
26�C������g�����D��NS��ID��+�-� ���8Z]H��ĳ�2���p�0�W����n9h��z��"}�;��,���zC��� 暴�Z}�w�\�"��=�z�Yܼ	 ��|���Z����+�	�%��*�����]�4�-sSI�^��PI�Ȧ���*^���B(� SN��R6��4�90�
Gm��ʎ�K��V��|,޺���2Z��v{�Ɲ���(�ĠH��u�4/�~bã��0�/���f���Y+j^�5ܻ��5�ph�ƙ�M�(���} ��5�Z�l�,�ޛV�����0F���e����<�6�Kc���Z�s�lP�)���~4��q	Q}���'�H�<G�`�~
��m� PC��j�c�.�bb���J���i^���c��c�CyK@�p�=��7ɺ��(�]�T.K��A���/�Ox)oҮ���~��c���
��D~�C�8�+g�.������!��??<q[l27�2��w�������3��J�����r0ldj��9�t����Z�~|b�&�sr���2G�O|�AY1,[���޳���=����~��4avo��{T���u_��/���ꆿI3���.�	�O&� 2֥� [X�7���9v�
��gT��΀^�.ګ��"��e�?�HC��MqP�G��a��%�hv�/��>s������1&�2\�I-D ���WS��Ȉ��-��*iκ�,]9|D.��{���e9�s<Z���2ؚ<�◒����%Q�R��(qGo9ܧv����OW:̸eC?�9�$t�y(f-�)�  5��X����#TF��p���*��‹�mRB=���(� ��@��?����
"�I�{��"Rd����^��r���K��ۍ���!�wX�V���JaO\Ҥk�f\�I�"v]-+�2RB�]������wA�VMQ�`��/~n�/�%�=�A�X���j�]�-�������>�v�w�/IjgD�#}�V�~���E�T/�I0NC��c��1�ȣ�"-,1���dp������$�h�'�w�WfW��� �҉�GT�0Ĩ�St��J0(����������2�����b��	���#�2�t@C�%a<�Y7x�Z��j�b��d�
���p&��H�����Kb�[#-Ж�� �Q���u�X�I�wQt��l%�ı*�J�s�oj�Z��+6$g,RO����Rj�1�ˈ!�?��#��qF8G�R~a��b�a���H�\u��T�T���p	T�˴K�W4<�m���C�z�����y�ַ�1������E�Fo���=��ޣ��k��z�����6~�Q�%\�,�@���<܌�V���Y��g6�:���%�r6$x����n&����0W���5\�5�ɤ�_�?#��P��0o�p���~������V�dEw�x>y?�]�Ȗ>%��96q)[jGiJ���Juwz�S��t���������5�_�UA!
��+��N�Ʉ�Y9k��iG�t�4.�u e��
W��m~�E�� �8U�Ӓ/؈}����rw? I��(��]�r=�
�Ă�#���Mlv���e��}���ۯvO9pﻟ�:��Z�c7e�Ygjr�T���(��P�3���)�V�=q&�C敢	0�OO[_|ȸx�bl_?W��A��ӌr��? �i?�V�!�q���<�؜��^�7W��Z/���Ƞ�ܬ���WeX2��~ciT���+dVui�d�q�ԧc[�x�1>{��)�to�����f�b�3׶�_a]z�Z�ҙ���H_�����}+蒓V��as)&:Y����Zw,~��g�G)F���g��Z��t�י�t64�o@��GJ�6U��h&ZL��&w��p�o�܏� ��E��;�w�m�o~Yԥbw�،�Ms�ɞ�ބ��AW:q�9�ʬ�to��e��~6�M�n�(�ʛ��7����Q'�ZKo{-�[�FҬ$YJy�w�#n��s7�!��BB�Z0@�F}�Y4��P�4:��!���@%��M�(�hu��췴���'�&H�o�\\�<�d��t��x!Y����
1܄���+ff��B6�u%��sP1�>*\܋i'��w�	��h�c�L������'"	_R�\����i�{��ċ#uX;��g��y�p���l�
���ORgj���>'N�K������1��K`�q����]��LAD��ﾡ�Bt����_!�C-jVCDq4���%s�Y���TB<J$�Z^�Yo���-ʯ�6�浟�F��~��t�����b����O�^�����}���]�R��N����7����/���*�>�V���X0���~,��R?@�w�-%�zsx�k,�g�Zs�#ɋ�%�c;�@�`ܖ&�+h���é7��3���;-�E��Gަ�E�/yqV�_~t=�����g'ڤU����}_7���es/,�G�-�C
�[_��E��
L�Z�.`�p)@n�uq�^�(7�W`O9D�&NC��q\oE�km�#,b�&�.�yQH�u�[�� ��r�k�.���NB�u��E�����	��:
�U&0�~��o��6�Q�W�q���'ǭL4���<Y���F������Yť���!a5��p�lu�{����i����!���C��i%����*h��w�I��K����kC�09��O�(af�}�s4�۾������B�c{��B�6��#)�Bb����+_��AJ�p%�u���fZԙ�o��N|�S�GlU�ؘ�D����p�7���	��C�hŬ��]�>�o�(9"	�LT���Т.K*����0}����VZ�OW�H��v��BP@.��c� ���,s���银�2GN#M`�>o'O�ٱ�l<�7��Ь0�f��,~b� 6^�7��x�0x��H�uc�\��;�����`X\�$�饄�D{�M�_V}�v�17�Yt�B�f���M|�r��xI��v?����)[[�DS�Zj'c~�=�&�!��
�3ƜJ���Rl��w��g�LZ�$��ؒ>�G��^�X����T\ksn�9����7A22{�S���9�l%}|&=�)���dӽ	ކ����p�t�'/�q[!a�[��d�J���l�8@h��d4` � �#�.�_���!��J�a�Ɍtʙ�4�B;-�j���<6�b�uI���3���-X���W�Up�o�m8'Cm�KoR����i�Ӕ��K�w����I�p�!YKnl��&%a].��,m��xw@��;�1��1'|���G�Ay��j�q9�G�@f�v�{yD~�h�l�  R�S�6������Je�j©,o��cy��+�xS܅��)=����q������4b@�T�鈬��ջ-��Ҭ���|(�eSE(�D����E=ʞ�uf�#�����(rkGu����kۂ������gUk燜��.'b�PICs���1����z�b\�>����'7V ��ӕ��j������n��g�`hNq��χz������,�pV��߹��E�������z։Í����M�i�Dj�����)~�5U@6��zʦ�8��a{͑O�&�Y�|��D3uk��u.GfdW���q��ӸeA����gr�oȪ���CՐb.�w`)��s���՗0�B6���3J��Y*��؁���I��}XsG:������
�nv؎�0��%ET<.�����F�F��� #N�"&f�`H��L�L��a���?ysG�J����q�d�����7�Ҳ�F�4�U�e����Rqս���_�t�z�4���q�+�]�:�ſVS����U���b�h^�3/^X
��\*#���Q�,��3ρ0�Sr��L�D����4W��ko7Q����8��Ѿ�z�u"6���A��	׿+�Ϳ~�zp*G���ń�����BL�moK�@�b�Ȟ�u�՝��!��8�g�({oc�֌}��E�h��r�q-g(��c1"{
b��d�VD��
C�!��TWX���k�&�p��p��g��b;��͍5�,u������5O��]$� �T�
�ݝ@����"(�XIM~���x��xCi����r� ��
M��P�\7"����&���Q�Z��������L��i�< �~�E_��E^]7%���L� ĥ5�}<��ڇ�kqQWY6^ ��D�imq�Q�??�܄Y���C.XH[��"���f7�0M�,�"������y�����貨����tWe�A�����H�қ��d�F��^<�"L�ƪ����-K���"J'�\�<WLT�����k	����~�ם��!A��{�w�#�V9H:�Á9�2{���6zi�P�C�����l�K##�A����s���
`�r-�w�E����C�{�@R�r�}#֧.��P��_Oa�N���-�a��	G�*l�Z��/Q5�h�Py'pIO��X���6��ʛ�Z!^�&UT�$D�M�:B4��o��=<��?C�1��c]��e�d��|���=�`�ql�qXCo�w�%䦥���$�a5�����y�q�Qũ�;N��ժ��),X�q�@��R-BX�/$���;�f����Ȅ���w�|ݰ@�4�-��d��*mҳ�����c����{��*�|�U�T3�0]��'<�'?��Zř��с�t��=���n8AOj ʛ�$��G?�*���hk }��/̊�o9��G�N[���<y5J�G�[�*ݷ��6OW�*���Sf�@.9����/�O�lվ�Y��[���"Yގť���UQ����lv�l��u�u��8{�;=��-�lU�?������@�z���XcGbl��q_Lʟ�x�����8�uN��-#_�����ݑ ��`�b��G�Vq}`�ddW����	��T�}e����X3�N��%��1*܄��eF3��+���Ke*R�w}Lb�E;�!��SPd�}�����(�6]4{`�=����_u����
C�B���{7�ݏ�Db�k�[��$;�_j�!��M�7�J��<�`�'�V��hl�~�`C3���Sk4��M��s(��榌8P��r�l窤�����2��VH��|4����������}�U�_kLo`�P(Yfx_d�� R"��#��Yu^�Vy�mT:�Ƥq���x����L�c����1�L=ܸ�d�.)�tbx�?f�ɛ�R�i��s?��z�R¶��'��h���X��_�Z�����"� ���k�y+�D����y��	k��b9|y!nt�����9�<�{�R;-昽��O�<8R$����TL�QE J�1\�i�����~��*��ҫ�j�^m��4�dp�E��Q�G	X�s|B
�q�M ��ֳd;�g���٤T���s&/����5a�[�hF�_E�U=�j�d�I~��lT����w���4�I@���v���h�mYk�������}'k�W{�%��BP�;�o�՘��֧˾8jP���#y��a^?ݟ�yu��E
�����z6��7�����R�ς��h�5?�潚����U����+n���+,�87�P��H�rS����������W�,�Hr���S�O�:���c��Uܟc?�&��T�iJN}����B�-�P��P��ny��VL2�_V灃HnZK>�%w@w��4z&~q��AK)�u,�����9/y���v��rf�~� ~�w���1���p�/�����R�Yi�4��k(Vr����[�z͸6����'L���@�Q�a�˩ �ې��Z�j�ceks	�2��J�20Iո��@в �g�<�- ڂ�i1Y@8�0ݲ�Ʋ6oL-If�@o��C��w$��N�>nO}>�!���Vp^��.��T�4�V�bg�b�0�H��@�,�-�4EJhZT�i�'uV��t� ���va�v�.�^�{�C+�k$D��M�#��DL�wl��g�8rYߤ��y�z��6t�O9�=����o��B [��骃�g�)N����k�>D�ͳ�,�JqyT��#���d3e��+Ct/��x�1����cP��DN�1.�l��^�/�R��EM����>}n�5�-
�0���9�W�۳����P	;�r�̰���!!\&�gIz{���5u�O�Q���D�:�j�y}�M��M�s��	� /�Fc���f���̐�Y
�"ݙs}y��2ߠMW�Uz��cG�H�>2�R����f�α�;�N�Hc�6�=��ʡ���?s��T�����o*�S[#��Wu�BՒm�|�y���Bʕ�B�H�~�Sc���μx���:�JJ��G�c�ǈoK�J��|W88�}~��޶݁�rT���ޙ����^d���8&WT��2��GW��t?,;��.9+N�:��(T0���c�c0_��"��҇O��{ΐ���-|m�[A��<��)(,��`v�(^�������e~�T��*�Đs�<��Nj��Ap����C�\�9�V�3���_I/A���
�qr�nҴ�If�;��[>��MM,vFp��\��Y�\���$�'����cl'Xc��D��O� id���I<��)�9�۹�1�e�+7�O}��o�+�3��"��4��B�$�q��PV��eK�տ��
gk��VR��3,�Mtk�v�[q0[{�&�񜰊)��6(A�C�.�$U���$J�L>u�4^�B��je���.�G�T.��?[�Ü��Ѝ���|>�ĕ�M̖�^��¦����Z�#�H�^����1�G�Fncq�{'�~&�F��Q�ʮ߃TBCg�����4�,Y��m{���
Rg⳿N�M]�l�F��Sk�i���k�mY*FJh�c�鉪퐵0�c�����`�'���>-+W��@`����ɜ��j`�������}@0"}��Do�4`��4E��NB� �Q/�/�VN�Yϕ��}Z[v�[b�{�r�Ϡ(d��#��K�s2`�xX���t�ss1�;���.|�e����`���`����q3o�v�G@��f`+o`�Ҳ�l�T9�O������� 56p?��H�qZ�8c�U*+��ƭ�n�9aɨ$Bމ�sœ6�S��Sq�<�/<���35�3����լ�^����zӀ;KcװnU>޶�Y���+k�Zǹz�t��b ���xb��*�R�Yx�>o>�>�WC�����a�)|%�B�DM��|b��]�=��y�ÃpS��԰�oGo�ܘ�Y�.7�ϥ4�	�|�ґ��Ub�<XB^x��_e�;��e����f?��ir���\qv̭Y�l����^��>�ozbD��@�H�q�Პ�E=��F�Y=C�,��k2IΖ�0��YW@��~>&��M_��`��l�k�+�y��)��]�մ�(�R5t�(ڡ-�9'��B"��[�GqҤH�Lm>�qXÊ��c��R�5Ö���lp�;������3o�{H�,�,=�,ĺD%��G�V����K�R�/p���K��i^��¯`����{���:�M�*�P�w�!�D��uMk������h8���8���iG�����5�ZY~��z��M��D�u�7���{�Ǎxu]b�b8�vi<�ح��5@�,MSZ${��bt��(T �6U}��Fk4�w��F����4� �e�˽�`м����l�(&Y���`Xb���b��
�^y;5Y+,����d:nK�L�"�c������X��#CΆ���c��� �l�c��J�d����0�gsR�ֽ���Y�͐�ka���8��Fz�XK����F����,f��������M=>��2�r%|�Iw��l���.AwZ|�IKr}r~Kw����n�嗮���Tb���$�g}v
�
�A�Ռ���讜�C$.�GB���M�?L����`�L��J82�+��7̹��z�ye4�B6��n�H@���P�8D3�0+fܭ����s�^m�8�BͤcObM]���M��F����H�vW�ܫO����>���	I��J~sA��F	fQ��'R���|��b�"�UWg��YW<��Mu�u�X��DE{4�~�j�=�H#��1W qD��ܞ�Jk/��f�jm 0T�%�;a�
��&g��];c�!gQ�
�^�X�"�@F4BӜM���|�C�2,��IO��p�o!����߃X4u�i���r:|!H�(@��(���EΩ�C�1���N����j�L� )0j�IW��7�SBn������"1uj"<4P)�}�;
'<��~��mzdz�JB�\�v�:I�j_瘴=농;��Vef�����"�~��@=�"y\�,ԇ�
�¦V�_c-<��xC`gC�o���Q�G�2�����/!�sM+�����-F���:f8#�^�K�"�w㕄�U�4��9��r'
d䋁� �
4;�
�q�79��;=����������$L@I�����L(IH���b`�hE"��@��%���|�:��7$HL��Rc2��,IuQ��O���ʫ ����>��O�Տ�
Q�W���2WL�B��}6 h��Y�}��H��Qjh��7R�cq&��~��Y�Z[S8*�U�&'k�Gr�rp�D.3��'<ao�j����(g��s��5_T���=D�jAhט���:k�s��6VK�V]g��-kn=�͘jxu(��f�yJ"e�5خ1�{��A��L�R�V�*�d�:�}�u 2��[���D�u,N �alS���\����g��M{6��c�H�O���;�	��%W���rMǓ;������3�N�G3�I8�b�}�`2Z�%i���i�ř:�۔/�B���U��6?��Az��hɘ�vb�M3���~��vL�f�tC��!h�
�z��H��#�#8������v�G�v���e��9��=:Q�j��'#���,�@8m�ĉXIN���6:h����ɩ�٨����!/�ႀ����=����2��@�Y��k%\P�<���>A,يr���F;�J��
�5G�3���C7u�� \\á,[�#�t������U^Ih��xG|-�LS%��Әwy��,�r�8fx��@��bTI���%�M�
�d�oSb� �����V�W�`R������ig�x+׾��j��yJ[�Z j�x/�Vq��E�v��+�]	�Bp=�/�b(S���M�����n#Y|z��V���������`�Y!}����SI7Փ���������Uub&8���˼uK��Zd����w�͈T�)4<s#��<�,p�izs'rx�n�Q�d��1!��$#�'|\���$	��"��;���V�g�>{����m�bV�����"e<�β7B���|/Hb��p�O�m�)~j�v���-9���S i�_Pȕ�i� �nx�	3*��b�����)�-w���&���f����OK���1#)���ڳ��R�[��*%��=�\z���%�So���d$#e��3���iv�8W�3b���)F���\�|E0M�ǃ��	|�k�z�}lzg)%��8��dS��ƞ��Ĥv.�Z���׹U��~�n��)���qҮ3��ٷ�K9U{d*�c��5 "��
���-��p����$O���&;�%`���a�����
��>f�Fjǰ��:h��pQ5��e~.����=�I�0�Mn7���H�{�pt�5x�ȷ�g�Z�E�H	$6}(�tOs:�Qqӟ�[����ӝ"Ώp�*�!$�aZ�6p/���iP�eEh�! �Ʒ�s�Ƅ�:&�uӸ�OC�Y�����n��_��������@��5��I�_a%56��c�L�f�����z8"c]���*Ү��Y8���AsđJ�Ӭ�ME�n��[ �k�Y�q��#s7������5��z��?�Ӥ�q�8G�#F���|��c�.�j6���	�o'����V	p���<�v������Ig���Jx�a�}�o��o�O�?̗'�����>ƯIA��!�D�C�>!x�l@�&�Uhؾ��b~�}~�!s�⡳"��<�2[��E3�)��{%-"(2�/��B=D�R��o�B�qu!��E��#��Lr������wZX�M��N�H��vI�$���Eb+G%i?���0˵`%���$ ` �FN#���"���x�B�T��0�hhB?7��-�->�M-��'7h�;�ħ�rF}6��Dw���:��@tW�9�����F[��@V 'Ag��;lW�j�R2St�tK�E頧G�Kw�_��v����� }��/#�;2p�E{�(|��x�'cթ��pT�}#t�{�."_M�<��^��i��۪��)RϞ�!��+��������Go�u|�:�ML8:z�(9�w��v��,���4�/9¼9��Bs\�dG���g(l���4��o��1�@�lZ3��t��1��t�6� ;�2�~۹W��W�ve>���cdc�j�|�g
L���g'p�p#G�'���;ì���/�M\�ىb�(;[���<��ۛ�$�@_��G[�N}#��&7C�Xh�U�4J�__��-�e }�)l|	}�W��yHnBc[�ܐ��$� )�������4�h�Iv^:�T�
�DHv�n��w'�v�7!)Ng<��x�3�f$ǎ�0�!�%�UVY^D��mt�M�����=+km��F��1q�o�&�v2F.�0��C=��l9����fd|9H�t�G$`n�au��WC���@�Or�ʡۃ� ?Q;*��Љ^�� �,�_�`��~U,Ex���1x�T%�S9�QMA?3���#�AH|����`��2�/o��3��Q3�KHeB��K:�c��n���9��'6_�o`1Y���RX=!��X��icPjS~|��!�w���{}������g��v܋�R�j�ƭ�[h�6�3?�=��-V��FH뭥*� ��U2���}�lǛ����sA����f���C|Đ\R�y�W�ٖ
W���v����b%6�UKu�!-�a�m�@�����W�𧉜����) ^�'P�7s��&{��Ĳ�&�?5��hPj\����=���.��y�ÊL����/������ =ë����� ��Ԇ)�q*�9��Ԇ!�n̩
\���1^r:5��n-[����� �T�`é�Eb��D�{�T��״��f���Ll�\l��UY�����aE��'�GST{&GM�"��c�&���"�c��R	�}�49M��~���Q�q��&��D��V�3W�D��I�q\/&�O��3�D�c�b$�| }g1����������a���=��Q�rx����n~�{H?�B���EVg)�ߐ���*Á�N�	/a@Il����E+�aˮ��-�5�D���0t��oy����ծK�욹1�4�AN���]���0����Ϭʝ�C-�Ng������ ����-���U ��@���\ǥ�MmN��
�m���	�O
�WZ��mv�\��|?l}Ņ�NaC�f�?��F��/s�T�[>R��j���	7"�pmi����Ȋ@ѭ^�ee��آ?����ꕥ�5�&���� ��c�D���U��%c��ʽ��}��щ��X����=���T+B{h���;-�%u�x�ڕ��Q�n)e5 �]����`z����s���Qe��}3�X0a��\K��*�)x�@e0�����2��_��͊�#j:O-��r�k���qjE,F�%|��!N�л��-yw��Q b��ȱ2D�K:�U�9���싱K���#�aw����o�m��0��P���]�t��O�wNe"��
k�����q���n@*�$hw��<�j�$�f�-Р�~`�4ff��k�p�ׂ�j2�E3�9qv�|D�f�k��d�t�g���t��:-N����E{h���͓Q���ng�	ɸ{k[g����JB����jr�Q��;ݥ�J���]3.�=izu?1UO_��E���n=I�4pe�h{�FRW�m���4��ltA�����aqN�V�
���ǲ�vyeQ���u�[�سi�Oxc���U���?�|�?d�� ����>P�N\���o��ԛ58�}�[�4�E��I��Z�䵅����+E9�>t���P�J�J���{��b��Y]|�;V�9�w
	�3`e����Nw�1��r�c�7媆 �s��q��8���#R�����/_�\�4�	�Qx�y)Z���_'B�a�p$Fy�)�ٌ31�������fkp*�d4�Ś6"J�\0U�y�qſ���G5o"�����������P�}'N�VW��U5~���h�>�uQ9h����B�ͮn, ��X��#K.��\��W��o�I<�����VTI��+�u�����ؐN{+��������QV����[�1r'g^�ϻX�YT.Pk#\kG�:�M�3�#�`�[�F<����E��`�O��܀.D���y �1>�K��l��"�&��K�R���=٭	<�_�!�|�	z��\Y�w~�� 5/� �
Y�~�U�3\��v`^�������B>���e�	�%����d�"�V�?^|��"���!��Gj~� �¯E�s	*���V�k�.ݲ�	���ɱ�%��/.�;%DMzFIʿ��N�f4��F���|fV���L�������'�p�O��$����*�U�-��l������n,/{��*$�qM�k����y����-/�����#ۃ���llQp����(��'��F�΁3��!v?,5Y�'��J��Kw��(낍���T����w�%�5v�M�_X� �5N�8��)���4G��-Ĕ��2�����D�Pڋ��b�J��F�-���R���α�,ע@�*ģ���"�+ZKЗ(xL����es]��#�#C�
��P�4��-��_�ZAT�ٟ��*��f|����OC邰Y���R�vM����,��x/�f(1�ׅv�H�X��:}:�D��C�x-.��P��1��Bη9�'q� K���q;��O���p��Ƒ����D�4e7"�#X�r'�E'wg-4���pIxY��^�v.t�^+����>���(z�"��[XpV�r���P"��k��3�=	�R�v] �&2{���my����⣒]�T!��RC|Xa�Q�WE�!ed��ǥ�Oq�l�16�oz�OAǙ���Co�����b��r�6�+y؟�k��&�+Q?%z��'��>��L���J�I�p�y�|� )���Cs�g�j<���*�XH��O{e�&�g������'T��%"�:FRJ�3a��wb|�)���'�:	ʸ��Z�*)���a��~��?Q˽郓��C-��ƽ� �}�d���"�음�n�)��.�ѥ�:�Q��Nف�ۜ�	�853��De�e]�I�|jDy�؄��_L�����.炦ӐuU�m�S��O�g|�)
����[�/!��с�\���G�<Ja&O�oU�#j�U�?`A���E��hz% ,�9�~�]b]v~yv`�p�t���_����	�0z�Iy\B�;U�/3�����Nԯڜ뢲#x��R�O_���kc�}�<<��F�*�;K4�?x;�pa(
5���r:>�/���{
��]5h�eϋ)6e�ov�(j(�5�w�Y��^;�^�i1p��Τ�+����v�}��*�,w^
�������0�Vݿ������b�ǧ��� %$S�hN�QF;?�X_��'t���Mw�I�'��@`a���'@ (��̟jy����(�
����5��]&�Q���:�Z
X�e|�H����-	��XK���؂�ɀ�FP, �U��7��R�S������]:�#�D;�ϒ.�E��!��Dcr0�Zd� P�W�N���_������ȭx�9 Ժ�D�R�z�Йt����=��@@#8�6��9'MJo�y�s'/C��٨�Z=k!)��I������^X�m�2�<��\����f�P��Rn�c���)$`�d�G�h�m����Hٙ�3�_ޡ�T	e/���wMN�p�S�l�?ez�*��tE�%OȑGB�x��� ����e�N�HA��wN�6��$�<�%y�߲�"����	��YB��� ��j8r2S?�:��S���S��8��}��i:��EO�ѾY;U1�8Џ�%ͧ����Q��HYI���J|=w�lK��!#�ɱğ��};cL��DD�_�\=�/�B�e��n�K)�--���h��w9����%k�+T�	�Ҍ4C+�F���T)�Ĵ"�Z��<ڶ���x�fa�J�̕筕�7�����2��@�w��=��Wx�mr���f�#?�>��f��p=�~�h�P�K��Kz�>ך�A�K$��e) 1-�d��^ �'��
��?j��)�CoZX�'K	\צ�d�L�I+�wg��� n��h@ �	��Jz�l��'y8|��h^��XƗ��D{�'�`�߱�/q���W,hs��On��E�
���eS���+Oߦ9k �G�8Cǟ���#9�	mt�_��=��m�6ݕ�}�~����ǶGM��֕�̴I�{��o/B_�g��d&���g7��ԑ�l�9eE�F:ɍ���}��,���s�͆~���H��a��Ĥ����t�h��x�C�^]��=Nm�Ly{���/��q3g²��zn��𽊣"���3�v9$�����7h��Uz08A�J��?�~����>̞2�L�p����9�y�,B̤�^�sc��U̽����.	�1���U�G8�Mw�ql�!g#��D���aE�j�u<
`���#|�ï������6U��e�dվ�u������1���0͂�ҷt�H���3�����FB��;:4�ۦ�0��⧯�C��#�+h��W�U�Ё& t't,6U��Rk��l�?��ű���43��Ie�ڎ������Zgc�O�����j�	ʠ��8���x�	��ZQlb���
bп�o�k�����\�E�$����&#f����X���At�r�}g�5� �8�=�=�+lO�n�3���T$����Ʉ��c,���
A1d�ӭ����d�s����I�k��p�����|��.�q�
���iD��>�����P����j�N������9O�2�i� V���~�- ��c����+`E�4ی�kσԌ�r$�K6�:o>��ӵH#)�0r��β�|zw���K�����~���w��u�T����[���mX�l)��] 0��w[b2�Ⱦ�xǡ���4%��jX���K:t����B��3v��� �e�_��[Қ�`�����y\}?�W,�X��tp�7���5nXpd]�=]����~6dkT��"�p��Ϯ���H=;#fz7�q"V=����D��y^`gnR���iXh�gs�=�
�uf��ԉ�ׇ���v�̡RG���B��}Rdn��ER=����`Ŵ�5g, :��zmRY�Y�wEY?
�c���ԙ���[̼�]��?��sT����3��Pi�� 6�Q���Dm�ܿ�e�f�N<b���V�3<�	 }[�J���8-B�f��ļ�f�뤓R�#��N�U��P5�Ո�L�?j�G!V�5wo��Ř�KT �I]�l�q��k�;ӌs�H���Gܬ��ta0��wGh�!3'�*��u�QEQ�)e^����|t�늋���x'�Jb��!� *�����d
 ���	<�hnM��,�;0Ε.�\�����"�CP�|O����0!�d�W�K��8�X�y�s��zg�_��Λi	8��9�G��Ж��H��ݜ�����_T(�{���t}��:&N����2np��Q�ݺJ��$bC�X�<c3���ѿܤs��^ք̿p�]��m�Px�N�v��8o���4:�GS&o�!Ӊ/|Ym���̞1�K�u���BNm����<x���w�&���7(����x{J�2G���+�f�tE!>�^D�.yCmO���Da�p�@�(-As�P� Mգ�A9�����U�պ��24��ت��%��$i'�6�t� !.�F��1
�oQ���
���iu�*ă���&�D��� ���,���zNm9=lO�?�H�>��<�1R-;�oN����H�)0�J>���
�Ŵ�q�2	�T|)_߉��� H=��:�$��9R��т<?d��.!8��Y&�p�Ѧ8�#2�ܪ"M`Q��D`v��
-}m0�/�;[%Gp����Bd�]����d��������yo[��'��bi�0�k�,�>��I?�qڒ����8�E��u��2�BO�U��n��m�U�����L��m�S�����5�c��+W���X����.-�[9+�O|�~i��>F ��^�h&$��7BŇ�h~j��t�³T����. ���p�.;�M&��|`����V�Sb�~��r��:&o��$(F�wY4PBNN�G�Äb�C3��������k�q`�� O��E�����@�@Tu
�;��<K�
ⵎ��\6�n: ��<ǘ(��q�U5�c�0Nӷe��FQ��w���*A�>��b�ȡ��ja�ν&'��#��"]�=��U� �ِ��W�Ģ���ү6�	�t�f�Z�I�U��[K���a�+譡)�y| �	��Ѳhh��z�H��S (��q�.#��S���/(��6��&As:!�I��@��V�R�pir]U7Y`G�xkߐ�������&�E#J��欿��?G}�v��љ��R�؊)�@��M	�۬�`Ħ������@G��P,�zep�OB�5���哴���+=."v���1 6I��|R�Lk��76M��2arCA06��M�x�G�O��g�9�5�Op)��\٫�Q��?�/ya��S��X�ͱ�1��jk<.~�b��-�a	ח�qjx �9�z$���	�g��� r�c�6��b�:`Lg�d��˯\��X�^�!�p
--��ڔE� �n�fv\�~�m5�B��.[���&��t������S�z�S��l�N&�E]��DA�i��s�`
ń�<>�}���$����g��Z("\�JH`���*J0 �9+T�N�R�/���'�uf����З�z�ÀH�+���9j��Q��0bqm�s���	1����*��z�V��ߣwm�Z����1�x/V��ʿj,L��v���)�- r21s=&�K@��6x\��i��he���y!ށ�J���Ϋ�|��հ@&�"�x��-��+��G���Ni�R6	v�� �����B���:�Ο���4(.������$�@:�zXj�`�ſ|�s]�p�JB�C��yMv*8��֏N�O��r�R����7`* B6�w<&�K!����0�(�	t�Kv��B_F(���mb��V�v�^3Ι#<
K*�ꡪ�B�'�^G��%u�NsbWYT ��͖Q.�¬h�)u4j
�KTI�D�D?�����5Bo36m�QFϲ�Q�����wCX�my�"�.b̶�U�W���*g�K�ٞ��>��:� �G�o��<�Y}�}��q6(�o-�$��Ą7D�a�{�a�H�2.AM(����5s�H&�!��U��(ܜ�I�����=-8�7*a��=���lyd�C�Ny���A�"]c�E����W-+mzz�X �{��Ҟ�����" �`�&�:S#K������@��$��OO�t�k��	�
�T� 8�˴�
Qz��ɽ*_xO�TQqn�ră���oLio��mů��B2kۑ#����>��ط@��*��,Z�J� ���t����X��X�NL\�n�Q�_�Z��T��e�`�&��I^�� �/��r���n"���}�xh�9��A��8�W�y��ES�<�c��@�2Y��������/P�c
�Į@F�T�T��ܰ�V���P���Z�X=Iո��ڃ2�`�"n6G���I�CS1�~���T����3�jA���̮�5���IN�ɬp��K �R�+�����G��iU^ �BH��'�ȑ�x�D��E�t��,��r���L�g!1�,��k�ǳD�&�qc��Q]�Ê�Ȳ0�#6�>H�M`��Q`�x~Iy�\r�Y���,S�Y]ITQ�l�,YI{�C�@=�{Q�	n�K����)ȋ̐s�����5!�VK����Lì�{�JZ��5A]�{�f��݁ꤿj���}��Fr��bY�t����s9WF��Y�c��7���$���Rk���R��δؤ�x�� Da@�Bi��^ѽ�g9Z8��R�F�����W��Ņ���%�RW�;��L��`�`��>���Z$�.�j�ۀ��4�&ST���!H��4�סL����.h���O����[����S2�׵&;΀�Q+��t*��\5Z���2x{_@W�q�h%�-i7��L�5�-��̓�_�B�A�V�'8c���Fr7~'��S��T��Y�}��C\���@flNX�P���d�֯�hɎ�x�y�^�����x�8.���J^�{���[$�%�]�,C~	â�~$��&�3ڦ���*��h�%��?&��f��̆���T���F\H�]\����쾰�v1�_*|p����H�0��p���mgp\[�x&V6K=c�t�c�#n��/_�'Ꮿ�_���W�-�M�����]�%��/<>h�$X��u�g$��;v�}]-e%r�ۑ���٣"����Q�l�ifX��o�t���9�Z�H�$}W�ǳNRQB��zZ���7ۘ9?�X�9aR��r��'&'d��J�ui7?��ac�Ob�T��z
�Ψ�HZ�����Bl���y�{=���*N�o�)>�%r���]��c��U�~R�W�e���g��	�Eo�<�*!��1/�	[�%�麯�6�w^6����S	&�ߧ�e`�J|�"%=Ů���{���IH "2D��*wu՗��b\p���A,�y��)�(��ݱ��e5 �/��p��<t�/i5� 8��kzBch��9 Dl�Ϥf��:�x�0��8�]dHKSu��OD5��n�{��3��i���A���i(�68�
.6C!X�G��AH��?�Y\�t����,<k&�֛A�-�&����t̾'�t�R�$�H:?"׬x��`�� ڗ�	�����khכ�%�D�n�xW@�ǆ��M���
Z��f�{G� ��]twR�"�,�ԀL���6=�b���_�ӽƧ���=��/~�{B?,�K׼��=��#)�yHTP�Ġ]X��gҺD6$4QM^Wi�_ e���L/�a�On^��7�����Yl�vH�j��y1U�>|��p<>8�b���-a��瀝፭$�&���ǉ�� �C�p+��b�Փ�M��Ȁ�8ֵ��j��Y&�N�Mj�O	��ኅ�|�g��cEc� �FŔf������L.�H��
7�w��l��f����}��k0WmLn&�.�h��\]A�>���Xl���H��� ����(_5�9]��k�<���@8O�qjy GU<=�=�<�'�6��4���tu.^�(F��.R� ��d;y�HG{f�J�!�A��(>y(um�L AJ��oM_��z�����A#8c��y����&�"v8u�~��}A������($83�)g�Q^�ndFW�#��4&ْ[�}�[� ߭F#Ke�g=BG2���������rٸ��*Ye��,+G�'2�E�Θ%Xj�LЮZ_�!w�$$�XN��BDuE?x|%�P��o'�ܸ��&篱p3ԣ���1{V�|�P+��`����Q\7WP�"kuE�yf�[�"8��͠e��:F�c��'�DjJ	¨��� �Ӛ_xW!�r�[���*�"Ǚ��d�vo�l[4e=�8�_H�I��=9��m� Va�>��A�S�������Vk�<\�wc)�]���04�[x���f��u�9��KdĄHD;j����y�nXP���"`�5�HQf̒t᠘uN^��@>�L/@���^�����	�XQ&�=���\�y�ƌ}��L��U��u�6���F�^��	[03���һv�4��v�I��q�sfÆ�H�hr[��b�!��5�ڊ��":�+�E!� u���6<(G�/.\2ڑٲ��MrI<�Zi�a�[L�� ��UFv�h_i��٠HFu���(�#+�9�Q��� su?����V�F�-��� 
A��e]5
�T���S��4Dr�km��͔ dγ-���l	80uyG���R�$/��"�*2��;�K�K��7C5�����-�NB	ۏ*'@yi��ø�#�!�>0/*��sH�^��Lw���w�3X�,^4t$���C?m-٩$%�3� 9�x�W�۫�GMs�3Q��
�?�Oؖ5�&Ӊ�3t�Olx��,������- !�x(\F���~%qݵ��w��\Y�V�B=^\�,m��!	�벝�����U�Ĥ��ފ��Ӟ_k:���cSM0kٻ�>���S���톌6)�R"�+/�������P�L�}��6�酑�5���6�$���l榤�U�֍����gS�1�s��o�
�,��I��|k�B��V�}nG��P�~��!�CsFe�C@����GEΞ����y�+L+�K��4Ͽ�B		�1�7�\��c����p�8^��#�KZyM�s�K�m�CG�ZhMnd�gZe������T�Fߟ�S� U�_�O�<ݪ �*�y��q�NSN�粤���:�:�����3
��-�s�I�۹�{�!ß�D��πZ)MD���4)���Z{GX��YX���i��]
�ru}��S��f�k�A�E�5�
�Ż�E�+ဢ#8G#�\��Gk�cEb������,#�w�[S*�1��2�~%��ڦ���t� �޾��&�Iy�F�V����m3ӗDRd�*�bY+�@h��֚)4E�)�_U����[T.m��^����]�����rSZ�Uj�������/})�#�l��4���n��u��E��}	m)� ͨ�ۈ�-s	�����yS(I�=�u�X ��ϮI>�2�Y[�]��v�ٰ�͐/w�Z�h��p^E$]�S|��g-��sYfΙ߸�
")�N��/��%��i�	�aL��j)���g�R� ��ݏ<��ǂQ��v�������MG�78Ǡ�~�.�0��e�
f��ǹq��>�o�T��l�PE�@�Sٮ�Z��N����,gr���{�q�a����vF�>�����ԇC��lR���QJw��]�ʢ3��h�d���������O�u�0�Av�Ⱦ,��O���y���(^�PU�:�_R9-di�e4���~l��fk��2�j:��Kh`�
��6���F���՘@w��a�!^����3��2e��TȽԆRH�iKQ�W�V��$3�j�l��\����dn77�ghO8���Kd���~r��s�5A�9�<��c�D����<�}
�޴6�Y�Z��(п���0�T�����0�-�&����2�;�Pݖ��q�ͦ_��6�4$��wh����`���}��V�޾j-�{��������2�4�+�c�Ό3Y� W,�<8̴b$$�Qyi���<�ZZ�{TqР����e�qp� �L�j����"�,TG�I��v��7Yݦ�-D��[Q�+��A6�V�q������T���4��ֲ��d��s*�&n��gn�[�44�AK���Rî���0�,�ʀ������50���/Zʧ� �w/�5�������0��ڈ��>��>�S���"3���N�m�$b�$[�ai�N��uR唭��|��`6�]����WA�Ų��Nu}m�H���|�_M��M��U.�m�_0�{����o���..%p��� ��df�gr'x�)INX�c+çu��Q�Y�8�>�qs�2/e���O�.?S�'O�V��֋pga���H���~$C�Z"(5�K���L@;a����*t�	؎y��)T�8����[�j��� w�j1p`֫
���Z�e�䓜sl�1�e�>��[�L/�<1�B�A��8J盝��(V|�g|P�k��A�ߺ$�[MJ�]8|��C�[�
-���BC�:�s�xߪm�m}2O4����R��T���e��Z��raG!��a�[/4�]�Z�T�+Z��$��uq��	k ?�q6vr��X�Ɛle�u�N.(�/NZOh�g�!�}V���C��J����]�_@^}��� |����7HT�3��8Kt�_����r0�Ї~k��|]��Oy���7JiQs�9{�6�z��)��S&n�[���A�{��璊�ܢm���eP��c�h');ڟ87p"�G_u��F8��8���qOD�(yyU{A���8�wJ��DX�4z0;}v��<���]6�~�/��FvMc88�>�ze?�E��%��8ă�T� }W�lo�tHqV���c��9�Z�o���cC$���]���ެ.y�.��-k�D�X�ڪ��l �)����2��I^�Կ�+t�6�@w���X��϶���i~��?�ԯ��բ%
M���#fAA�ȼp��%[�u^���ZT ���LʷF=��kl��s�a��ri�k:�[���Z�k��a�>BD�%`�C��]e���Lyzʡ�,:���<�k�	�BJF��
�I��3}c�(�;.2[��k!y�~��m��Rc��*?xU�Է���t����7�J_-��u�ъ~�	+\��$"4��|}����m��*������0�IL/3q�G�0_z©�Ћ��k����"�,5S4��L�^������l`݆�� �:�%��4�=���S��:�UI]i�"�3���҅g[� n�zeX����th��������9����;���ȭ����亵n��%�"�G|s�I5V�?�V��N��}���8k|B�h�^��NmxF��0L�­��e6�`J�$���"N1���Vc��.x�#�~�����z�4.�>���w�0|�)�K�����g�80:�ڀy������	O���F2�+�L��ݹ)a$�6`�;��������Vޒrx�sr+#��r��[N/�,�̘��X�;�!�;��ۀ#�[@�`���oe��Yh1�ϊ����@��|Ȟ����~�\�w�D�?�/�w!���cG#�I��Lt��:��= ���Jm��УI3WoGJ���}�ȗ�wq��I��e=�ݹGی�>=�ZV�w_@y_r+�.޵�*)�s�
��_��&7i��#�M�F����R0L������'by��������
�2~i
T���4f����1 �cwһ<��t,_c�g(�DH.f�1�.�:	�k�BPW�[�+����S����Ҏ��6Y���1����"�����V��� :/-�WmU��O�8�=|��N8��]Θn(Ͳt���,���L2���_���:�q`/j.\��k��/��=#V�4�k�=��C��+'D�\�ϰm�y*��z��#���[�#w���(�?V�Ao;�L��AO�E��I�ݚȚx�Nұ(R=I^�+(Bs��
������Z����al��]]+�p}���WLR��(4�w�<۪w�~;w�FDr:�U9��/![{�7�pк�[�A�1���A �	}6~v˝�e'��.Bua�#�x��-�^�����H�AC�g�/��G���8f�M#�X��@E�Ee��XB����7v�^�6�Ne��u �O���E�i���;l�nݡ�=�-��z+��6�a�]�v� r�rqi���>g�39֩dvA~�="� ��]E)M �AFk\��lh����΂4kIBrx$���U\��[�"�}�-�x��r��0�2���fp�W�r�*m�Q����D�p�4$Y���Kݲ�����	TA�$&�|N����R5�Z�	��N�8�D��z���Q��hU��0���m�3��9�ְ�H�;MX	��/�CCAt�r���j�!�c��Љ�/q�����Y�t��V(�!�B�.M�\I�?0=��`�)�a�ƻz��O�p���N�bbu9�����J 9�E��-�>a�)�-��z�a�Dl���C��_���~��{g[��O*1x�~w�1h΂��,�� � v���~���bA��H �0��:�,q=����P�zv�/{k��r��W�!�1:���[#�5�P��NĤS�H�v5`����s�ݑ����x*K���d�:�R��b�)ꝁ\�W��~8��w�4��@����M'�Q+>���oaǽI����ƌVz:�[>u/�NLL�J*�\KW�"�r��;��k��q{�j��a\�!���x����t���6 @���8\X+�\j�=�Hel��S�if���{��^L[Db�X��5��.Y��
�^u�4\z��R�3��~��`h���M��RJ��A�#ւ��:�C�ͯ�\I���ؔ����"C�l�L�̥��Ү�[�W�)@�q�|�zc���.C���{ji?۴�3T��>�% '��O�L�>W��0 )�^�L��^���I�FEH��;�}1�7����/U�C���O�[3F*�7>uy
 �o1��95&"kF��d}=���-q������*)��f�Ɔ.8rr^����X'�^wj9sN>/k*���z"y���Ś���� ([�PZ��x��И��pGp}}��ӯ��m� }�8U\,Y��})Cre�Ң�(�ɜ8�W�4�8ZQ� ��)\�(2���Ӕj�c����n�$Fg뎠���d��M�sa�>��]��JR�/�����Z7�F3,�U�|<�����>��= r
�j]Φ�oBWk�sc����H�
���(:Xo:�(;�r��A����/q����Y3�J�^vp?ER�Ņ����E�$)�ȯ��n�'%��"s��"���ޗ�㩸�<�N��K�\Y��K����ȗ�;V�e5�Nz	�>a=9~��y���*sd[ȑf^������=���!H������w��NC�8K�e�n������J�����#����)�"q,N��q5��	4��y�ۋ6|r�O#��b��o K#D-��	H��Z�6���L������_�z��ڣOŷ�b{�V�{
�ø݁G��Gѝ�����N��� �P��lU�܍o��b�Jl�J��1�u۽�^;�򊿀�k�)��굊t��M6�G����[�q$x�D�N'�W~x�~15f�rŀH����;�f��Qʚ#�e[~��O�Hm5�%du������3�uNB����Ԓ�|�'�t��&QM:�7�J��ehz|��h��l�m�)}C9��7@ۦ~��k>J�R�i$z��ޞ+��њˋ�f}�;�b��d��vX]��Au�F�s�5���ݟ�|aI	7�}�9V��.�$v��P�.����|��\{(�;ӎU��~"��+0�<�+��;?͠Z.�"5�$p�RBǀ<m̞�Cb0�����gm���U��&�\X$9�9|c�hz�Y���L5?��C�<c��'��1���W�|lI��z���H�[�C�r��∮��ſ*%��)PI	I!3�>Mc�=w�E���܍�gT�e�[�f$$�5��k�'�c���#1ן|�W�VQ��k^�-�-5f⩎�`�o'�>�l`�|v$%%'�㹑��H6������:�QF�z'�3�cb8�MQ�Z&�k���2@�Xӱ�΅3?A,FO�D �~{�-�c���W'��]O��1�3�ǩ���\����Ņ��Aæ�M���]y��s���K�z���ӽL���g�ԑj�o<wH�{$&"]IVGR��+)�Q%���U��BS"}Gv2Ķ�0�2ண���v~W~[>>���ߐ�_ (��ɖG�]s�
1�>��E'�r��v"�Q�%J�Vi֟H�t�O~g�?���v��y1�l����zy�O�a�DG��V �i�&�ײ���4��`�X��;�q�V[A��U�O�-h+PE�E�5ʩ��зا6?X�/��^ɮP;�v:��͗p{��؄5H�,F�b_�n}�AT��B4���s�ۥB,�"��q˭[�h��_UHxT�Ȝ-Y�N�ï����EeL�����'@$P�$��_���a��ņ{F��j�*��N��+?���3�=v�
*�`㧞�8Q�C7C'�}4���?,���j�S"���5�o*�.�3i���V:H����v��6�������eM&�IP.7�.%d7�m.ꭓ�P%���+����bZ�؇�'��kϳ��Ea�?0��XIo��N��xZJ��H?�JZL�H���|���M%5!A�*�����=˻{��0��+�hK\I��i���J�����{(no�n�X�G��X�M���&���z�7b��66�v������;��x��j�^�x����~Z5h>w���@���:�l2��ׄ*��h�e��G�{��|�;���i\t^���P��-�g3w7�-�ϔ%���M�=�T�7�����������b����YP���7�LS6����%�KWӒ�d&\Lڿ6�M�x�*�ޣ�����s4��;���{\�V��)�>��z{��<.�I���l����3?mCp�y�$�p���������~d��ʰ�"��t�`�'ϧB���'���	ߑvŹNfQ�׺&��ZtLr�����Q����'@�T�f�[�_�b����c�� �|Q��{s��Q�ۆ���]�+s/L&�"W�?�=y�!7UsŢ���@m�����!�d�Ǒ��l�FK��3�ږ��oy���xu$��tD�~"����WTJ_��v�G桏I�C�M���\�O�Đ�z�[�?��6�h�@�w�D�@�������i�H�tT3g�K��J�0#�g�j��� �	����Jؒ֎Y��� �Еsm�r
k��$1"'�	�Z늤�Y�r	m�՚JHnn^E�i	~U$��
�/e>rrư�v��=W:X���~��J* �dD0˓B<Q*���餐��H�uB��Ԝ�@�a��4�#|8�!Ig1�y�(B�7�0�8؈��{OzW��m'��yN2�
��#U^���b����"&[y:�E	��'e�ԟc	����V�צ��Sd�G�1�@�r��7<�$Viq1��G�2d��9��.��d�A׌�WA���`9r� �}��������-��O�T2��7��Gȧ|]�<j�c+�4
7��ǂ;J�E�O�����{�wG��Q#Ɨ�Q�THӁ�f7b�c�h�Q��u�sĊ[����p5�����=���d��4�.0��
���x;��2��j!rl�S��q�y 燱"�&N��f'�@KN7��\d���V{	#}�o�P��@P�F��گ��O���-|,{aP���S�A�e������2E����l5^�F���� 9? �tNlb����m~��m(�F�x���1ب�/)���X����W�L��Kk���}]�V�=���wh�f气�-uD���1g������t�I(#���^����LdJ�&��Ct'��#P��#��n����*�D.��L�X$���������+��Pb�{g4��K�Ba��8p��]�pS�0����L���$6�N>�~$�3�߸�>i�{a���	����9'���`�`������}O��"�\������s.8Ԧ�:���!�x�,�<)����|����4����M?q&�ؓ�5z�>;S��_�r��IS%W4	�(�2�++v�8��/����ԯ��/u���8Mx�R�g�C����O�~���H|����k<�)$����*ԺW���gS�s��w�E��ڟW�z��B|V�AGÖ�;ؖR�	�[6�I�Q��!���}:�J�`mDkz�u�-(浏�[}TZ����G��豈��{A�X�>H�U4�V�w'�`���0|�K�VO,Z�T.��+�:G$�d� ��!����賦v��3{Ͼ㸐�7�(��t����x�f�ePU�}���KmlY>|������(k��)��#�6��X���4�x�jq�@%�Ǎ�Z��~|��B���ه?���q�?ÑL<��gЮ���z�:��E��v�:�[>!���_�,$5�N�ߵ+�1bJⷱ���D�L�#���ϦX��?�Y�v����s�BZIl�?+��{OF&ly�t�:[	
�����Wأ���)sg�,m�K����h�GK7�(n%�~�k���o��*�z��u�Lꠏ0qF�C8�}jI�;����{G��x$v���	O1Ŧ0���An��q�fI����p+�\-��Ew$�������$�^0I�����Yf�f�6�HP^�W;d�D4����x����dY�� 2|%U�׊�LTS�d����V��ID1Il����b�'$B�Ш�0�D�ռ��)�U	�>ڢ����K��2�>�D���k0Sg�:)Y+c ~3sg�K���p�Q5U鈔2���ș�xކI����o��8��Z�ڣ��G�XW�����U��)�e��N)i1CV�=8�O��HC9�L�5O���(����|��)��j��Gi�y���qk���dz}3]�_RJ����%Ie�V6.Ԫ��9��`�9Z�����	�[Ӎ�?(�Xuy
�z,�άD���Q�s/s~����2�Î@W���&��g%6�2��0�ny�u�S(#�nU?�pܫ����7G�Єݺq����/1ĵ���g.�L�q7-�����A�6�um��'��6d�vŇ:#��>�`�0�=�aŘ��I���R8Λ��P0�6%��n�����P�Y��9����l��9M�G~����Ǥ�C2r+B��P�4�!�ķ]��֡��c���D�vpk�U��?� �8�q~��7sNx�-K�`��|3�<}��SA�JT���3g��
���~2h����v�]�2Yls��\=���>Zd�DP�8*L5Y���ւ97;pwP���n�eۻZ4�2b�BRI7RK�D�H����KW�-r��x��V:ȗ.��yi^��VЧxj\�t�유���#e��rgt�o�y�
���#~|�FاL\�1�ገ|������	M�"OXX��Dx��r�$]��j��&T�G��'��+q*�5s�^�k7xZ�++�B�J�8����w�~�����"����
דլ�S@�h\�;�0��d 6g���)1�L�a�%��>��,�I-��,+�:�1�U�eVoe"q�C3ג&�[� Ǟ�p�,�ڳ�6>$A�Ɔ6�<'�����G�'d��USgk���W�������7(P���P��蜂aL8<�'������w��_[�h�=q� w<w�j�$��(�#��5�u�@�(G鴞��C'CF��D�ϔ��"S�:�r=D[��P��f�h`|�3<�Ή����ᢏ�!.�A�񽼇�G���Y>m��\�A��T4Xr3J���e�6�ك!茾�_2~��8��QhP��S��8�-Hy���|���]T�'�Ҟ��A���o��@ˮ,JK7n�dcp!�4{�9��$���g0��P!:!�Z�'����~}!��
�$w�"���ܝ���0u�cD�hk�G��S�]�#���Z@���W *vp9�t*���ӻK�^YET`֑��8��y�8�#���:����4(���N8ܯ۔�J���������*�2��p�}`���6�e�6�ʳp�����g��M^�x�6�V��1Y��4�{���R3�V��'#�Ld��x��DP�|�����@�|������m�(�y�}�t�=t˗�s�:+��°YnV$�h ���P���X���RE ��~7z�8:^Kb���-'q~�b� G�K�J @Y�m�[�]��$H6��x�s��ɚ]O� ?�)[�np�2k��H���P׺LF�.P�$)�b��ǉfx�����i���x�d���5
atC�N�$�n������@�����`��b���9�LZ� �(a�j���ůa;�A$��F��ݯl��A�KE�3�p��ɒ� Fg��������)MA~�{r�8a�᯿��w�9��lw ����TE׿������pË�QgB${Q��r�VF��3/��lVe��:�Y H,�m��ӫl��cUn�(��S!N�+��f�5�%C��&��NǤ�g���`n׬,K���;�]nLA6��T�
t�����z0fH��ݛ��T��2��$46�k��A��v�!�[�d�E�#p#uf�]%�:m���(�/��y������2���s���ʌ�Om��j'^�a����.��҂/j�'4lXgk����
�ɹ2Ò��I���:�G�m'X�5�n�֍��f8�/5��@/��L�����qĐX���i���b���`����"N��ΐ����y�!*pr�ҟd#�P y����0d�U��2��a�Ņ%�a�h��{���3v**��
0K���ݍ���[O��yS�_Z�}A��w`��EQ
��d@���M�vU�9�m�������^NM�����|L���G�X��^�����Q?8c]���C�[��5lC9-��Y'=��g]�^(��:�_G!�Rf'gv�U�nfזQRk�����a���FB��a��k�Z2�^��<n�5M'�p>�̛,+��A$�VWƖ��Cc�]sI�İ'F�q�	��e�|Um��z�	i�$����o_^G��L��6	Q�΍�	j����?h.T��%`�A��>�BBr�8K���c��*����?J�.�s�জt7u��7�`mG�ܓ��/;��M��}��aǡyH�b�9�[�޸���J��~��Jx8��R �����r�I��>�St�.X���ƿǀK?���k��Vص�r��q	�ŧ-�VI[�7M1L�b�ze�,ɲ�����d�QV/�lRe%��&2��!�duj�L�(���:J&(�jO�X��5���I��J��kvɮ7�eW��[P�6��-��U'X30֨3	4I~���܅���F�m������(�Ȗ^�&~~�$�?��; �_�����/�q��ny"ѧ�6�0[�W��5��:�'��?����2�Ǫ������%���&^P���ҷ�	���5�S��3enU5[�so�-�,�`�s�Cf�E�>ƹ����P8@�U� �,_cA�(�m�J�FK��,}����	7�ܒt�
V����@���«A>�'�J��)�D1����&m�Y?v��ܖ#���l�?T�g�&[��^%ړ��fA/W�4|H-B	!)�ۚ���x�?(bhL34dFb����Ke��\uz�T�!���t9���Hg��B�+�'A��"���>�3�&;�#��	Jp^��̙�-�n?� ah|�+���;��@��T;��Y�Z|f�i{a���"o�7`��-?	��T�z�K�(F�y��8u�¬�y[�z"�pQ���lRX���ԧ�Og_`�n���sqd"���FϦ$�zL4m�G�e@/S�ߢ5���R�-�RU�U��9���9�}�+kߙ?����e�,��|)s_�/�!ASw��o!�*�D�0�j3=}͎�W�=��t��"ᐽo,��% ���ɟV1 �㿦��rj3��]��g4X�jd��%�=���Հ�,�JKX:H��/^l���QG��E���ݴ&::���BGCH�!zaB�|�zL<	�;k�i��g����S�pw=����R�|4eWn�Z�D��~U�]P[-�͓!�G�X%�{��^,�������z�4�p��a���#���R6Z�v���LЪ6��F�7��/��Y��b��S/6n� >�c(�u�� 4��S9-0��6}�[�,�����p�|H��P����/��5��e��~v�1��_����*��EO��[ź��Ɠ}wm߰��X�`��zM��E���5�^UC2�^�C�`�����k2��E ���=ZA6����ih"�t{tV��wgڴ�̱��W���TI��~�H�~�o��q�y�+Y�>U[�)��C�y(__�*|m1E�4O׹/'���ėM.j�^@���#ǰ��<�Π�Z���W��a���E�E�壠��V�����mE������s�.j�*��:~Al3*�dD�W�$)�@��gt��,Mͦ�� ��µ�?�7KI)&㚃!�D�yd�H��F��������練}��!Hg+i�Tl��^ʏd�#l6��Ξk*a����V�Ɩ$߬�>2�t(7�+�`E��G}l��oc��4Nܬ��/�m���PI�m��G� cD+�1�g"7l����U��>��P��Ar\y� (�b� ��e�X�J*Gw�a���K�6KQO��u���v:�,�Y�Z����-���v=N�i�w�[T��hAR�9�� ��������N��}r�?W�e��$eH����KR˝���V�=P��:���O�̋;�O��!�!8&��"ǒ������,��靉7��Y�� RX||9�U����?����5ĩw�s��%������j�r۳�j�1Ϲ&\�5�u:*���@9piX;D���x?��WO��/?��ly��I�����1j<\�e"Q-���"��G����6�,�)���k��f�^01]�B�.y��΅c�g��VV�Ek������"��4�Ɩཛྷ�
DZ��?Ԏl�9��ʘ�F��玩�q�2���LHOR0p7l�K78�6����o��ƾ�2@��a�A�}A�Ѕ!�����I�TKK���w��տ��9�sǿ�p��̶�#g�UK�<�	v��{�Y����� ���̋
�9�$��J2�r%������r�
����$n��溫z�	����F,����e����J�[���K���s]Y�Ggq�2�73(��ɝ��\�?0!�DC9.��
��^K���f��].��%�c���Kv�����Q�z?�喼��+fS�z���oB?�;�%���9�m͝�v�O��qi`�X�!&~E"&h��,��Gmg�BҴ��m�Z)G2��"��\�#*�%��O2������2�_������[d��D,�RRX̛st	@;>!�{BBY�b\a����f;�B�
ē���l=�����P0bl
�y���5mq9��,a��AB�K��������p����+�����FHؕ@e�O{Dx#���U��9���͖�z��m�,xw�|�_hǺo�5�2:-�Tsp�sAVݦ�ú�����a��F28��L�`����58�H*��of�����8�c���UbCg�����f�boG|7���Pw�)(8���%�5�˾���<�,�E��9%��R��W�^5��V�!'�!ߟ�9���Tg��,�O9�5Aݰ�!�F�Sڬj{���?E�����\��&̊��ܿs�W��]{���w¤X6���\%��vHP	��%,?:�UI8!Y�0ʚI+%�w/�֪����=��zO�y��@>�Tݷ���3�yы8�JD��Է����&.�-���wt��	+�m ec4��nh�l��a�K��O-I�J��U��l\�'�b��ay;, jfi�d����ì���	���.7�`f�Q$�p�34ܦx�#��(�y� .Y�A,^(6��yg�Ѽ�m��#�<��{'�*
h37�/�i���ҹa+8�B\X�T6�ɽj|]�$�����5W�#�ԯ��1ט͑��X��z��9&�/��۲��	�b���4%
��P���F�
Cx�.�B�?���[��[�/��mF2��p`-\��6( #�vOTu��F��B.��ά�d�rH^.k�Z�BD�M����j�B�2�h��,�hgNakٙ2��f�����6&�
Np8��{�'	�d8�zC�p���J���ڍbW,��E�D���'�[����m�>8��Ŭ��,ޖ�^��]�mw$�P����w�y�em���ا�!��g#T����[����W'�a 0!�}�½��U�\���-�u��p�R�*��l=z����0�y��r-ۺ�ώ�$T�gg�����{�z��}�1��6ӹךgԥX�׽��0�-����˫����I���~2�ƒ���a��ԏ�[|�4j>�Dh(�g�x*I�C"��L��*I5Q�l���F3E5���A����sL��q�)ي�X�u���T-��䚾��lP����M ����!
�P��|�7,����<�̻���x��S��晼�h�頋��h#S�.��>��1a�U�"��K�nS�T5���6��?�pǓ�����[|��$���s7�)c���v-���Ȟ���a/��ۄ��պu�� �k�RQa�7��C/���~K��Q�+D�c����}V��S���~��h�🗼|04�٦�$�uJF^�	��~���뎑��_�v5�<8�\-����S��LHa��ǑS�����P�0Z��$v����@��{�����1���������9�����ZEրY�r�HN���[n]d��̤�w���'�B\�Be����$f��.�5a-�5d1�f}���!9��g|a��d^)}:�1XI��Hc�5���^KCe��ds�j�!>(P���b7���z�3�4"	t��j������,CZ��C���N��L!�u���C�����������9��ػ�p�r����!�Ň0��"� ���O�1��
��s2Z.Ah�Pw�#51$�2<