��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>%��}w�K�P
����$"uI���10;�f��� u%J�Ċ����t(�k���_�ڭ҅�q[�Y���hB�1��
c�,�'�`� @4��B2݅�0�$�;fb�l�!�Y�l����&˄���ؑW��n%����zfT�)�u|nv��b����u�V���h;­�f�q�2���G΅�]�.��ۆʄf��9l��3���}���N,� ��f�B��o���@��&� OM����%"���w�0Y/4X*��?�U�8��l
a��iC:� ��R��.>1�x��4�.c���B��FZ�����1� ��e��|	qǫ./V�)�H�4x���>�<�f�N���5�l�@�@xK�q�BN6 �2R�c�.�p�� �i�,ϝ���Q㤲�(��k��������^�AN)��1$a(�C�n�% �O�}��|��+�R@a<��0�D�Tp9�mA�/�T�e�����u=�s�C��]�_:_��QL�?�W���̆e�ܺӐJw���0�v�#$���?'�}
D�]w<��|k$�¤���|f�a�j��?gi!h�!ز|PC_����X�SO�(τ���l��1�-�
�ek�����݌jfJ۰�榅�u�-H��DQ+W��qJ;���̰�4C�;�L��� ����-둙qi�L��ӗ�&��D��t�*�UX^:���OES_���/�I|6 ����D�i]�":����H�_I��N�	~�n6J���KG�4�`ZltodW�������&�2p�9�oc������#��}:��GW޽��VET'}�_U�:�R6��0�yqƝ9�L��a�lsGU%/ꊝ'a�N̕�޷�Usng�P�4�p�Z1��:!$�v63D���{��>�a��A�p�8����<��K��Q��E�79������\�h���,C���$�"��*jAAr�:���OP����SfE%М}�� ������%�Gx�L>i�>V2�����ŨU�E1,QJ�3��0��4Z�.=
���v,�'N/Wg��}eq{�hq-�Ж�8}�տZ���@T%��:��!	?��z֨c�`+� Qd�pw=�`&�c�P����x�����ԣ{'+A����`y�4����e!���(���KF|/���;M㋻}0���&�<��Q!��-�[��̘���f�o}֨�l�����\W<m�wU<�i���]��V�_0O�e����dd"�J�z�1��c=n��e~ܝc ��r�K��vY%�qt(��~8�yxw�V���Ϫ����|o��5�������b;�����ڰ)�z�Z�\\�"����s�8HDJ���[q��������j��K#�za׊խ��p���:�R��/��E�W�4�D�R�}b��`�p�W�b��dڸ=�cp��~�d�b,FK6�FZ_�mqLhA0��<�WJd?��[1���� �rԒJ,N#�n�YA����z�s��S42!�%�����+~H���9���1DOY�d\vե�w�GM7��}l���ޕI�G���1��lBU�)ܼqz<��j�L��}:��:n��7�K	���C�	�}d�L�0��2�7���݅֬�W�]Xc���5�^��f<��ɗ���x�2����^�����t�:�Y:�e].��O�(t5>����N�Q�m\����Y�>��Im���0��^�<\���'e@�&��k��y����R��UCN��ziȠW��5��	�P�>����1��U,2Yk�����5�-�)���Z�].�z8O���:�{x������ѤFvX�w2XE�������d�tf�g�4w`IǮ?�������	��L�>���G��q�>��\�U<�]�n4x�x�H�Tb�|T·��A)�0
�<�F{��$�Y�	��՚3��*�zV��s�8-�.��;Q�-�<<յA����ڿ���%�(��RH�S˨��IVj1bt���g�肄���۷�>}j��G�@��+q�S�8�F�e��t�vN\�N��Y�MP@����F���~����1 �>m��c�>N����I+��Դۻ��G	�g�Q��N���f���,���6��{˽*_#Bn�r�N�.ា�>b��~0U4 }y��qK��-Ҡ?{p��a+�'�+�C��F�m�T;�S�#�$g�Bu1K�Xcc�7���4"V�FNY�v�]W���ApD�NZ�	/�'v�w#�%�&��֫5�[D�ђ.�Q���޲�� ��q�rR��.`Th�¡��4H3	��l����\ Sߴ:�`�<;�����㰯&�z��H�ҹq��{9�����ާ��Y5�kezT��M�����R�o�pݼSHu).��]a����e+��C�(���zo�h�U�J��G��}��� 9�¯�+;�W��I��v8��7_�s:�a�ˁ"�.�Y���f0c�p�1�t�N/&�X���?�X��_�u�U��$2��\>��kwW@�Ko1;��m�#˸�� ��}�*}8�FT��j��m��h���c��.�����GK�-?H������-XHҡ�G���c�H����h����*��v���d�����"ym��n9�{bץ���(�T���_jl���k�O���PP�"�MqՒZ�]ig �g1keĝ��Sc�+ç�L��g ��7lUH��A	���_ѧѶ�V=�=Y��DO%��:75��n�k� Z!��y"�l�₮k� �`���?{�I�j�ҩ%ʐ�W([��+��.��{�JtA@T�7Q�cG��� ���LסM�7������9�C����L�W����F���g�%t=�̙"����m�,tp`:��Z�R+���c7���/�䇪����PH�"Q,`�]�/�E��"�ZW
�C`-�FU���C�W�Q��x��W�@�v뚨�c�i���������C%��jS�_�P�ɸ<ʭ�8�Y���i�PV����cSM�����_@1.�z��\}���Lg^�˱�g��_�g��KX 
#J��'����%@��6�~li�3Ycs$]}��)���lЏ���y�|��Ӄy����
��� `���"��h؉�A����,�Hpc�B,�C�C�U��5K�f ��-��,�=}�2���~ʗ`�v/'�ӵI��H��^3�	}����H@P�+�B�3��$�C�V{�<��$0�F���1åN��S����d.�B�I���iN$�d��8��~�LE�]=eE�/�j.��Ar���IGT[L忭�I�s�j�P/�2�G_[���O���l�(^�{EUš���֑���)�V���=��|�A,Q�&�&Y�?A��2[�Vp��3����&!�F��STa:�H0ܬ$7�,d�y��=ˑ������f�#�������J��*Xsc�Q��M�L[�'���à#�3�v��t#l�X���ANV*j�z��0QCO�n��Yw��<�y�R�8 �#3�ְ2��S�������RJ��J@1�)���}$�z��r�O]�,��;��1�
�>�� %Ͳ�+�y�����"�.�]q��I�5n�b�
Ϻ�1o�� _��)�)M�`��y{�w�i��;Peԉs|N��� �Q�x�?'�q��M�Э�|`!{E�{��� -`�ߩ� Cf7J��:G�`��^�XRn����6���rJ�ċ����qb�~�e���7�2���vl��h.Y�ʭA��X΢}�
Q����P�3��̰*�5 �,-+vh;�N�C���=ǣ�쮌}�h�4�GMZ߿#>C��</�o�;��0�����	<sۓ+G��Ou��
�m��T�E_Џ�On.=A�u��YqW9-G�A�G=o���U�S�����8� � +�����"9���u�ٸ
T��
�X�Ż��W��w����Tj��c
�j|F\�vȡ|���N�������ZM9T�v����j)G]0�������`����a�06N:bگ��ɸ�+�l[!�\��r���tM�D�y��7�tN�BeԈnϱ�Sh��s�]��y������ޖ���H��?wZC^����UV��)�	(�1O3�!�Q¤�v� �}���vT�Im<��vؓ��
�����=�H�1��l�z��-�fW/��<)^�Ջ�x��|�5W���zp��ָ Ԧ��6\D�(�������xI�O�$N>|{�Hm)^� �)��U��ߵ����2��}s�N��)�څ�s������=�[��$:�����]�X��F���I��m��ͥ���rQI��9��3([�B-,�e�;ތ�n�G	���Yd�q��������&�38���5�86�Bgٰ[@��b o����P���r�G(�;xr�ո�?NV����oF?i���fVG1 �D��=�D\�6m�0-]�6�1��e����WV��w����}�0>v6�$^�7�[B��9�6�b'v!���T������!��sBҸ��D8���/x���,���j��cE�;��A/tIM��2�8�d �f�D�m[��in̗��"\1�]r@u_�������	�j�uuS��ra��s�uw��z={+fba��2 ���?*�T_+�i2��x��P��%0$�K^�x��>��PA�0y��1]b�؈�n���/�N3�]B頵�kĿI����l������|f�U�>do��S�lx�051�RM�����<�	I��Td~��4�����ǵ�9�����ZL&lb���.ɶ��K�0�;����bn�f�=e�M��X�}��3��5�?G�\�V����������F��ߑ��>}�7S>	ř��hYX���ņ��򋷉ez�I&P�=��a?�Uu�(��Ӕ�¥Gу����0�B�zp����e�����\#q�tw=z��`t�a<��.N/ZĴ��~p|��?Ĥ�?��ΗM#�7 ��Q��Sk89�a惙��.u1lD�y/N�3:�S.�UB9.rE��N�ԧ�y��q�]�0U.^�ޱ������(p�G�t����-�o��ʷ!g+��n%
��ɬ�����
Q�����я��N�Q����Q<oj�Ƴ>
�d��'��_��'	�'q@�nr�.�2Lob~P�e�^�FcO�� �,P�_�Ice���}�W(�]M�A ~;�K��@��j��"��SWZ���Pa��?T6�ޗ��/m�G���e��ԅ���E�����ķ?��㰌H�$�[E���-௜�F�A����am��愈R�1��R�m\&C�n��#	��&_��:��c��P�ey���~�>�G^EJq��܋�y�1�\M�+�Q�m×>��P2�Q�gy?���Oϙ���������t���Q�[�m�ī�jP��1�����%���.��o�?�x�U1mQ}-��/�|���������a{�.�6��Q��rko�c�	,�L�X5vӫ�\�w��A%���j�e3%ĵX�P�:���)`����l��I��"�XRSO����8�<�=��c���{���͏\�C�"���Ox�６O|�kN|��k9���g�š��s�v���i�{vZ���ɱ�b��w;�Hx��5��no�n�m� �b!��)b,�˻�6�ϯ��n����C<����%u��4�@M��<Y� �գ�,��2��b�z��V� ��������J��A���Er2���	��x9Z�X}~��_�oM��')�0����\?iN�L�9m�`�G�|�`����`����������ً���;l��4�<>T���)�O�N<(U��wGU��hF1�{a-%ᗾ�F�j
z�?��2�;~�g�ȗ�C�a��&�p'VF.Ғ�m�&P��g)AmJ�T�8��-Z��*�j�q����$�b�����V��;}ׅ]�L~��"������[�v�`���F�ёM�!�t��������&�3+�"L��gT��ۚc"��(p�����.�+�<]S�~����������js���/����G;�ϓ��F�,����<�����y�(��O�|��,�[�J[V)��9}}7C	�x�:�������P����h�\cg�ED�Ln�r^Q"G�eg���TblU��Cڞ
f*,�r��[�Z&�PyWq�h�A����|i�~3�\�?$�B)���2I�����˰��Y�����Ek�ڃb���5\t��R��R
��
H��cɈ�A�)g�t"xiܩ�^��NAp=t����(�q���uI���Ok�D����B&4�܊�N� O�Lwrdo����e�!�BC�J�Q��d^rKN���2EqJ�΃��@�����
�4�A��?�
K��@\0ѻ`��1Fe"�J�B� r2`5Նw�T^�q�x�v^�'��,��"K|®�#K����'� ָV���x�x�� -�8�
ݫ�|BG��
�;�id���</+�C��s�� db3I=�2Nm@th��]�E���
�xyw^�5��!���}���ߗ�A�A�914h�y'�"ҧz�+�(;�W,�޴su|���<�����θD����/Tʎ�Vv�rC�HY%��B���~������a
$�� de��X0ᵣ�eS�4�]����X�i�T+#����Lע"�b�*�Zb��ɸ�{F��(گD�exϊm�@)��X"p��O����R���q��M���.�jE�M$��<k/��j6�=\���Q�|����Mλ��.P��Ȇ{H�;�Y�j���(�>	魈"�a
1b��:.�@�[�s � ��TL���cn��ٳ�����t}
q�1�Lx:~ ���\�+|���ۛ�1O�ӝ�K���ʺ(�s��NS�>)P�CN2�,�"�o�]sAf�!�X�+��[�&T��"�m��'���Q6̓[�q?*.K?w��h��b|���Y��@��O�4���,u�O�q�m�)ɻ݀FQkM1~��Y��ݍ����RƤI䥽Ѝ|��ϕ�.U��b8�6��6)<���Q)�Z����1�=�E�M�p� ��7 
��2y�{Q@40yG4�dE�F���~�"`�g�Zq"E�hE{i�}�do������8�	v�Q܌s���盝OI7B�t���93���k�C��BO�o�j��v����>tu�ӡj'�\�DS ����w(^��軐o�쪹aѧVH_��/�]T�����Z+� }�7qW�`y��-/-(�Q'2(����#�th� ����y;�/B����a�K�1��b�+U
�%b�[��c�\ �?Cp�5ճET7I���_��CLק�2��Xc����0�|+�^3J;�4�m�_�7��g�����%���� ���wf�4\�9F�PI�u~��ǽ�ɓ'�6]90VL%33Һm!�.�2SRg�E�	����G��ʒ`e��v˫��&$^'�$d,j,�gxS/��;�7'��Qeg~sb&	�^1!�5�0��C�"��N������E��O�'������cJ{V<�hp�y�bD��n��5�/B*��}zD�r�Q�L6�a�Ɠ�:C�-s�32�ûL�M*��T������QN[��eo�&�e�H���?�Kg�H}����4xoe��������`��+����8ڽ��_Q݊|^����?��}���=�5�~��{��$�6]ۥɪ�o�X'dU�K����
��Ē�I�Ĉ0p�n"O+�a�	D��U;����N��(�n�_�}m�x�(�2�1~hz��Zy��x���Sɥ_�p�'�>����a"����~!��,��~�v`��v�V��;NjGG�k1*���+.m��U�C�Eb�< �)J��Q���_m��sK�q�HR�Ku�k��V���Y�	G�=ʟguh3�y����S�PZ^�Il����yf���Q��y�iBcέ	�ٸ6�~	��z2��B<�}�Tܱf��O�`+z���x��8�Թ]�k4N��i��%+�x�)��Ȟ���euo���"Y�҉����Ұ�J�l��E���"[~�(rZ��r�'�F�`e�^�M[�~�����Յ-�}p�YWX���)4�f�в:�_"Ƒ`�P�^��%�\��ɇ'I���0Yf�<���z"AvӐ��wԒ�B��2R������*�����F=��P��S ��
���C�\O�u�#NĿ�?���پ,�L�>Q���k4�^�{0�W���4qt+M��%��FW��|��}�Z�O�WM����vr���M�̸ȋ�  ��ޣi$�(�S�~Ⱥ_�����<�pf-�F4�}�'���˘�tra�0�s��V~�#y�gЏh�>`��d+vŃ+3p渣%
��hE�=.*_��*�
W�T�1�"�UB'�@Ҏ�����ܙ7!����=赙�{�"X���d��o�G����Ud31�^4����M��f`Έ��`�ڷ�9=g1���
U�7��!/w�ɜ�@]g���Ղ��v�|}��Ao�);]�Ѭ�,%�,.~�D,p�x���:\l��hn�x��RǍ�\?1M�F\����Mx�Z�K�
�_��<�U����+�E[��֥��2�^�}1yN�:���!�S�HNĉ|�%���{�gtޓ�t`u0�H�"CC=���>�3a�{�4h��׊%�<��90�� -Y]$���ct&8t,l����8��	��S��Ν5��;ɁP�C�e���� P|�$�\��'}^U r�X�^�������'�n/p��'�_��EӢv�+�`�Yl��~������J�4�-��a�b����e���}{�]_.���_MBN�]T��\ֈȒZ��?�h|Kq2]��@h勻;�[�ZxK^���Cm��%Ǭ�+=�C���H����;T�@���or&l�R9է���,yH]-;����	���8�"0r�|`�16��yP)%�sI���W�Y3E�$QG(��/�~���,_��qC�?�Bd��`�8r�#�'��K4W�$$���H�O�ɜӣSE�((��1���E��E��I�0���<�]�=ɟ��oK�0��*�bm�G��\���	�}��L*:�C�V��b���b��,0�$@ֺ�5� XB�=��)J�f�lb-o���"�FN־�J<�1N��s6�[�7���M�Z��֍�r��AQ?����؋'Ϥ�w��:Ѓ���2�B$z��ziT��!�r�vv`/w8@�����:/�T�{�,��a�I�ec�ԜD 3�Z�=�3�~��C���t�xwv��h��uY�#'�mC59��b}r�'HV���q8M5��D��iYl�c�1���dH�0��M}nVB�K?�7M9j��Bl���닪~��E9�0}��S�O*#M	�p
ܫ�CSۻ�U���VH��������
�P٩�)��Y�K)�?H����1ű�C��m 6J���)v� �z��U&��L� �^�>�t&v��4���%�%�'�C�?��2�.cq�+�2Q0���6;e�&"�5�p(��ub��%}v'��N���ݙ��d�0{�n
�v���=W��aȞ%���eW�R��z�9s´s0�R^6��R(h�<��qe$!�o���~dz�#�f�2��ba�����ȥ|H4css�%)>)I���.e-鈑�����P���n��X^R�495ќ�,�zP���,O'��)�"}�ܣ\���"��&�*���;O�'lё^  .޿��w��a���+ѯ=Z�o�����Zk�:���O���@u���#����Q��>U9� ��b���;��H�>�oE�[�Np ��i��.�`m����B�#T�]��QZa`���F�/ ���r $Z�Ӕt�Po��ZS��҉�f2�ZV\��PDP�x$x%�V�� ����YUgm���̰�]$u�]�n�z�į90�bdh�i����g�B�d	�C]�/"!R�npG���L~� ��[	A�>G�B� �z�^�"[kf죾g�AQ�U�1h�_��4(S��۶x�������1l��J�Y�s���ER9,�!,b�����n9�s�k�.��.	�G�Zq�b��H����x\�S�u}�7J�6�_5���6�+����A�e�i�-ٙyQ;2-�X+B�KYdC���ƛB�Ӧ����5�@@�B��s������S�#��B��vw͈$�M��tNv���v]ڍ���A�`;��2���|-)mi����Zi(d�|���A�R�"�pp�'��S1��G�,���o� �O<���M=/�I���u?u�"1�y��/�]T6�o��Ľ`u��@����Ҕy(J-�Xΐ�[�\��̇~s()�* 5,�Bd�huBj3��z|�e@�73^���G�O�t�Cb�I:��#QDK{��$匒�������Mܣ���1�J
�%� �'���f0˗�:y N�4�/噢k��<�F�1�j����W7��P��H���KR��aU��%X�wx�V�A���]#�~J:m�J����+u`e>B�~E�����.<�hΌ%����T�/�y<���ؙ$��tGs�1�&g<qV���!��7�!�.t�D�{ktWo�/�5*0�^b��\�	|�|K*Mԟ.l�����s)N�a/Q�}����=�M�В����6{�s��;���p���[�mQu15D|8Z�B8k.���1��*_ܝ�B�e���/#��ߵX���u�������Wf����w"ާ% ilG�K�ï�`{2F��QT1\�l"��������g{h0���wͲ^t�0�Κ�;��m¦��j�H ���otO��F��t����,� �ÊE������y�.�;���^!m�����g�g�l-O����땍�dV�N~�����E�S`�u�g�Rә<��5i���w��~�9s�Ɠ����kE��䛰
���w�Y�N��x��̃�^։B jg�Z;�zݦ�4�� �,��eR�cﵠ'U���e��v��@y��+�3"-N=M���ky/�=�{(r�q|#�S���|&�M����PY�lځ����?�cM�˪F� ]ȌLb�"�x<y8P���%Az0_��0���zEǕ�Σ�6�1����E�	{��܅�,/\�yGZa6�Y�̿���.ٝۜ��'��w7c�����{��<���d7`����y�t��rgqb�zG�âЩ�3ږ��=;�*�+�<~<���%����4YK}�#��	W��A��\�_`��A�Ob�td�+��%)N��8[������f�a��0�sV���J}�����k�0�C�M��s Ս!u���Nx	�N��M�l�dǉ�܃�s������/�b�G�� ?�����ߌ�O�Q��\�m�i���8���sϿ��