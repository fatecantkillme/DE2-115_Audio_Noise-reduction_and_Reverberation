��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8SjfSު�U�.Փ�"o���Ol>�g�t��"��+_k-vz����;@�[k"W�3B�|���m�xbZ ����="�8 ކ��Wὣ�3��'��.7 /�ȆIc�Z���ja`�p�׭jO��F�����L�m�m(L��=��+��ڇ;��P`.#��١K�'|��C�J(��?�R67�d&�a'�۽��P�t[ü�̝��WS]���nm>�wˆ@R�U �I��6䳷��$�`��t|��lC�q��0Mc���Gq�w	/ƍ�ţ��kt�Xх����������G�V�mΐn/i�M�R����9N���E�\*�Z�#��5͖[��|+B��޶E�8X�VmL}��v�\�uM�]!�Uiq��ʌ����B�eX���(x�Ж�Z�T�3�uVaKGZ��.4�����q�hc_M<lO�e�cvw�T�\�E��igM�m�x,.	6�L�Bѳh�,y�LS��N�����[Bz%�������ߙ�gk8�?�K��O/J2V�FGtL������N*��歚d�����u��2�XHV�򄝰@~��2b�C���vNx�^*e�!Ԩ�yUp���nX�8R׹\µ�X���m�X��N��U���	u���(�F�Í� j(.�F�����gYm.��� ;�Z�&���s����7�C�	Xa1����5�:5��.��Jo��6�t��-F�s���D-�n�^�n�4[-8��j���Q�F��EƜ�V!���7�Z�A����˰��w�����[��*&W �pA�:iv媫 ��F����L���>�'�������Z4���WC�#�sͮ�3�|a	��Z`xF��q*S b�<�f��+o#�؄ZU�q>LTNYо�Ӓ����Bj/��3����h��/ʳ�׵j���3Z��:D�����B	������>$�����tE��i�msL�%�����\l��f�@{a��D��p�I�3��`���� ��رi�ɚ����1,`�~Kģ�����z�~3y��g�2�]f�ކ��3ӳ$�2�"2���٠m$�N7٣Є��x��j�}c�@]m*���L��>��ϒ@!���=�[8�p	?F��4��@#B��ܪA�@H�8�6�gJ�3�X���u�Wj^�����ƸR0q��0�]l�>:�L~�;�<��ˆ�3�fl�h�V$����WF�p��� L9@�[�Hya�%����#��(_�t瓧>I�K=fž`��'��yx]6��
�6"�$�K���{+��+�§PT��K}"���Z�gf�N�i9����숯d�ؚnZ�j�s�s(�}�#ދ	QQ��8뷔g&\�/ ��nJ�D�h�J�{B��9z�
�%erwũ�@NL��C���I���M~��z�����>�R��XN��7������,��mBF�������'f������@-��3z3��~F�p�����|��U���k���=4)�D0��kI��S�v�B�:�
elj�P��6�[�����R>�USS���J���)�Ӯ�`xH��;�3�M�n�ί�|wj�^f�֔Yv��L�{���7_�*S�pR������&�U[�1��PR����?�@cT򡄻l9ŧ�@��ԗ&�V^������j�=�w�m��[�xu�7�jO��#¾DTw�%=h��fGJ a�`>3�*��"��&����TV��E����v2j�;�:���%!� ���Li`|qiA�xW��
���h`�}��՜g�2�^�����*���:X���Mn��r2���0Qx$�%� �Y��uy�DA�����5�;E�v0.�F��פp��Sٱ/��ߡU�6��1��q^0O}��Sb:���U۳9# Udgo�Y��dL�2Q���uT���a5�Lbp[̈�|��9|H�N|IO�{9?@�$�9.���M�}�vBI�0t@l�tAK�}7�`}JS2�h�"k���Q�7ʑF�c�d�
���;P���׸��1�t��,��W���i��C�`�S��������GW���c�dhw���>���-��|n��&�4�8�]��ㆌ*}��|���������Cs��U���__ԟ�	�G룕�W���#Fa�A#II4�\�<F�U)Z��"��^�>�]"��a��u�C�!Ҵ:��T�ב1�MN������Σ�d��#��{:'���u�Xѩx��B%o��I�R]��.x��2�D�*�OW��&<؈ߍ����, �$<�wr����Ef���ǜ�;�������Ն_"IEq���}����ix�o-�`q'@ʂ�����	|����="��c�C�΀D�a���$J�1�c�!|�&f�,Q�+��a�,b+�u�4�v�m ��~�8E��~��7�1�;�˘DwSV��,�72]d����s�{�a���J5�P(♄��L!I �E�c�a謏] �D�TӜ�o�VX��P���B�۹�]�ڍ�Ց�/u�w�O�$��\JR u���H�'�W�U��^�I�`��k���³I��'��"B].>�+@�o�^Y�?�D�+���%H�Lݪ\K�&A��{�/ir}���q~��-��	4�?aO�t�3q��3���H�Ȅ{5<FM<�s	b^	
q��ƚ����[�w�G�,{����?ۛ���	�M�#4������,��r]��������!U��Ȧ4D6|:�f�_%)���L����~G7Fi �`��
 ۶�C"b�-��a������Z?;
\��x�n��e,E�j�{ajf�Έ��+ ��f���^��(�쳀N^��N���+y��]/^<yt�~/f��Z8��i$�?MUL#�Y<�gd&��9rK� $R/5��e���z"�7�S\H[��(�&�Vog][ /{���h*��ۺ"	_��G��oà.�i��|�����]��EZ�X����B�
6�y��Х쐡�w_�Z\%���aI�
ru�i�j���xl�����g`���O߁��Hk�hzU��Ƿ�i4���ϿZ4)�-*+��)p��=HGB0�z'r_A�`n����:'/F��c·9 |U�f#�*f(�؂7�= _P�<��\�+����I�_zWV[
�������ׂzJ����w]ZP�1�����Ρf6wJvY�VR�W�>�"��k��B�+X�+E�h��}\�9�?�O>}���[A�	�<���a��`1��	V{���z�L�j���|�>�G12y��q�_��Z��uF����U�M9��hZ�U�5,52����^�g���]��wƝ	�OKA� J�ۻa�m�ҫ���f�'._��s� �KX�n����5E��O�z�!��d�AuEW���C� ��+
������|{�iu�P�ِ����~�|*څ<W?S��j�D�y��z9�C�S��������R�9p�D���{~��q�	���6GW��H��5�W��(�8Pe�e[�R�<J�iO�6��I�_hc��T����M�RL̀�����$�.��NT�8�h�s$�	�ç�R�f�Nj�soC7щ̨[�o�	O܏&�Y��̒�l3y���Y���[�>� }m�MV>5K��@�ҲXeS	/�K�3z��zt>G<�D��7�eV�!	�*�U���Ѱ#l㚳[�q�:�x�C`�@_m�3�>L�e]$0׿�0%�ܕk��X/l��\��\�w5�6]B�g垭����E�-�bG�@M�=YѸ(�l���J@TV'������3���l;��g��nyCU��rq��\v䊈;^��6��3(=N�M�T����8i��s�3��8��t���������]�W�&�� �!�G��ȱ^_�!r�0k��2�ͨ�8��`f��M�c�+[å³Θ�(*���H�-��Yk��9�F����&c@o�?��7�~q>TGO�������:����k�N޸%���YX�wJ�N�@�W[� ���4�p�4͗���ߕ��CE4($R_͙ͷf����v�4��K65B;~������)�\�mW�چUR~�ha��65YC�a*O%��8�Y�-��CL����
.Zm�N�W�'�!�ݴu~bL��Ca~��A&VS_�� �4�-��źN�j�ht���J��	�)�~�ۿsVջ�� �$bm}�-�����1�
�Kާ����4����S�G7}F�Y�����&���D�*ĴPF�����9��@�&HO��6/h��Y�h�o;�.V!�:D�/��5�(�J��w%{�&I2N�p��ێAQ��s�=T�� �[y�,�#P�ˋP��%�V��(����J"�=x쌄���\�؛��?VD�d����6����Q�}O#�P�;PƉ4��M�]������v����xab�w�l��p&�5=6�TZfB� iUi1���Y��n���C�������'c"> �x�u�b���	�X	�P��Nq�1����az��&�>�L4��%u�DHTAa��u�'<p*�|,����R������6K�l�h��Lh���ߺ#Ԟ�l�Ͽ)^A�}���~�̕�|n���(O���#�mx�y�B\Ҋb����Gv��n�N\��z!Wb�dV�\��7� �(ֻ���g�k�kgZ��%Ž�7FN������������EP��`@�p�A̠r>g�Q����S #�� $p*Q���A
�D6�����?heN!�`�s�a���xm�Tԧ�����1n�%�ED(KȔ��b|`�
>D�4�݊����pW:էٓۑ(Y`R�h����&�nքl|��ޘ�4���0(I�5Jní*�/z�q�N ^�^�k��s�=��(���|��bKl:�2�!#��i"�wY��� ���ޭ����A�8B��+�)��w�tS��	͚��W:��]Gȇ^�G�l�XǠW�䋣 ���iՕ3��x�!U{~L˟����U��ش�O�b	�»|.k��	߫�{���qv��M/L�j�.a�!�mON�E��9�	A[��X�T�|2�m]��b�H�7F@��3�޽u,U%�{kץ1O�J�t�]t[��E��[�5r��Or���=���1�&�����-��W�e���G�`C��,��{�v�ş�Bcn��y5�6����UO-r8���$�>�t��E�b1�D\u}��@�]�U[��;�m���MOY����<y�d�x3��4~������F�Nq;���	~�����|�2Xb,���O���#�_;��9n([R�7�hg]�'?⇹(/Kf��FK�I&c�*�{�b3�u�V�ro����,FUF�l)w�ӭ�]�u)ϼ�����5�Դ�,C�h��X=E�i��T�m��s��8A�mx�Mܝ�aV�J�kn��G�ߕ�򄒯�fTO}p�ʟ3���!Ҁ��x��b�n0�Wm&���&R�'{��0'�v��UVZ ����A�8S`:E��)���/���ؼ��M�w#i��#�v�T/���7^9�sD���rJ�%�'�T��С�SC��v��8�͖�u�額����dڡ��}g)F��(��6e�(⩙G��OT��/��h)�3U�K�!L)T:2��t��9qXsD�'w^�P�:�8��ṑTC����k��6zD0��nF��;e^<dl�3$�B8�3�zff��K�/���0��!���S��R��i'�Sͧ29�����0�|�L�G��Z�C��Na:�]�:Lai�v!�&7��B1�IXk;F�UNlp�[©�ދă5?oM&	��5E+���Ѿ*b1�j-�sdI#��s���:O��}��y�,A�\H�q�]�C�����>� xX��=�-ᆪ#
�&=�Rvn\��+�/$Jt���2�ѐN�c5�.��z|�=0�,�5�@�l��$���V�x�X�M��є��L
U�H�99�E�-�ض2,���B�f�}|��@S�7�gҨ鐁�݌�\�oA���]���.q{�)r����Q�.8k�X9�罨]t�Ql��Mc��E.δY��EV�(��3'��o�,:�pU~���R~�Q��$V�1["x7֊qo[��^ڇKFzWK)kN���q_�~��k�L�&��aH'����{<���ʐ�oy'�+,lB!�^j�+�� `
��k;�X�����G� �{h����~��ԧ�C[]t��~m�9��Z\˃�X��� ��F����.����n�(���N����^���u�)������v��蓥�;@��Љ{��2�i����8��z*aX�$��J�������9�%S[��:b���{����]�0TYR���s�V\ܩ}HȠ��]h�n�P�ϱQ�.�d����J;X�c ��m�V'���o8P�V��I�+0��u-;�0S���]���l���J/P�|sA�'���5�W�ͬ��v2ǂ�������ʸ�u�D��<93:�$}Ƽ%>�@�$��j�SV��]
�����c�&�:s�r��8�7��\������ߜ�	�W�y��<��"&~ҽ��p,����6�8��m#�3w�d�b,JN2a�D��H�2�!6;�p��eh;��RJ�t�R�xo*�:���:����59��gv��h�p��������G0պ���Rsx����?���|��`���h�~DI�v���B�%�wSq1C�����2���g��Zݨ��IP�����������2��zƗ����%8Ӫm}Q|����@��B�&6�>+̖^��d�2��dy�:�r`�J-Ɨk w ��$j�����Knb��R�Ql|_��,c��	�n�kL�'�r�	���K>ӣK���Ξ��N�;|�ͷI�I�Y%��ʝE�k��o�''�9�PX��u��k�w�~9�06F!+��C�L�)��j2��>�I�����t�2&,ɏ:ѓc�-�����[�܋��Ɲ�v��F�tKK��-铘
��`�ho�ӷ���G�eU'�0�ǋ����r*���o���Q*D��?t���0��G)=�7.!����M��e5�Ԝ�)6���d��$*Ve{�c������Z�[GW���AՐ����4�]�*�y�wKP�DS����<��ʆw-<_Fخ�/	��a�.Y�su�RP����,!j:�Uu��Vc峻��tF���-9�fR��;��\�6n���_+���P�ǟ���uٰ#�$�b���1xb~�пp�$u��r�R�EkU�9��aXQ�5��G0>IϿN��_
���~���TI�k���\
Xz1`��0=���G���6��2��jo3����T�	�;}��D�].�f�.X�&W��:X�P�5��x2Ks ���MN��x:9M�`�κ6������,�d�+��]����X���}rZ&���H���/��y�����Ծ�w�jO�B�}�y	�&O�-T��;���]���<A��ڞ��^�����V�߮��~/}�c �i�z|nƼ�J^�r���N8F��WE�B�}8�"�*� �X��[S?G���s�#2B����
�U����E*q��lM��<8�i��j�7�������G@�N�au^�8���U��جg`�����̛t��8x��wQ�li5�ك�靯���]L��Q� KyzM�r��s���	k���C��6�@pa_27��+�Y[�w�M�$T4Kb����M�tm2��f���!�(�.�7x��^x�<K�yE�^�E~���ZM��&�������?���(�\���yg�OYn�]��y�-;�%I�,8�.�J��	6q#�^���9Y'�����|��������J{� 9�3Z9�+��b+��P���V)��08�o�E�O1K&z��N�QQd%�����F �,U�h���x� :���X�]�s����t��UB�3$�h�-%����5$h���ވ~�G�#8.���18�c}T��&q�Ow���Nuح3U�Jm7��c)��X?dt�~�����W.�����;�I�� -~iG3g�93���N�=�B�l˃����ȷ�Wp��ui$<}�� �3��[th<��8�^�L�`@Cq`�±���Mt�7Ϩn ҫ�
�hJ�<ؚX5B.���^�`RȽ�+�T)�p�^��1�����tF��J;=跂�1
�ԋ�	O��gW��8��4�����~++�Or&�?�ql�O}��ߑ��X�r��f=��p6|iMF�}`jٗ[g�PuA���\V��iۙF�Ħ�K��D"	�F�uwcUōQ	�(�bp�r�+X��ƥ�כ�����T��"��Zx.��[�"�"�}�J��\J\��D�F�;�NfH���@��VHy�;�z=�]���S���}�l.W7]��c��u�`yS�?�]�>J�#/�a�~a���̽�chr����I&�2],@�y��?��B7�����G�ϯ���b58>��=YdP��f�քk/Kz��e�3�=���?0�IϋFֆț����<�C��Q���c��9@^!n��r2 a;�JK�� �mb�]�W�}���? ��|�a(>�]��| �uj���N2��Ct8�!��8#�`����|N9��"�Wړ`��Ċ.���_c��6B0Z-={�8m���J��
S�r�����~~���+���G��}��W�@��Hz�ay�#@�	��� D"m�D�~HXnJi6DK��^��1��0L�8'�h4�U�)q�|kT��OI��7vMs�	�jk_���$�#�JX\&���,�H�*U��^��˼���e��m.S?n�.�<{��X�4��P�}�z_Le��-;�L,k�R��t.��������'����oO��Y}�7����-;-�f���g�H+l�q ��Z���N���n"��dB>IՓ$`l4s��-]���q��z�Y��t��1O��Go#�n`�;�k�0ܩ$a���:�7��d�JF���4)� W�Il��Yz)�q5>n�q�z�6�Tڵ�y����6U"�>�q�I<CH�ؘLQ򋶶�~%�G/4���}�m��|�Ǜ��I��kv���O�cw$F��ls�u����O'����{qخG���H��ijC��t������f�L֢���)���ԕ�<���e��8v�o��j�=�f�i�i�7�����d����s�z>|2�jTXGzw<�B���1�EK*�ȟ�o�K��őf�o�!ʳ#ހ$��p0�yu6M�C�,�����5洽C)z���۽�:G|̂
���̬�k��|�5��J�
��/W�fM1�J���^Ӿ9U�^l��|�2UG'p�a�`��&��ܞ��=s����,����2\����#J�iְ��_ڜ�%��j2�1���rkD7WJ�	���v�O�:�!� ����?�rFg�7n4ڹw��A��WR�l���� L8���+�ȑЁ�9�Y#;��DO�]����^���`���e��~.=m]� ����@�Ȩbi�\z|c?V�
aMlyi�-v��0��qI��Ƹ}t۵̝h=�'�IJݥ����4��K�u�-�P%�i]e�#��yU �W��|�:�s����r��-%A��>-�7� ��p�.}Z ,2ʢ�nUh��,ߐ��:��R��_G��5[O7lYW�[�-��fE�m��-|�%%|���^I����}�5�)2����i������??83հ<'��1b(�؂��Dg�lw����1�l�V,9�։`c�CC���g*�?P33�$W�����eC)2d@��ee���lD��E?�� ��/����7�9����{�}����~8��?�@'��];1���"�u����2�{���cP�K�zF(H)2��Zn������RҼ��s��[�
�QL��
�zJ���-��P4�Ɓ�����Z�����%�p�TɰQP���_����0�4�Gk���"3��I�����T0`8���^�_Z6I��ų��C�����#�|U*b�`մ�@�������'���/� }Ar@tך�RE��r�Ys%1P�0o(������~�z��G��/��>�%:K�
#�QH���#��3�X;��o��x���5"ah��X� !�� +jV�Zv5��z�i��hQ���^vS)�ʷJ��Tި����'j�}!���r"VA�6P~�-Eyrj$���dOR���d��R�r�ܢ<����ӡ�r���8uF��f�J�Qs��v�b(���"�j5',�YI�1b�eq��mr#Ѷ!-rr��͂/���uʲ�����?w��b�G�-�ߺh_k$W��9�u7��qC��d���L��;�u����\�*�mH�鎪�?%�Z���,ɯP�Zc�Ň�fg���׻E�����tS�,�(K�X�	�VԬ7��S��^��+
�Y�r�?�4y��f�=�*��)��6!A3��J�����!L�VvE-���R�Ҷ��95l��U��Pj8r0��st�3+�V��'��eǪO��R+y[�X��`�ksۋ�P�~��,r[�q�^��a��Qz��Y| xH��$�^��6����{��V��!E�e��k�I7�,��!
P5�e瞘������%�d��wr�@��F�'	��tQ�̖��e��W�� �邒��5����zb��Fi��:���h�ʁ.Xm�����KV?@���5)�B���=����ᬅN��F:_��M��P�gX�_���޻><��q4{�wr�N]���O���\��]F�Fɜ3���K�DDiJgS���<�B���&�b��<��0�DޯBω�)|��F�f��f���>�V���>�0�(�U��bR�=3m��gp9$g~������K0��A�J�᤾�tgD��q��r�&D�Rg�Z�T�x���@^+Yh�0�"%�/M*mө`�7��^S��q���m��^q�ٱo�KR�퀗�rzX�)�ʹ��)o��ҼD��^����[)�^𝖂ك��DH�I�����u	,w�+;P�>\�H�U� R�,��k�}��GI͐����z��3� ~�Fs�P!�4����%kH�r�\�h^(�� :�?/,Kݡg���V$��;��:�HG��\�G(�JB�א�u<�ZL#i��#�����5|�^i����GN��{����0���\e�N�Ci�b���c�xh	'�����/l��%R���8�xR)�L��b]�Ϳ5?,EA��#��w��O��c��u9,.oQ՗�4;��e���nP��n�P�&�3]��>m�e$�:G��h��8$���� w��v{�� @mNI$�ЩbG�O�+)�4�[@����nE�,}�����t �̯�a�y#w		��2�ş�m&� 'Ev2E�:�י���&�e�'0�?���ي��B�c�@M�'��]/���zN\Y!�d��=(Ծ(u�M��@nG=����q�Ѹ@!*��'�7�h��Aǫ�ݾkB�6�#s�OX����ۀ���%��T��[\���p�2������pݚ�۴�!����2 }b������K�&�@�����x�3`���1���i���`���yM�1攣�4r��N]���+�(k>o9ȧ)�#���g��s���,-�ڷ2M��P��.�Tr.��T����]7����y����nZ�Y.���5CE!����k�n��.�-TX)��������WJ�]�zs�����q��p��at����[��V�k��{S��N��9�nL�cwS���6�����9t�Ґ�h���^��yd`O9D�F��g�o�k��(G|�E G��_���7��W��X�\�Gf=���=S�b	a0R��������ڋ�F�R;`��+�������p-Z-�-NLY.�� �lWw�����|bb���� j�t�hY�0�+Ч	c�D6��vn�����ɊB&cE��~�+_�d׎�^i�y�V�<kQ �+,q�	l�L����#���w��A
MH���j��n�����%
�-F���~H��7M��5���,��-�s[;��ɘ��~O
�<��\�Û��w���ץɴW��;�w�`U��v���CV�!֯���SS�p�aO�0۵ViIH��9�����zE�~��@- `4j�MM (QG0?k(����.��=������.~!Z�Py矵ED3�E�qM���q>����T��Q�EN���3i��38���pE�K8B隶|�4\'΍u\�S��ߧ�;����D������d��h���l�d�x=߄��z�=_�؟K@�a"���Q�G�d� L=]�ws�Y�h�� �+����l��D��m:A=�E/�����E�GE����ߘP�T[国�v��Ce��8�L� R��D�������>��V��ׁ�?x�����OeF�g5�hk�q�W��� �/D�g�
u�AdmUu5���\�{4:tj���X�����j0&]	@48�oi�X�8�M��/�q�]��˶X�:��������}aAyړ�.cD�/�J:ˇ��c%�3�g\��ȓ&��0�_I��O8q^��k,Brr;�TAޕ��80��HdBQ!!��LZ>*�XU���(��Ō�U��
�{F�l\*��ї����Y� �
-X�>��� ��}ʁA�Fe{�o�m�.����Lי�;a����(0��Һ��2��v�_y��]��P���Af�~���>.a+�Hj65�A�N��,ع3G��߈�9{��%��V�l��̩��+�9�V��ά�dV�`��n��F���)<�����"�w��'j�=4���H�ʀ��%��>d���;&�K�X
T���@:v��$��`���j(�
>��5�իn[R�%F.7�5K�g�fp)0m⩰ror���>�mۈ)��h�԰�~O��Oiq�*���� ��H�W��D?0-��dKP�Ӡg$��Y%nD�z��*����ܒ�j��xb�n�H0/��؏Z�-� ��;�~�Kn7�s��7Z!�nQ������c��z�5 x�q�_��z��wJ�U5��7lv�+��2p?ƣ��)^�_�a���ਅ�}*��|x4+M3�rh�MO�|�7��=%�l;?���0<=�z9�t+!��gs
��A�a@t�o�~f��c�	��a��!U��j,��k]b���67?b��ó�)��lA�+��[�0��\��r>���+J�|���� �H�.�r5�D�M��險"U�o=x��
�fl`6�}�њA���J�����
,�H&��0��$;2���.d-��Jj��̴������X2�Dhm��)tIc4���Y��%�x�dl�İS����>^(E�8wCu�.�%˫��v�5�����g>9�qܿTU��_�˜..<�RѶz}��l W2˄3[/���?F����WQ��Ѳo �2݂SG��g��*�P�bģa%���chD�K�������9R�g��-7}�����������|�I����?*�C�){���{�(�lݴ�i gDg��0�	�3I��Oy`Aq�	���tU:e);{���
��%�lL:��`F�s�������q%����^`�
a4*��/@4,(��Rb���%����?坺&6S�i���J8#�NKMʸ�I�c��+���uǱ�Qv0�ɟp��&�ѭ���'��..���'�ǧ1m�5���:e�p�{"�7�4�Sr�.t�6�%vN�ڄE�9�Wkd�u4Ơ$�D ����d�I��eVC��y��<!k�9w��LW4��:��޺E�b�PS!�\hn+��k����<��ܛ�`��9�*���/����c��E�!�.�7X��`ͨ.����zS�5��[Kɬڎ[�qӴ	S�pf��N^�.g�c��;�&r��ݔ�=j�+ ����v�}Y`Nn�ހH��h�E��H�T�����i�Μ�M���);~�h5+;$�|��ڱޡ�n ����V:���-'s��n�Js����Y;s7���&;�{C,d<��@:\^t6ZZW|BҰ`l�[j���#KA��Ei+�9'�D�s�f���a6��������֑��)3� �8��?����a�k���OR�`���P��<.��$Ł���+�=�Y̪���i���5����~U�21�1�/m�ee�%P&�w� ���D;3J�"�Q���0�q&������%H+&7�t��w��Zb�n�Z�h\⹶I�G:�P2��`���:o��i