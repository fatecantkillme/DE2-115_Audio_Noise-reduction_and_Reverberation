��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<S��!O �&�>z��AS�:�a��L+<PR�nh��	�������r��T�h���I&�}��4�udhС�n���T�1;�tZ���E�#�x<�"c���:��i�/�-dވ�
��Z�5�	�n<�?.r��6���d&��?�܀��y!wCJ�0���D	;�v��K�hrB!ˆ8I3ջ������#b��^Z�!�ۏ<�s�9��!�Zi _w����U��p���0ڈ�o6yY�u��16�ؙS2RveCbJ���u�X�'3P�[d���K� ��w(��3o�2���T"��z�+�"akY| 2���������4h"���8��Y63A��� �W���B#�.��F�����eR*���=Z!��b7D�����c�t��E˹<[�Уc1���+� �����k�+kʈ�<(��^�W��bS�7�Q�ٛ��1}]���0b*o��N�*���{��Cw�F$ڙ�Ǆ��Zɨ�����~�E��}G!^"��`�zJ�=Y^�=O�K�!O���J@�"�S��z82û�����(��C6;8�����@�$�	t�"#~�N�Xp��ٕW����M��	!�$%�ck�l�H:�_��ԹfA@��И`�	@n�e���8�V���x�Z*آ�����a��Y<`�E��Ն�q�H�}�*� _9FO���̟=����#�!�y��|�%�H`u�W*a�	|U�Q�g�L%s������	m�4#���B:3�a��O$��&�:0��mq5��+�W��<��C�>Ëʣ �j�ɻ"�3�B�sV^�>��"-�L��� ���RJ����]�l�Φ�r�z=ӽ��hnW�o,?,�AY����1'9�����M���=��X�g���87�{�x|ǒ^�z��js�l�/���������l ��H��*�X�F�iw�F�cT^�eŎ7.څ�:������们:�Nj��q2,�/�PԼ=z��ir"����rO�ep����a����y4{ة=��d3�Q�_I�c��M��\�l~~��%?%;��0J���z���/��W�u�+`juı��������ʎ��f�Ż�hxT�#�HX���0aU�Ӵ��=@�ɂ�U��G~�o�1�'�#XnO��~�4���d>@岥���o�*��A&oӂ����M�.���K�=ă8{?f�E.��Wj��dk�?�+g�y��5�Nq����I-��֧����8()Q˖�g�(���m��7r���_(�v���*7A�_Rj<[���-��f*H��tC����)�J��\�y,(iWz� ���e����X>�tu�ظ�����ǟCȺ@OD��(���?��3�+���1W��#2�=dg�œF�\Z��㬳j^�"N�Ve��<q�:����7$k�o�� �n�ql�W+.Z��'���H�裍�@8�4�b�"�i�s�<�%�*��G������E����i,���ƧmK��J"Q�� �}��W�0K�XDܹ�iE
qyc�Q�z+��%�Y��O�6(EN����S[���=�1�T�-r���L8�#qZo��C�ڹ$�3VM�џkI��l߈Y�s/��W�1w�e��cf��Y�;����փ/�n1�,`���wب�d��써����q����쓍�7��� ���V����!W&�����<���<�N��G�ð��cȗ��0��b��[�9Y3�\�	5F�6pV�����nԡ�3�����T�3�9!�,36�;��h�ũvQ(�SKny��!��q;���;����}��%��N��Z��sW�H�j�@.��:h�|\�~#��"S� ��`'�4�*��;����|�>`�D�!���+?KT� /M}`p����h���i����R���&�IP���,ׁ��
I�q���z��aJ�I�r�]L�2�G��r�*�`���[��sr.�uP�2^�AJoJ&	�Z�c-�#Υ9���|�#�2^��@Pe�':q��q�� �ɥ���m�H��g�ڵa��#籩n*��z��hiN��N	?$L&�����)b�Z��6\��*])��U!F��r���`���q�F/9nYbVF�2m}k�=�I�}d�x�~E��2��Z�vS��_V�"���-\}�a�"�5d��%�;N����c^�c���V)�6.�<�����.��b����/s/��FC�T@9:�#`Vƣ��5���c���-$��X[�1���͕7�'~�Z-���`�8I9�R�<W3�B�HoA]�<8�Q��m��؉��MS��žl{��G��S��MY?�[����z3�Vr�W1$�Ǌl$wo�ܬ��N��'�s�{U�������V���(�8:=��0k�&���[!�2�=Z�SCaD� �A���t�.*AQ�J�1<8�����fauDd�ΰ�7�����C$ �xL���w3�_�c����[r��b�����LؼdT49����ai���ʚN"q�Dl0���(�b��Ʃ�p��ѣr��S�z�~�NYwѽDF��\2?q���)_}��1���U��^��0�<Vg�������T5ԁ�C$�^E̴�	w?P
�q:�I�4.Z�*Oϣ]6�V��1,����5�`��M���{wՍ�|NT�
Sك�r\s��`Ǐ�,d�*�����
	�������t�`�%����L��ꝡӼ ��#>*|��P�T���$�U�ؔ��j�3G�Z�֗���3cl�x�	�Z[�r��m�ѓ�NKa�"c�{zϽ��a���v?Uds�)�F�����!F4��{���1i`i����rC4XZ"�W󖬢r�Cp�����Zf��I�k�qFZ��qҴ����kP��m�TS�U��S]���K!>�_��U�֥R�TK=���ZtcH���|���ׇ�|�AK�\�eS�pה������.S��o�0���g��B[�D����e�-H�Z����[��?gݟ��%����~���m\m�H!�H
��v]R�������dM�P9���ý�IV�H���I)n����\�c��%=Q��Y���h�PPB���\��4�P�I�y�����@l	>��{CTD���!%,�]D�K���/��9��|7��2�:l(���X��_	���:gW���:�JPXA��~G�,�-��p>iMZ4,J:�������h�����Y9F����
Y�_�\43�9�.�����qY)�HS;ro�z�L��w���5C��I��4/^��sJ6�ؼs�c�s�F�C�1�=���H6>O��/�I[kG�·74:�km\��?r���d0������&_�b�:_��:�a1(D��P����3a0���\���i)�Ms9�v�B�M��9�@�4�ڔ�D'���
%�6�����P*J���M,�o+	������K�\� ��("+�U�&>x��/i	��v�/��~���lT��5MB����Ccr�$Vi��1o��2���DW��׼s	%�H�i(|oh�ʜ�58pͲ��)�$��Ī�ߤ�k�B�Rp�m}3'��|f}����܌��Pj��xR�C�Z��*2�v�j������`��|8NC �M�o�"�in���ʶ;�
#���|1p�a����*�EpxK�A@��%IC!�w�FW})��y�6V��_����N1�Y��NV`��������O+�ϧ���D9Id��:�j��8�Pv]�̸K?2d�1=x/��n5<PnO���ψ�N�}���?�LGy�t�̊ֆ�8�@!��q������'F�$�A�\��1�pz�:GJzp������r(4��9������	�Z�¶��V� ���`t>Y٥��(�D\�A�Ū_� �1�d�'�\&�J(ٸ-����32?�-Vs�׏��h����cH����d�|٩�����d�(��W�UD_��xz6q����9���P[���<.�1��Cȩ�9\Μ�4�b�q��MD�/���y��g�҈��C�ʌ�M��fX���������BA)ʼdu�;�s=�/�j_Hy.f�=:�[Ƽ�	Av� ��U���,<o-�Č��
GO�> 2����.�����ϭ��b;C���64�1�G�aMF�����̩:��ߘ���s�촋����JYv�sZ>K�)��[�H��SߧM������Rty��s�����H��-�zG�њph�#q�:=��ο�]�0���f ����;��ྮ�ƙ�᩼����*��a�XI���������SiN�Zf_D���{h�%oϡ`�RJ�%X�F;���}�ŪT��F�P{;��)��Rn�%?1𚱯���_L.�(�Z#}�~9��m�=a�����A3������>��ߡ��7K|�g���i��l��k��-N@n��n(L*�r&�oD�c���R�k�$ڢ���<�:X������w x��׎����.!�F^�,�Aڐ ��r��6��Z�J]xD8��pk|{Ѫ�?ʵ�m����p/2h�,q;&\k�F��.e��t���Gm6;�A�.�]�dQe<g-Ya��q�����3w<�.������iz7x�!mǵ�Qo��f�I�B����VA$e8G[\ ��:Y:����J�My�s,���n�i��}���B�d���F#_#w��)�Q3(8�D(�MT
@r���pз˹'JC�<gXMn'{��X������c�59��<g{X�+S����q��]9q�@��x������)���39�3���T|[�O�Pʍ-d�}9�3v×P�(�v�����ʀ�mW �r\��b����y�v����X��P�r<��� h�=���wJq��RZV�yZ.,�P(}3j��V��Ӂ�?;n5��F�S�D!�cD�$�tˉ�jW�#~��m�����Ht��;��P�15�&���cXԗm�n�A&t_��n���"RY�����-�z�����o��=y��/͞u_�;��i�L�v�`�>�\��9� E6�������=� �����e���<,J������I􎉓��ϼ"�6(��8�i����-z'��+�����p���͜�`A�����o����ۿ@�z����!�[�m�ǩ�w��Փ1!���U`ݵ�MA�-�L��l"}�*���"���A!�=�Y
�s������h�I9���f�v����c�J�P�@L�m����!~b�O7����4B?���NV��%d~��q�/[/P6�s�5]�۾3Ե*��+��T��{,�#j��ط�S�ESt��B�=@��p���rg!:)�o��	�Jo����Q�<�n$����햫�)��c��f�+��O8�tǫbn Ƹ�r��� I#����2�bvR!N��|G�����_�A@�M���c�η�cw�<I���e�ֿY�^�
}b}��iaz$����(ߐV�M�7���7��a����lк�0�Wg�`��I���>���IT��\�����D��G;{��y��f�3��6bs����DŃg\O�=~���;�5&�^i�Q�z��ɳ��q��՛+�4�Z�z-��?�E�ֲ�^}��y�ay�bj��M���+7���J���h�dL+�p9`d�ؖ��a��3��/o~�s��)߲_��-,S�s���(Ӗ1��UL�xq�G�����UN��;P��mQ�S����:n���ҳ���iB;N$�<��S����/�0��P�c�i��1�dw���,֪������N���v��[Q9�OLͭS�w4Pr+&Y���dO �ya���ϢZM�P���Q��}E�X�s�*�c�}�m����s�����ރ�۳LB�#�stc����x��R�g���@��8�%��K.CJ��Wɨe��e����	���j���T�:���7��W�q�H9l�P@r��@�c���^�V�/a�O+���/?~NI���%���'Sޖ̘����ұ�+T#ӗU�^��k؇4�Dn�{渎-��1�|��}9� ��~qqӧT��B��5xV����!!�.�z=[��VA;X5����s�/�~C�s
F+=��1��h�Na��٫R�u�q��ŵ[�|ӇK���7�5�Ʀ�{RyX�.zߎ��Np�Ï�
'Nj�B]����q0&Kd4j����֊����Z^��}��
�T�@9�- ]�|f�ƩE�g��,��+>��������a�>��a�r.ZZ��[SQ�h�����1(���n�.�И�K����dXb������&��; >�yrR�P�8z�f�!I"�iR;l��wq����%�tz\�������"�l��*�J�g��&9N�1���.�G��Y
�[t�?%dh�
��5IK渨�w�M����	�̨6EDvݦ�m��Q5�OVh�n��x�	�j�=ېf|-߬��^,�jt2�:���	sR��<���qrk�Cv!�G�xJ  0,Ą�/�+�7ha�����;�X{�s�U�k�¡+���X���������9p��fRȌ�/e�{�I� �q���pg�Z6�]3I�n���7��!�����<��<���$�YM��'3 �� �vz_����G��������ҊÇG �)u�k=- �X����HP�E�0��?��1]kCSn[P�K��E�VX�jD�fW<��5*��{O�`����[/;�8�X>6�v:��%��X��
��x��p>�rbWN1~9\@�0�I<=]=�>��y����:��e������oO2��lyD|�pm;�K���Ռ���юr*Y}g3u��J�<����@�\�<�����Q�M��)�Ez"�wc)H-X^ϑ�B"n�g޶��~��c��ԄB���I�1hr+-�&mHZ��i�}���jp�)�i���( 2�TZ�yA�*��<J�>�w�{Ju���$n�J��~�4,� ��?H���������TX�霿;o�����Hfb��x�W�񸸮*���s4���tT��49�8¥{q�S����~�kY[��	��fIBϫg�"��� X`�r��9�W~���\�+����vS�'�ģ;��=���" E�Ǆ�k~�I婄���俁}���4H&���|�ݢ�8����\O`���:�n��Y�Bz���F��oR��,Պ5�MKd.Y($	֞����;)�2���<R�7L�.Ak+�M�z���T)���
k��#���v�7�SN�m&�\;��"^��J�����w�S1 �z���W��_@mBይ���B������q��E�I̷��,�~P��!��
�X�z��c�7��	P��Y��7��$\*2�'"r3T�>�#�,��B�c�G�X��>y���D]��`p����|��/�#\d��4��N��~}��,�xͧN���:;?�����	mk̲C��(�g�ԏ͛<�v�S���������'(Q�>�F=�m�O���P!�E��<=�L�?l���� �G4�m�G�U�ǡd?ؿREe䒜'$n��3����f��e&�zlEae��B��1�@����gmc��k|j�ζQ��A��.��GU��kX*I��W�"�}MCj�m�,���ŉ�!'���ߗ����#ذ������W���!/M�J�iNҖI�}wjƘ���TǕQ�� ���\p�߲�m��~iZ�<5��0(=-�'9mm�dF�6[>�HS�*���;��%>L�b)0q���p$V��td� �h:+��Tɉ���͵~���Oӣ8���}��ueK�Y��7v��d+]-�2"`��2|gf�K�:]w��:���?�c�k�xe
+�'�G�Q,�b�[x�����9�;��_����.f��F,��}�3���z�$sq�1]q��A�j4��p�܁�͏�s�����9w#�ǉMM���z��]��T�<��z���Ӓ^֖d7X�R[2|5���H4�'N���1��M5h-r;��t|}� ���e��]o\�� ���7���J%ע����^+�w	(�χ�v\���@�tB�.W5[��f����Ld򜸒Q�<���p*m�[N�&���(䪶���e�S�ag���ȁ������(�-U��Dp$mV�אw쫌�M���p��s,:O������RY��CbS��Z-�������%����]�D��Uh�i�[���@q�(�*M�L.�a�o�s�;�P��q�L&n�߉�P?�Z�Y�5�E2�Z~�_"�#D���Z#�v'p��(ă�;z`�$�C��a�1�kF��!�]�+��%'�0�=��P�l�;�7���hS���p�\�n/5��/��]�s�[[�/Jg|��HX��_fiV�-Dڋ�Y�����Q��pxP��a0��Q���ل�2�*]���$03�;��*� �fS��Љ/��S�+# �؃��������ӈ��j�$#~�>�S�29o����y�\�)^f9/_!���+�c�@W>���QKP��`w(Hj*f�nhRj��'Eʡ�^u2���o�[�r�Y)���Q��d�v5 �r�	s_�pȅ�P	Ma4�!H�9ED�QӍ%r���޾x�{}mD<��νQ�ө���(/DB��fp��d9,��0Ἂ*5,�� 4��ؕ�0͒$�����͙G]��j:fy����6���M:n��#�����Pt�j�#|b),u�3j�I9�؂����q��x��n�! 
�X��P�I���" ����C)���k���|=p��n����g-�b�闭�y�Ǚ�e��:�V\'"�'�Ct��mޔ��J'7T^\�g�zff����c|ʙv#q;��eJ���gP�;�5Ⱥ�SuM�����{ Q �EW�U���Z�ѯ)��A Y�f��\9��XR�~1+% ���E�g	�}��t��a���e���XC�Z�^z����'Y^t���MN��;N(`C
x��h�;:ET��͍���>��s�?��b3xX)���< ��H�voU�)�����]bj�u!�G'����g ���R����V'%]��a&A����H��o/�J�!;�Z6��yb=ebb-��4;�������yH-{�).ll��8�}R�<KT����-
���
�����O��Z'���m4O����=�"US;HS#�_~S�K�ɉ)�n�H���j�����M�k�O�P�i�4{Oٟn���> �N5pbH�����mQ W���
�<n�}s�O�5���25���{���eV`fYv�Z��V��������I��p�]�O��x�o��sE�ǜ�S�5�K�ϊH[���'~7R&����+#<���8v���nj�Ȟ@d��-� ��ͥ_����+C��$�_����uf"l�ZYj��P��#���/�f���q��n��w��ԑ�1���L���1���nq(��r��՗"K��/�k� �uDl���!�,�"D�f�qg����k�s��Va���b9͂#�Rr�/�ڠ��(�Ɗ�ՓňJk����,��n�D�+��o�x��&����Yk���oGA0z}^�0/�-�vbQ���Z�\�6�ѐ$7��]BG;.GT��U���JBM�c�!;�{n�E��V	.0E�S���j����KG��w�����E��d��:��H(����J��,\��L�����b�z�U���^��av��9���s�)'���\/�.�6Ih-^��/^(C�y��8M=�x&Q�F�eX�16���N#1�LQ����a���H�R�g��#	L���j|>?YG�7Ng�_����|ŧ}jw�8�`Kdi�� r��"��cP���SV�Y��4��Fg��%7S�VS��%�Ƥ�-���2����a�9��q�.����ZB~1aw�\
�.;�4����,������GD����:0I�]�+���X��܊��i�d�sb�z�GK���)ÅƇWO�nk�(���\g�c���냥��,ǣ���X_�A~Vp)f�tԠv~w�&��.��S�.Zg^}^��<=<d9F�'8�>���������ݚ���u�Eٳ4�#���y��K�&�4�z"<����gw�N+%�_�&���@բ�6�M.>$u|��o�o}�P��ҩ��׮r��h�ؕ�D&��*�OG��Հ������Yvظ �O�	��� D��0_k�)����vxx��}t���|$������Iΰ�;�݋����:|�(��O|��.�A�h��TX0��ڙD�L���-�/J��R���ҭ罹x�2x�>H�P�D�B�u�-d���K�_qP�Uot��,H�����°#�W�i�ԟ�o��φB��o���8-��J���D�"wJ�H�Ic$�#�?�� (λ�ٗuB-�0�'�J�4��6|l�������*(�ƹX����?}bÿ��g���8;B�"L� �PJ|�?�#�l�<Lu�nX��V!/���2C�l�	�Ab��ި����6"~~��O=[0q��ݘ+Ĳ�6�u��?��m��/�����$�@��rf;�D����Kc'�bcM8R��S�JD��P�	�i�D��D��
�����@�(`�܀#>��ߵe� ��ϩ�>U��B��T�3=���&�\��N
���_G{�ƒ�<ɷ��$��Uni�xZ��i	��.ǭ�<u#��˱��ғ�pOs6�uD22p����X{��@�i/e�Mw�:��h�[���ї03	��H��$Cx�W�q�@_X��'P�ͮ|��e��a�����;_(on{���F.'Qd��b��i�f�]u�6�Uz(�3i�;!�l�B�JM�L���!�G1����?5�(r���Z���O��)�:�(E=�~�,̨�+�0Er�����U3R��v1u�ft�$�l��(t��/�B�'��?|��]�_��1בe"Q1�#�X{�����U{�V5�c`�M��6iu��-hX%����bH9��n�D�*�dY�Xǡ®� ��I�`�I��b�&cϔml��[p����MQ�Ah��V|�=�������^��t`D�A��TW;)�04{V�jR�_x$��T�,������e�f@��e`P�<w�~?�l�_�B��\H���^u�Z��c"��<�l��iҌ��eN�|˖�Q��묙­:�W�X�����	��r���9���W2J��[��D(���^<|�k1�M��LY��8������7��b��Df�D�~Q�h��Ńd!i��m8,N7���_��WH!M�9~����(6ּ(����CT��<8����j��`ȇ�?���^u%IP���9&���MS�e2������u�1m��+�!�@5�W� T�c���y��!��c$��4���8�|@�@<2
H�d���Q�Up������u�щ��钲K�͇�r�YƉ��!�B��&��x�@��苜���BOS������뀜��������	� d����1��!e
}V�����x�N��*�޻PxVE�pj�^��a��A��|rĘ�r�&?S�M���f�Ќ���Sf�cǩ�	����C"�C��&I>
�Qc�ϫ�8Gd��W��5�ڲ?�Kü���e �b
�T��RӞ��#L^�B|�an�?>�*1y�HQ�"�g^;������(�S�.w�v5a'�f��d�]��Ą+��lj�k���P�֋8D�]˺#����IM8֘[E����yXŨG'z�K,�����g�0�N6�e�+����1;B@����S�`t�ԣ���UH���Ik�gR@�ͩ�,�a72;'�m�;>n����u�	�W��})����k�o�iꂲm���SRr5f$�E�ُ\���9@��}ɰ�@wL)ء�}�K�}��R�oko:}[1��2S�����9��r�-�4�;��s�4-4�:��p�O�@@����	�ju0�Φ D�{�rWL�>C��1::�>G3d+���?Ge�D�?�1���F��o��B�`�5��3�� �E��N�����b��I�՟�oz����бۚQ�|������Zҳ�B�˖j5I�~�swt6~�P�+������I]N��`�x'mP�?3ϐ��R��
��U��ԽӋ%��~u�t�Q����SL&0��S���xN�j��q|l>m���%�T�z&BO���VYvuV3�䓻���X6�W>i��h��T�6X]����v�v��,=��,�~(�`<vN����$q�fu�b���h�0��hgm9P�-ܛ4���������P�@�~5�b�3��|b|�@�tS�K�Dni�t���.u���3`��r*��{��^`�-�K&�*�bZvђ0�8�Л�Tq�թ�7�5�^\fSR�s	1 ]�͘����Œ�1Se�K��-Nr�`<	��5��\��EfiͿN��|��G�OU���
'Zp[X+A�=� e�o˘Ҝ������'�"r�:;n� ���n���K��*RqwZ!��B� �eֺ@���Ūg�f��V	���
��ŉr�;��3��n�R2�{c	�3'���}l;�@�QRC/��Y����I(3���3>��%@�kq�/��-�z�<,~��: ]Wc�����XC��~�����F���yє��QH�^̕s�w)�T!=�hs�k]�1��)4��)��"R6����|ek���t)2�P�d�R\v�C���x'�5�i�:2�I��oͮ��e��}u�
�9��"t��v�f�)�Fok�1_Xo)�C�Sĝ�:|���u�.�Ѡu`����^��6;��ZЄ�Q G�	�I� +4I�Y0K�H�G��~�S}�`$���.W�M�x������Ъ�����i]��6Vr�w]~_j�_y>Vf��w�+sIg�&`MtĮ���IA��q�Y��|<��z��P��b�yD���X���ya��,��I�EN�Ϗx�»F�C���FQPU�9'z��?!��Hb����d�K�(���w��e���$�C�j�}�t��^�R��(�'J�Xk�l�Z#��y������B��$�_��!��%1�ݝn*g�ΘsZ�������Tv8".U&W�}����wN�.�=w��:�?�8*��ڑ.b�/@$���	��������oKJ)��8�J��tic��H�] \��唜M�v�xl�ॏ���7X�v��B�.+�e�iv��I�~�0r�W�B�>b{�1�A,}��2C/2r�P:�M6U����'ΉvJ.��|�֦7ƺ`h�<�0)�nME����� ���Cu4@��b�ѭ@�W��L���4���c��O}Rc���G�TM
���6�3�������Ӫ�<	Q��7��>HHݤ��2t�H�q9�AՁ�J\$Hf9U�x����%Y^ub�Duc�u��H��E���sptrT�����^�*�9��'���i?\��		���I�s��#���P\����?��$]��}��:C �M�.[��������d��+I*�랮�ZH��w��)=��!�' �<�i��=�Z/�_SW=���<�U7�7{��&e�`�����*GjM 0LZ�BG�ZV����%�������U�S
���������}���j;5����;ĉ���ױ+�O$����Z�C	b�-j/z���� �U�)����/}D�~���ޛ�aȵ�|I��{I;�\���4;&���g(#'�^S��RЕ�V/�trLN�+ �Z�}�|�A����PK�ӥg�,���0��7�����Y�d����|Q� �a?�iE\�Ow�*��A�P*����Mo�$E.�Kq�`��ob&�d�C0h�?������_V����4��:A�8sA|y��T�{-�+�ԶІ�3N�]d�=O�]֬NH3��}[Ƞ�����'Fj���s��m��3��8�4Z���.�F�+_G:2M;Kdt�r�����Pɓ��CT�l�<�s���Y�c�4<G�d=�$�p�Ln�.��|�<��"�k�_����-Ӣ��֓�u����o	���K�vM�l�{��k��H�[��M\:��^S�V����O��Z�}�+ Q��'�oN�xH׉��;������%(��_"ʣJ�$�Cˡ���UoQ��kx�^ޑ���iaN�JDbhD%O��WGk�9�^ٱqaQ:7�6t>�'5��hp��b��
��ZD[l���a����$�����ܜ2�&{���i��6�I�w;~t�6w]{����"T������ $㿃E5O�*�#���r��yH#ʬ����R�9L�9�!���}*��̄4�O�=�!��(r$ɩA��3�<{[���敵qV3����A��,�H��C5h:O��0����*�q �BJ���z��bV�3S'�JEX#"���LH�v%���PER�l��s뱝��s�f�A+ϐ0��Կz-0e�TL\Tˬ���1�b������E^a�Bws��r÷fm�%.�?�Ex`���B�snT��� ';���E8�k���-�a��ﳱ�u�'Bh��}�d8���7�� �T3������ḫSە�om#Y��??z6�{DĿL
����x����GZʐ��ͅn���r�֜&g�����z�����1��۹s~��J��K<�co����M�,4 �[���^ w˙戓q��	�@���`���ڥ�xn��I�֬�}χ&���ʟ|�Zjj ɘ��I�N��\�aV�v�R�nbh����-��d�c�}��Ta�@yf�BP��Meb��#����S��E�kzE���5��]�Jŧb7uC���$�Ұ�D��i �L��Ʀ���q��H{_����_{�ܟYۈ�[�Ă2ţU��E�吲�F��<v�V�Y�1ڶ�Ί�y�+뵇�����WZ�W�S5<�����P�D��QR�85;s���fK��;Dg�F͇Y�^@���~)���������+G�9��F�h���7�wԺ�Hd�+R�dZ����hI?�߯l(���R�Kn���t�n�P���`ΐ�����g�p�5�酿%Q�#� tZ��z#�(Oѱ��О��δ�$1ƕJ!��!���oB�0�P��2*�XJx�甅���?]�UC�zx�Ѷ �a�M<�0���2BP����!�^AU�*�Kb�>z��	X�1�.b�c� _ ��oR���z�*~`�RL#t� �a�0�1���~��� *Œ��M���Md�"9%�X��#�EյDd��N��@3�S�w�p{��V_��RK�� =Jea��bVNp(�,�A��� c�1�rY+�����Z���i��lGt��o[6���`����`1
Z�ڣ,u����!N���NXz+�� q��'�a~��ޮ9�t�0q�^ʃ��C�M��1;�*GE_BE"v:�Z��\R�ꇴ!�x���y�rEn�x��Yx�&�W�(`�G��p��0�`B}�<w� �Fկf�Hx�.��B���
6R�;�e�{�@�sT�hf�3Y��pafv5���u��H�܃���S�S�$*{-�\�?���Z[�����4����kɊ�D�5�U���i��ǁ�ʝz�1�?+�$�#��ҹ��s7-���5��g$���:,�������iS_8:�o#�]w *�G
�aOk8],9˳�=*iUx4�
v-e\��fi�UI9}�B�K�B��@|,K=�"jG��<$��$X��K
ӂ� ��_	������39��2�j�Vh�6I�L�A��{,�7}me<F�%�� ꒕#����]	�5��_ʊl,��6�Zj%
ypQ�j)�u<D<��у-ua����bK���gL�:Z�vz	^(O����0�x�a�đ�Q�'
������У�f&W�$Ev�\�+��X!%FZ\�>-�-N:��z��t �4��##�OV݅͢��'�e��G&V��Yҝ�T�
�(Ye�Jx�A�UE�g�U,�PsG�P����t�\�Q>�t	����.ca�l��zW��Ƅ�>qxc
�/r�"ߥ�1�%.���5f��7�/?.D����lנ=�`�F�<�� `v����V����� �7]A�t\��vAE7����x��/��){YpL�N�ߣ�(Q�s	�V�����(��H��Lu Ma(��}(�Q�����7��T9%V�5���:Q�҈�KI�#�;�[_�򆮠�&K3���.b�(�L�XW���ǸE+�,��oI��=���5�ܠ�y<~�5[�+焯T�.zC�z��/�~X�x�6��n�6˾��|U��;��-��/Q�1������*A'�oG��G\~("\]x[&�:�6/ɸ����v�|uTԑ�n����o���Loz���ܟmȉ�Gcow�OG�/�,Εx��������,�"[�T��t�5������M�P]�/]�����y���TiJ���<��$́��fZ�.��V�\�˛�7˸�ho�'��)=�,������� Sȫ�j`��/6Ө�u�&�_d�؀�f~�҄�<���ҦZJSb�B8�S���_�Yo���>eU.���U���νsm��mZ��Bu�M������'V�E|CbH�콘�X<���.3NVr��7l�iYi��12^��Mm�mO��m܏�q�1z�{<���zq��ɓ�mW���8"�,*����oO��0���(������F���D���_-_� d�5��jW崿��ە8Ңmw�Wx����^h��Cy���ӏ���,B;���I�P
1�if�U���?	���Ƴ��
Įc�ڰ��8u��T��+�m��A��IT��'�D�J�:g����6L�"5����.�?Q��.����_�bU_$@LB��Q-�Ӯ�����OQ���+9z���Ƅ�̂P���wǛ��(J"'j��5��RƟ�J��{�MH�8O�>��+cn��@HU˕B������Vm�Ȋ^������n�f��D��h��Y�����9��U �����:\���Yi�ֆC��݃$�n���@h��[^�Ŏ�y��i*;7����k(F��}�C����up+�V�����^Ǣ0dپ���u	����`���P���wܜ�`;�D2�C]V��.Plz_"����O�$�Gj��Hʳ2i�>��/}7&럗rj���Kb~��2"	ӾR"B��<"�X<�V�8�؜���%���
�j�\����)K�"�1�d󽛔�q���������j�,'�0A��T�|'ؑ˝R	�˘ �in)Ʃ��#ʾ%j�kv,�tb�GAs���by/D�Q�D�o�k�$G%oݬN9�<5py^)��~)�ɯ�6�E�í+�y���s65�]Z�Y����*�4�����I2�Bg*��j�Ȏ�[6����z���������~&�<�2��_V~D�GA@|T����?:u�#� _��
�~\���zv�Q��c��T��흭&G�e��7��#X�����>�-�g�𓑿- ��|z�����6��~e� �K�]��Ϊ%�1�в�!Ȫ�:����Ͻڃ6
n���	9he�=�?����Ѧ����z��Ә��왺\1jF�K:Ϭ}	)��x0;�5���L���2/��a�Ӟ��*�c��J�`~Q2��@��K}A�J��o�y8�ۓ�ګѩ�t��������{�pSW�r|Q�`_���7�.D�pe�B��w����:4x���{F�9ֹs,Z�B� ���}�2�I�H�K����I�(�ǧp�f�L� _D��#���N��_P3�B�5ݒ=wXCd��tX�O���MD�����J#̗�/�Dേ���7��Cz7wI���ܬ)~�0ڙ:�Sa��9�o�"b���KR�64,���%LcM��@3�}�HK�D�,8AX#��~G9��Ν��3�)��Pwͧ3�e�*�.
8~��{��0a��g�R>�*�3�|�גgcr�(q���_$,��$KN[�h���9'\<�Đ��a�8�y�&_�O��F,M�8�����C��"7�h�Ǌ\�A����BT�.����'�8ZtM�R�J���)kxO��DE��&�+O��6�7�4�� ^]�kz+���ї�#a^���EsR
k%�v���3���o��BU��%�0hW[�xO�{�����FG	�~�u6[��ݫ�c�b�)�W[Br �hME���|x>����n1����mg��"!%��Yі��Y��p�� �|��@����Oo�纔{(�㓟�I��XU�U�4g+U]�n	J���>�k?���b��A"�ٺ���<	iӚ���p-ot�s�XB�f�T[j���C�
��I�W�K��)�%����:��)eSe�M�X��/b�q_���%�k�׀t�i�$ƽ���8���A�����F��TI�\�s'Y�s�	G[�[�g�&6�<ݰo֛,���PpO���5>*�h���o�A���N�~��f\�O��x(Z����0]�O��ES��l�OS�F"�V�c��^�Z���3~yX`i��]p�R���їE �r�n&U9cCA=���IͿ�X,r�H�8�p����ޟՆ��m�]9��i28V��O�P�qu����>񒱄��m]�� ?ƫxE�aY�!�ٗ(��&5 *P�������6qx���s!�΢��Aʿ�5a8�|�`�u;JcFY|"s�Z	�	��N�̑�2� }�g����2��@O���@;!i������l::z{��)�|;��:^ؚ3<�:�wd�Mn���b�������B3Í��ĽȖ�e�4 o�����:��0 ��$�h����HL�5�`��W�+YH��|)�Ҏ0�}J+�n���&�@I�)�+��T�"5�aZ	!�(b����;5R�\+k�C��"�[���c�Ь�8%�T�F&�un�Q��IP������U�4e����	�p������ﮆL�􎚢7�W���[�@�?(	,9=���λ\��wȆ ��2$��P����XZT�B� M˺\f�H2ٵ&���z�ɐ�2�0[S��\����fE�����&.$��w����(K�"NT�7�m�ٜS3�1tCQ��}�;"ڹ�-� �%�A�2{�3�����J����Y�R+��NA���z�����n�+�˨��g�p�x3:v�IX������XK�a{����5��j��>������wK���Ki偬_%�����P�pڎǫԡ��p_7�� ��^���.h���~�����Q����2� Ж�е��
�����;Eޓº\�1[A��֖Ige�I���%�O�����q���b*h��ɲU��r��b{��݈Rg��2oF��`х��ﭳ����;����tQ�?���>8���͗�|v�^5�=����a�)��)�� ���"Wz���n�E���9�5�gK�}t�f]i��F
�tw�
���V�>��l(��S��9�����`�ۺG���Qԅ4l?�a�6�5c�7og��giv�^�N�X�=d}E��"��|�Q�,�#B�����%�S�� ��ӆn|��A�����'"��i�d�y�sG�j�*�|Q��څ�Y��ƽ�F
��P��A-��O���qF��&q�G'�|4���,��VҰ��u�'��caR����u<�`��`,hg��{��÷�F�K�tN"�	ώT�+��|�VN�^�s&�s4Wkn�G<�[����;Q��	�T�w;�X�1m�4��=�a�^?8,�c��^��ǭ��Z	�F��t���)��X�`2q�N�5��$�<�Q�j�D�N�ʖi6F��Qd*���r����*�CkJ5d��鍻��&Ayz�
t�|t�*�X�&/Iù����i�	%�zQ��a�-j���*�y��ĐL�"�[Wń�,�B�8
c`�SI'3�d�q�9�fn���6P�R��Z�'f$w�/h�@���ş�:�B��S��4�{#����7����4_
�T4׆��O���(���/�|����eU��{���F0M�5�φY�8������M��RN%T���Q����j�9K�WM�ka��w�i��H���D��g�YC#��%��.? N�n	!`�˰��WϜ��T̴��=*&���t9�.|��F��Q�.v�)2��]�=��q\E��X��{��H!��#X��j�93l���`��-��񛚏�;hf��|�A�GV%6���	=�}�0U�k9T��� �R�H���_�����6�E(�SoNn��I�.k�NL-w�H��K5�6���NZ]������E}��Q��c.��d�Vh��Ĝ�Iy�����/��Qb2����ဵb'�s�LcT�2�-��aפ��.�`�UGrk�U��G��?��.J��v�l���e xU��RDŌa��xM�^��P���6H>-�SI핅�;� 6�p.�E�=�`/�"yhc�u��+�@�a���U���7g(��EGt<Q}��Ǹ�ᒍ� |~pa�R,i�������z	{�-!_d����@�Ev��_ܸ&��_������@RB�� A_�W+��V��:/D��E��c��UI� k�Q����z���˷ԍ��Bċpo2����s5���Z�7j3lX�e\�����!��*U~�`����P�2�p46S���*�S���ʃD�Va&�o[5=��'�J�x���
�՜��ݩ֠M�<]e���j�6 R5a������5תE��݊�e���ƑB?��%�x#�#0ٔߪ���O[E�@�k�������T
n~ꑏ�_1g��%�T�++F�=ɍݜ�Y{"8��������Z��(YZ��bZ�PЅ���k��K�w� ��uY?҅��/ԫmH}��Z��"$�P��5���TF������!�9&�JXf�)2T+*]ն{��ό�ț��L��}C���3���Y�p`m{�N)L�[����lIi9t�2�U���:�����x"S��9������yU��׍����0�q�;��a�\�#��x��q%7}C `��y��ʾ��im6�ǥ_8��CY{YM+s�x�a�~4)�W�}�n�����5��U�q�D�(���-��u2����`���U��N�Q!��z^j���,����W�YL1k�%(�;��tcF�U"X�aD��O����a?!b�>0�n���֠�G�����8���M<�;o� RΡ� !��u��D���?�Oپ�,	A��@��\�p�|��<�13;x��׽Z=v�$\��m��
2�d�ZH�Õ���^\S��̩$Yq�-�����m�4�5AS�μN~B�ʝ�y	�d���Y�O�^֔M�r���}�;��<��c<叱�Y�j�t�,�o��а#������������R�(aJ@�O\	ǖ���<`d�d���UxRE�^DB�� �n��������b@\ã�V���Ѯq �-�QC�����mE�Y��}[�{S����p刯�h��۠d\#��bNp��������U����P���G�楋����|�������^������&{�O$ױz[Vn��J�}�x�ʌ��7���zM7�f%��x�)�Cf�j^65'l�\K�C��H�N�/��:���Ad�çj3�E�������*Dm�TrH�)��@���P[����C?N��Z[��"�Z�Rq��`y����;��.�����;�֘װZ��xp�h�F[t
GuN'�Bd�������Gr;}�X�\�'�<8U�=g�ª��>R�TZ�qIff�"~/l����������U}܈Mq�������{�]�l`���>�!Jt��y��4�s�5�:��ڙ��`�Ɠ*]��pD�Qָ��P�敌 B���D~��=��E{9z�8K���^��s�	t|~�D�D�������Wd��udxk�=�Y��Q�����V�|��)��T���ޒ����S��wg�A5��?�ኝ���ɨ�)���m�f3�<p�UM�"i��6���\:I���M�U�#uM��S|�a�:Q_��j��Y�P��Y��⨀��vw��V2�q)���&C/@�M��e�O����W>{r���/�Ը�R�v]����d$w�d��q&�]�c1��ڞX�G��Y4�;���F��iq�{�;#�M��Tʄu9ee�a�p�ö�Q�Ж�����H�N�[���|}� �" �(��l�^h��`N���I[�Ͻh?l���,NC]�-�[��^�{�+&P*��N"������2Ђ��¼H��d<W�D4Z��}��֯{����©-9cN�F����E���,'*���"?ŋ,q7O��{�c��J�{�:Q�8j��֒�o^��}�s�W���4�ۻ�\,�`-<Fb�H��1��
V��0�W+�5��4����9�#s�z07ԡ@oU���:�t�4J �\ ��/R�T��X��*�,�d锖�O��=��Dy�k��=�lx�څ���9�9��/�{Oy��Z�l�Ӡ�Pl�����o�)||���%O�f�7�4�&Կ�BD��bO�X���U2�Tk����-�z�?�-ԥ��}D�H`w�D�8��d�U�F]���o�1���������
`��j��o��p���E��<K���w޼sN3$3[eo+�H}w	�"���óqcֈ���r���t��H(,������~o �%�jn�M�QʀGҐ��5!�da���Q��?�� �� ��i�[�d�EE������ĕ���o��*�������.)!��Y���@�/?�Ƹ{�9ڴ'+ZH���y��:�GK�a�نj(�]f������Z4u���x$�Ĝ��_�txiN�$��S/�cH|����LXb7/_&Irꝰ�����U�W��Y�K�U)�c��?j������[��P�`v���=nc5�aލg���@N�P�l�وI���b%f�d����-Y$���A�w�޹܀/��^���pɴ���Q\�h�9�!	�e��5��/�-;)�O gh��~�{�����ri��G��	�����t3��KN.��21��UV�Jb�X�S�B�J���g�l�'�	ڣV�_�}{C[f�L�����kn����ac`�V��0K�瓡�a�$��E`�����Uq�`�J�6�����{WaC�4��r}�RGq��5=\���W~����>�ۢ"���*���=�������"!�/GLwo����H��q��U��׋��LL(��eL�i���r�I��pr$4M�OrH��GF
��k$v��JX��,`��wq�V!����o�%�m�Qe�j/p�KC`����g�����)A�����}�|rm�4C>w�Vp@pp�s�-9�#�3;wV/�]������+����N���@�ՕIjp���[�n�H>�7��f0�����<~S]_�6i.�bH4�MʪZ(��H��}F_ʾ� �����m{4��Һ3i�gY�UU������%�F����I�1b2�s+��Qs���蜜d$Jǯ��j&�nM�-xd@!�����W���eK��
��):H��R�b�l�g�����'GR�xz@�o���,۞�c���`yU*㾟�Eӕ����~j�a`w/�Q�|�H�>-;�{��1����ڣ�7u�vC���m1�J�H��<�q�Wq�<M��ᱹ�-���=DcJc
k�^��R�v��_�0V��d�4���p����wkw���
�jSo�Qc��DҩV��	�~qM�1AnD��I���~�݈�g�9Q�އ �"K?�`J��o�w��Ը�F��6��t3 ��@��I8��u?K���?��e�S�2�������be\M�*v�#��'@d/�g4z~��.��k�n�3c���o���,� agh��%}f^6]��Q~���>,�|�q�WW�=�s���D�#̪-�##`��q~K�zZ��ܾ>��� �-�Q��a�%���G���nZu��XH�ɘ����P�+�oճ��}����g��ӎ3�r��Gf�㶀T�X���q2P�;&���{�/)�,�Nm	tb��1��`̖Kl	'z�n��x��%�ſ���,2�,{Ep,�;����_���u��?�@�Vq�NZ�s0.p�e%!�b� %��G��T@憩[�2|� 
������,.��ڧ��� ?�
-㕍<2�� ��Q��r�P2��S��2��a����Yfϫ��i��UYW)h3>�hC��u��G&w����l-#�W6zO,Y��l�)q6}�f�7{BQ��%���߀��?Hp*\P,ǢS��������<3Tź��y���;�,�w�k�F���p��.�JCg0�8��߽�!�r6�r�i��:㬠���-�Qe��o2�~Q8��N�}���~UV���+�۸$I�bs����_��q���1?������p��0[Щ3s/���p���"��(���;��c�i�:���x�|�4JTm�U4�a�	�Y1���'V�z��P���٠gMo�yNY�AAOӞA��~��Hg�Ɔ�Oj7o'�MI������D��kOѠA���,���譡�����ů{�T�F (&��=������\�Q19���w��.�cb��)���f^3���2��	ݱ������Ȕ��J�F�j���hw�J:1�j�r��{G O]�N��\U�����M� ��`�	�o�oYj��I��3AS?����1��e�pʻ��sRJ�-�U���PN�\葳�Z�$8B�PJb�S��=���kk����*ejW�∫�l������pX��U7�⌘,oF�.Oa#�}Lޖ��ʤ]y�/�,9g�R+��9|��T%N&>a���s�;I�P��*|�jiZ)x��(�?#��mo����~��n�T?�X�p��9��?BD��kZ��`��>�f�C���w6��5a�;^1�t�!�4��B�	ں���w����]H]�����_|�G9����5ܱ\��ꪀ����r�v�Ua�SK�G��o�<�K�!^ro�-���<q��L*�Tk�L�6��W�e�+~>���Du�6Y��ؗ�Ӣ��U�z���[�)MD1�#N�{%��ࣁL١O�i�Oe[�e�J���2��bmk��d�蓽�[��O.T]]��c��yK��4��Yk
��#J�����Jn7NuCO@�����=2�F��]�if��7�,������\���Fm�9�f�`xV�Lf)?k)f-�h��4��*�%G�L��D��B�0/�gϾ7e�+�Ѯ^�۵'��˘�%���m��U�I9z�ƺ��ܰt
cO��.���1�<�R����`e��{�$UR�DO��� 	��w֕�X-��У�5#ffO5ȡ�x�M�`gv�!�O�vŇ	�]"�/Y��Ko����³qJ�-����pB�����w�)jڡ
*�fĜ�}?Ru�,^Ł_��ʐЗ�l���/��-3; Y�|�����4�W��Op!ȉ�����s�����R���q��$�	�{�H���6��֩X�8�%��dG�?�"K��IGeDz�t����a��\�^��$v#�����V�ay�����27�z+KfG}�s�-j\8	
C��I��'�D�����fdT���=� 1��S��{�ɡv����Z)�-��T8�"&�r�B[�� ���vK�=�}@*�S�k?�J�wu�c�n'���	y)��7ʎ>��I�,�6�c����|-�-3�e��),L%C�@�,9�LfQJ��y ��<��V<�1ÂD�J�D�+���-ea^u���@���4�w�x�s�e�e&����0�YƂ�Н���Y2�F򵦝���,��ذP�7�QU7&��?��{\�X�y�����}�"�-Z�8:�����V�Lo�T���ru�������Sմz`�#�B�M,*0��2��qqw9�P�K��9��E��H mrO2ye�ZݸuI]g�<�����B�x_��}9�P�j��mQޥƽH\�o~�`��n�lT�7�f�A$I������ �v��������F'.��36��/�����T&�sQn�2ȭ���96�XE�Ā�W���p -��74~x�����ۦ�#��
��O��Ag`$툝)����7�8�G���a����|��P`����80�X�q�	)��3IV��n��z_܍��'[8��bS�r�^!�|w�a�`��$vH
rUib ��.�i���Z�����Ov�u4����_�*��˿����@.5�1Y������^�XXD�����G��q���=Xe����+��:�h8�%�E&�;V�ݦۂ��ݤ��u)�Î ���6]ٷ��4�UC/�����v�ЈӘ����`0%�h����^yy�i�����;�;��-۪{.%Ԏ��nɿ簏0��������jp���ê�CL���/]�^u�߈��1q���ɢธ�Ą�{�I��h�Zu$�D� ��IQ*V�x�G���B�(/�_���)脺���FQ�_g�k�n��6w��f� (��@��	O��N[��̉�C�dq��Ƞ��n��]�1��h��	 ���������-K]�``�7�KW?K�P�o��5��b`(�8��vEC�G\K��>p�c��"�v�+l){m�R�Z7��
O�o�[�Z'Ҹ�����+`'�-�Υ�$�̠n������WЄ�!�#lK��aP��"Š�>"3p��\�x��6�7�bi���Ym���OJAX�I�$�v� j��qPF[�b���I�#x��tn�vg>o��@E����f,�0P���-d�`�2�R�@J������F׌6Q��]����[$�AOe*q��1;�������.K��q�<����;�r�5:k�諛��җ������͞hWT6"MtT��D��*N!�XBl����"�ȼI�����}n�u)�jS�,W���~>��)eƳ#4k֕�Ж����U��;��ۏ���t±�
���-M�S67�Dl��ٽ�y�����bq���e�g��2�AC1$�	juƈ��v��ə�Չ��USՉ�)<�f�pOb�
2�j�_��EQQe`�a8�6)�z�h� �i��u��!EY�#����oա���K6q�jl���#��-��q�p�%�Ӽq����R���"
2�\��!�:�����x��{ ��]��c�_ﺹY�'��U.9W���U�LQ�ib̄�!�Oy��m������`Z�C=9u�8�kxp�|:{���u�ATw���2��&��Sl��ۻ��uQ����W���?�]s\=���nӹ�0s8�K�*�������|6��*�+��SL��#��/�A�#��)���$	����5��]�H}�}n/��<�f����p���>Y��!@C�Έ*ȜL�W�RD�ěkʟ��/�0M�R�~`�w;�x���S�E2J�ɳ��+2�B/��ֲ�ޙ�$=�du�����Zl����Df������&�F���7M�>p$"^��_�����p�ڃ�N:"�PnoTk��Y�l����k*^��ݭ�)1�F�<qH���.�#�R��뾬(1�o��X�$?�Em�=jF-4r-,�'(����y��q� 0�;�gG�Jț\?
���� rSC��,����"�me�e>C����M׵W/�~Ye�
�@��3�2 �?�xTMƸ��[+Jf$U_,���%Ms�{"^�]X��>럻�>�jy��ň�����
�[��w��M�h�L(�%���?穌�׊�!�3�J��a������s�u��O����s�\}db�׎[HJ���p��	\D�������4�D�@��!	neX�,ٸv���%ŕ V�� �^f�+�� ��@��|M� P �1/I�Mcѓ��0>�^����SS���Ї8�(�y)S"�U��5;��UthǠh�F��"6k���:����&#��ɚ	k��b@nV�)��nD�t���/!/�fBA"Đ�Lv$����_��_?Me+��m���,O��@�m�+��N`�h���+PJ���jq����o�Бa�n�7~k}P֯E5�Wd�p"�Qr!�&���`w�z
uZf�"�m�T�l�e�|��	e�7piȗ����հq����頸H�I�"�5�ճ.z;m����`�!��.H��q˸��S_h���E�*;Jz5h�r�>ɫ���vU�r�C�C&�����Hʝ� ��#�ymԔ�G������M-��S��P1C�:3F;�r/"2����Gl�/�B�S%������Q�&����r��!*�0�O��Z����^�=���CO;ef�x�8,��=)�����׋�D��0����^	���w=}�1��fj�+��|���C��7���M�ވ��r� 昬��������,!]�[&�A��v�?��� T��pA-���h0�!C8�Ӵ�?��8?�#�g�~�`�I$���AϽ���jK���հї���i�Mz_;���W��`mR�³elBP�NwȦv��_S�
�Z�Ԫ�e��0q�*e��T���"�_�%�>ɟt�)��P%�JW�"P\��ךT� *����?��\c�Q�Ί���>`Ǔ$���&����&'}A���@&#�!��c�!�[���d�����Wj��X��Uȵ
�����-s����wM.F�8�~��ժ�i���[ 6s�p'm��>��綽	^o�N�!*�N�㦠�C%�J��֬� ?�Yo�%#n�ONf��$��x����L'I�b���-�?�z�-C ��������wAk:w�O
��]B��#Y\M��3�����JUd�~A�ۍ�9JAx��vX��8�"L��"���w%+��v\&&Q2)�Es��:ѽ��#q�ڒ� �h��e���nYtP�G�b�*�����5.�81;��!�pűh4 ��Gի���^�V���LiE����WM��b���*�_ z����vMj�N�|��@�����Md���*H��P�� �?��VD_,|�����i���!>CBf�/EO���u����+z�i��"�d����%������6uG�ޤŢ�]�#f�E�Ůݏ�#	�.��8%f8z��d)��mm�Bn�����)���8t$��w���Xt>���Iw�|�ZO�����:���E�h�������I��6ܓ])�;��"��-��lb��ei wS��Z����hCUhV� m	��~��G��:s��'�� 6WJ�z�Ui���~�{_���P�Ap�5�d
n��_��4P�ÅrLɮ#[���єڻ� D�����f��+�w�����܎4�b�,�8�mĴ<g��9s�0�G2%�n����[��P5b�L�V����O$&�����T%t�<���6-𧤜4����!�#F.2	����U1��yx�l��as��\������?���'adʽ�A��Fb�HP�/��:��{I� �zńU�?u�cCb "L�D�N��<�BT�p�d��b]���P��U��`�!Mi�P6��&����z0<���W^hi�P�<�������T��	q��<����(xaGZ�EL�Y�v��7	^a��"H��4垚%��f i9-c[��)���q�B�X�8�2%��^��%do��*b�W���n�S�H�'��i<·޾�:P���n�azV���'w�g~Pk�$>��)b�-C��@�4=? ���3x}���
�x�%)R4�:>,O�]�\`�1<'�����.*@���Y�]�k��Ħ<vj�;a��б�U���..c�Ba�젆�:8ހ����z�oW��k�*��OX�f�|���D&�tV���@��u;�	�^s7d5� �M�m/��g=,�*�ݶ^3��ͱ��vV� */�aT�wX��"I��w����L`��Uk�LY�@�VqtOB1oz_�谥Kx�"Z�%0�hͳ �LY�����gTnp��� �EǍ̼�BV�?�Ki8�N�)9���yBٵ���]����������5񮆥���4}7$*��/9WeR_���p�.�mT�]���/�q}>��8�'����ūy���s���L���P�[I��jm)�q�l��{0�����R�n��V1�O��*p�$XX�I�d�?j��|܁�]C�E��t�=-}�*��B��LP)q���C���k��4]���8&q��?��`؆[�;S���y_��[p�F�ŧ�w%耴�@lN�61�=ʃ����+w��G�����yN��b�"~�?���	 ��Vi���'�T$������������"�EO�h ǭ���B.fr�Q���ƀo��5�*�P����o�-�t�O�*��sC�@��Tc�cV
�6E:I��DȽ���`��d��	0�;����>APQ�ViB �~?�p�+X%9�b�u_�8d�!���r[�������ce6��{���Z����ߡ*�q���<������_��N��Dl��l���y~i�� "Ns���������K�Ngajt�"]��rILb���u���ԓ�5/��׉�ߵiؓ��.��:Eo�3�M�y�����l�j��\Չ��;��B�M����4��l��%51���n3���e�Aޒ֖!��?�+���7ۂ@��|�7�H�q'8k��W��>E��P%ʽ���U��M��|L\��0վj˪-�}G��r� ;��G��`+v�f\IKUMj*h�KkD�=3Z��A{.O�W
\7t��K��5#�-�'�4\"�'��Y���GQ�Щ�\�r���������K�5AV�c�,�:�aj8��p�i��s��}1Z��=��f^���M�tG�Ze�k�q�����6Ӷ|p�ɪ���S��G���.��������r�  �dFQ9%\�GD�~62�w��w��7O��R���l�]+��tg�!uS���/���_Q��6�v�ā-p�$�O�����k?`����.���E��s��E��Z��8��JFK�B������n�-su����p����ӂ��MX�M��^����Ϲ��6��қHd��S�u<�1�eB��U�
�k�3j��SZl���/�W�p|<o Su���~���+�>�.fe�V��߸GC�	zh�����U��S���&�.3��L���Ł�i��6��>;���ܑf���D��>ڱ�'j8ߕ*N�0���$ASIlU�����ܾv�p{th�/Ϯ�W��{�%vN�*=ڏ[l/�1��`nQ}�ݡ{6֝�M�Y���0R�;cǉ	����]�2�JHbČ����7n��g���[���������R"�j��1��|��+8r���u���Vo�l��22;���2yފߘ�9�)�K��Io^���[�F�6GR�fnP9Nw����ba�T<F�|�N%��
�C�Fв��f�'oŅ�Z~fm��} ��X`_� ��5J��"����˖�-��(��`����׎Y$�@=���ׯ)�"��D��7��ϗ�!Sz�����Eu�	4�!d{��2�����Zӫ��f �t��z��:���H��'��>N�{�����3ߞ�����Ka_����l�x����L�����~J�@�L4�0��U*~C3`��"��ӮrF[����	8���S�X���H�ҫQ�
A��&����dJ^��"��.�;v���17�g }*�{��BWԏ����(f]q���H!�Ð�7�#(4ں�Ü���i�g��G�S�����Y��y8�t����w!�>!�`�����}��]Ҏ��a!-��J���\l;�P`>۝R��Rö�sa.F�J9a��H���L�;�?��8�ՐL4�?/�Jb��I{�����[�WF���V�����������C��ҫ�;��3.�q\P�D)<�ްܑ]OM4�r�/d�g�#����S�B�ۖ��>��n���0��`����}�A�a��p��u	��2H�i"*!�/:t�[�4.�V![���f[�{�U��g�����@�G�����N�t'"!08v�*�
�C��sy�vY����Z|�v���UA���N�kl<|��gc�?��%\TLI���Z����;�e���}!���b��-���|�M����)���i0��e��H�7J��IѪ�pf'/pfn���r�/�w�[ȩ�ꃞ�J� TNbi�f�p���/v$�3,E�'S�9��d��nG��8���/�z�7\)a�)|��Ő�W����;�Bq��!�-"��?��RVhx�t���vB��Q�_E��*�:�"J�����o�&f)C������p���e�H����.�#�5$Vs[�f��)��_h���}�?b��Z���Z+�-V�IT���4[�:25�e9x/�`Q�yI�/5`��V�ϥ�ѷw7e&{���X�nklR�� �Ό�T�����T�`��: