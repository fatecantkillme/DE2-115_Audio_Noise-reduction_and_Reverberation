��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|̪��q[�d�v�?�X$���C�O���s�#��\献l��ȸHm!�R�����<gʊ�O�W�}#�4I�����:�u�5���`���1)���V���͜]w���B��<�+S֮AN�G��J�8O�ER�����ɾ��gt�����z�,�<�X����S+4��y�S��<����|�$��ޘM�r���a�^C�2��|�=|/�>��@��ݴlzI�j��;,�7���� �[�ޟ�"��V���Q���cP�� ��$i�$�ND�*���� �QWډ��59-�rA�q���0��L��/%���4q��̷�?�3�:L����_ �0t�Mԙ�%��7���jbT>zT��Ώ �+T<��-Sϰ0y�d�j�����y,�V��Ⱦj�����Rc	�4jע�+Y hb�t%��/���j��^O��������G*)[\�aH�� R�jݣݔ�a��H\\����L-�C��ĢA�/4F&�4A����Z�!��{?���^��f��ŕX�qƪ�'����C^����E�]T��Dϓ'�,�U^��+#T�~㏉W0��6��ǂE�j��j+��]Z�p��������M�1�F���kp-�˶1�]���?Y>�F/E��?�����̑+G%Lq�Ҽ�ߨ����in�'9B��A̚n���Iv�x���6֌WPo��::%h��O�_z��D�	c�3�G�FD!0̼�!X�WX#�ɤ[Xr�i��kY����'����w;�Y����}��J\Hڭ#1VsZ��u��bp���ګ9I�e�d���c�u/�" J�h�ť��m�b{x�K��r�;j�`nXӕ��A�+(RW0�D��M��]�)(�H���E0ۡhk��>dګ-[R���5a�Q��uy���B�#�B��B�x�r��cy*[L��`p��"v.��Wj֎Ҽ�}䀡��2��_W{ �^�#����ikVɭ�����D�r�y������*�����p@���� �1'�L�ȅ����^�g��__]��%�פ&q�C��]+��&�I�����w���Gs�5J95Iㅥ����v��VQ˞�?mSCY<�X�4$`yt���'���V�R��(d4~�շj+���3w4��1��V�Őm˖	]�*��!�;�׏�s934�C�I�oɇ�v (L� ]#����#1��D0Nͥ ���v�c�r�6}h�.d�aꞹ��>X��2K3m��|�᣼�lVr��}�~������
����O&Xo�la+�
�ǳX~U��ܜ(����z�3˄��Cٵ��sۣ!Z�&T��.s}tAS"�gN���䦶�Xň��吱�N8h��{Mj��Q�k6JZ���1 u�$4��Ť�w�՞�u�Ml
̻T�5�e*�6�4A߉E��ψ=����*q�H�� �K�'��#4X��U�����1�93��L��[�7�R�cQ�r�p�@(irˎv��;�t*G����n-�F�c�o��u���bH�n���B���q��z꠻���,����6��6w��2<���s{�',�-Ĩ�c��a(�ü38�<���u�<,b;]@�Ay@�����:#G�/#�C/��anݍ�T�@ ހ��\2�t�� p��3��=ke��NԤ�Q�_�V==a/NK;�ꞷ��u<����dP�F3����E0��1��&LV�*Y#���K�?��_� K ��4�@����(s�r|kUX��f4¶Èd١bv�
��H��z`(b��P`�p�V��`�3KƘ��+O��>;}���G���֩�
V8Vҡ_��դ�3q�<�%�&��_�'��y�y`jU��5��z%������$����f���-y����7 (;2�u0�5e���}YgC�y�3Y}����fM9tj�ԃ�,�-�X�Nh�b�(C�=��LOY��H:WA���'�W��s������ĮA(}�H'�����_�b�yq�΍
�����mY��P����<N:���WC��Wd���6r������H�����C�Q������Մw��s����[}���lsݮ�L�0{.�-���LЭ�`��Udz�"�!`�ۮ83+wj��∪��ע�
` �%g��[鶬��"~���W�I�/7Y!Z��u�S>��J�J��F`�:g���^��E[R_K/�7n�����r�B�I3[�u0A�3_��m��� O� �J�K�n�����{3L�~w�ú׍q�R�о��DZ<\������4p�=3��y��dk�J�E���%|8��w��3��Ӵ-V�6z~@1ӏ�~��BA�Űm��82^�I�a��FW#)x���zy�@�7"$�l���y�G���m�g!� s�����-x�-svb�~�����N�@uJ^�@��m�_���կw�O�_k�-�h+6������vڈ�v�!;�H	5i�xKp՘ݸ�ů����f��pT:%����LO恵o=�4�F�GkLۆ.	�ڈ�(�,�{�9�Q���o�9�1ktHfY�C�_���A�/Q�xJ�L�B$���j]1	�џ(��X�y]�.PC�O�m�?�$��A<��2��3��I��p^�E[P .ۿ��9Jҏf1+�����f�*��+,�mU�r���ZD�L_ ��`��K�����e�`�D���0pI��Q܏���.ps*���܀~����$
���[���g����N(��A����SJ���ȘP�7��^��.G�	���U�faT�1�	N\w� <ǥz�Pҍ3��x����8�J+�)�qF�`�S�4$��<�nP'���	i�X���x�=`
�q&�sBzSB��@�(��N.ag�x)f��ƽ�t
��ɇ�f�*2�+�J}��@`�
��m���|��t0!<��s.B�7/�q�*��3iB���Y��MUR[�!�'�T+�
ڹߩp��%�x�x�.�׃{H:���m	1��z���گ��a�����M����v���,�A3gf-!L8���c�c�BǷJ[������p�#���'f'.�E��݂�G��A�Ow+kz7���v ���;�ؘ���뾭V��H�Q嶢H�P?r�����!HA�h3d�2�BH��/�/�5�H�VK��,��g�$�{�����_�~MS�&�0�I�"����'H�:�����%�A|�����
A��N`oƸ{B�r������jgo�(�`Be:Τͳ�&������{p���C)7�Jv$Jxɼj8�F�'����L��=D6��|;��W#Ș	�[�����qK{���1sۚ����ұ�*�4�͠��g�`���S�ňq�&��?�o`],�/��H�g���V��Qlsd�s[_���hB��F'��J�B3�!�yb�R8�nc�]ڨ��6]Z}<U��Z��"�\M�+Ndl\�h<�p�����#�A��K�{�Ș5�Tg����Er�>( k�}i�*}�W����h)�Q�a 3�!k�u�o`3כW����
�@��u�o݇��`�dyMwG�I���O+_N�
���ɽ�����ӭls�'NB���O0?�mt*�H���z 3J%շE|���-1G�͉�3�����]N��;j��,�05���f��$W#��s{S�.��u�F��v'��L�����PG��Dl��\1b�h�O{T���t�{q�� V�DVM�Y�Gz�sQ�4<p���x]W��W�+�v��Ё�4���A��	��Z���}��[Q;�(Ր ����\P�;�����bf4�3A��<�.��Um ��[�2c��Π}eЎ���I��86���@K�@���em�}�gx�\���'Ϫ�s��������3���¹��f&�J�Mr�˞r�zE�ct�����Ż[�'�]i�ƴ�MAF�-Fxc��h������چ7��jF�kM���+T3=��ae*�袎��4����4���'�X�?HwH&D�:�Q�y�ܢ'�Z��{$�[��'�2(�ݵ��`0��H���u�mh������cI�ᤔM��4q{$���V�AL���!�7K@�LO�<I�������xu���Y��|\�a��"^�kD,�����XE~��4�(�tI�~���I�Jw�v�����D=k�J�Z��2&9ӧq+����7��'�n���&�15/-3��N�b[��LHf�%J��2��ǀ�7���� �nL�;>��l�lo�^��G./��xkL����w�c�_�M"�څ�ǀn�"�e��J��䐽���⬞�����S+�>9��2�B�zw_W��B+��.����䄶,5��p�>ko�u)r��,�lb��M�L��F"�7�h�D�B����dQH:c:P+�xx�,�K�.����/��78؛hrc��+	jF��ZE~u+maF2 ���=�1�Qd.]��u�R�jiB��q�E�rA�e%OȢ�-��Z�
D�.�Q�7�c_�'X|�~;�`�G��YH}����v#���Ӝ��i�.����׶8i���<$�<����z�~��Hڀ{�vƅ�Ė�W�$k���<�@[���ò$��1+�j���w�=�H_��7ZK���Ù`��_7�:��{!�0�Ս�p�
�^UT4zY�����J����
K����t��m�c�燮���M-pŪ������+�:#G{�0��-���|���ʤU�`~9 +���M~����i�������'��@�M�2���ڤ������/�G�(���g%zw@L�Pܫ���!`�'8��ƚ�6h�p�� d��S�<"��A:��L��NP�ćs�ia�-�� �3cBR}��y�z�I*��ZP�/rI�R��D��˭��AT;�ht
Ϸh�X�w�E��P���O3�r� ߧV�b�U��B�g'������­����F�RQ��(��!��F�_�(���2+E�7�k�K^tENp�"`��"�b��r�ʗ��s�G)D�2>ޅ-�[`����'ޖ`�������l�Є�Lk��u�+"M2;��lR�邂��p��
�$(M]�W�B� ���;�Ou5�K���+�Խ����[�?|���He�� ����µ��=weԐF1����^gs��[R��ˋ�'������t�ɑ9%� !U�nEK[�l���O�q#�qT��Vl��>��7�e=�&fE49�p_���Hn���8��<A4y~@=0o �ew��_�ހzh�$����kp��#ę�����<3�Q�0��:"w(�KF+�&S�9�&ٓ���/