��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<�y'�I�zc�2����@ū���6k��E#���ۓ��V�}UI�q�h��7��|�����]�^�[�n��s�Gpm���Dh"}�����p�53N�V����!#`�����C2�N�E��Z_�a��D������ةƇ��{�M-����_����?o�krx���Rt�Kj��֏�����4��2R�i�B��O�ZM��V=�Ҩ;�e��S� x���ʪ��ľR����"I	%��	d�5�Z\D�
�r7ϦP좡�O���*�M�W*}�W�-c��$��Q ��h;�e�+tT��'Ǫd��J�`v��%����\u�*Ր�/��>�����Ӗ)����cS�f�h�ߠ���C�kjJx�.�P��8z<�@��~�@�u|戳�bƝ3��W�4Z���ѱc��y��y�A�^�#.˳�)�[ ��lz6��4�$�f�U���y�L	�Q��r*&����6�2��GaH|�霾l���:���X�ݯ�͝G��3�"������s+x�DBUy�=�������eZ\{�:���9��-I3H
-�_��=]p�)pM�QK�ɪ|�AeGh�VHc�Hj[{���"�ʡ�|�*O8��xp�W!�p'g�Z;kf��6�|�}��떩�<�(�6\Ҕ���\�*�P�wWL��#^�9�� 	�q�
~�v�jiU����y���=�y3���6")7����@(���JO�N�ŝm��%�>��Y�A/��}��@���ۑ��¦2t�����4Ty�.�++� �"�1
bD�_��W;�b��]�9��,�����*�I;N�;ug&:8N����0[~���^?5b�z=�ϛ���>������Iɋ� N�}�#�^�:�pwo�ԁ��p���m�_�|�/��Sr��?�oõ��[{0�8����N	[�E�ϛlm�_	�D5{�?W�P���x|[e֔4���>�ڇ�����f��$�߾-�5�O��=�l���0��K	���@[(X�N�۲�_ɖ�=r:M��}���Mi~�-tJ�Q�Ld&�Z"�{
_�^_vE4�b��έAuĥ�u�W��=8�qz�����E؁A�$���ſ̄K�W�^N��\3��;Q?"J�Űz5K�m�U��E�詷ϐ_	�0�\�ß��Z%Hߑ�ϰ.ܑ) �t`�xaj��e�h��ΐ��'�͞.yz�5|���Im=j�֛ ^�?�Ҕ/vaj���A]���7̟ψ���:�7����8�Qg)1a����{I��'5�BOs�;��i�5qn�'��UOͼsԎ���.mO�]�R��oU$�\>^��m�µ�G���Q���Lĕ8~x�`����p �$L��Q����%3$�(w ���a�Y�h�j)/eŢ��o�eb�����"3��l���47>�s9s)�V�5\��T�G�1=TC�-F�z��Or�Sr��<C�rF���p5��ZW�G��"G� �Z𪷁g�C��*�Âs���2*���?�U��dH��^�����e� J;dxW'^�HCɗT�0���?��4U�2�P�t;������̍���>�I6�T�V�r�D��	KF�C�����\�܈�gv�Ůʘ��O0��� Ve!����~$΃�٧͒�"����J�r_�O��V�Bҥ�{�L����N[m��aʿVa	����3�nJ��{(�LUh�6�#?�7�o��%�V���h�>�tirl��n:m�eE���A2��>�cK߯��������7������0ϾD1Q/�&�F�3��Ϭ�2���J����ǧ����i�G��Ƀ5;T�Fh2���}Դ3�̞���Ĩ �]w�e�b5�C0 ;�XK�+�P|�C�e}�n�Ah1+Z���#EX��i��7$<�8��
���T�h��Zŧ�8�+�t3}N�bQBeS�|\�zc��a��k�y���9�_F^3�Oo���W�����U�e����x�_|`,�3gx!���C�1ap
�f���;�قbdmV��ȓǷ�Ib�>	8�I}Yg�+��s?7ʻg�BUs+���(:K�@�=�>y�VH�|9�iX{�O!4��)�ݢeZZ��`+|���.;û@[��I��Td�y�a�o�c��|#�r���iT#���!@��'2ne�GMu �!e��nAhԝ��V�x��� �3}Y8�A8 �s�8Wx&��o�
uL9gk��vXc�d�=� B:s�_)S���6r5ྉ�����t�YF-G:y�qx�US���c>��թO��*L��*� ظ^g�E�х&�,���~#M,�.�ak.��)wU�������_�JBsZY�|��:��,��6~ ܴ㚬ދt<�J�s��RI�]�������EM��[�7{�����=���uH�5�g"����>*8���u��LW�f
��C��x�$��hz��W��g�Sn�x�B徵r %�-dG1�zf�,�(B�N�=��eF9Z�-��6�0�a���QZӂE��^���Q����q5�)������d�۪��� q�y֩�DcG���Y����E��pŉ��	),A��'��K��n/��][�}	� ��n�$�Z�u^B���~�����:� %���#�O.S�LŎv�{�s�b�G?���1�$o��t".�:~��i� W�Gr�Kbϧ�'ׅ�k��v�,�ѕ�k�v��I����QBi��B`+�ٖ5��΁n�D�E�Q�l�=�����j�B��E)8�y�z$��mC\�1��$����MV�N.�Z�>���v� DLԗ9�*���MkK�7t0uc�|�W`��KJ@�| 	�c��0wH5�Gb��	O)��a��?���y�p�{�,���+i-��YM4Fb��s&�|��Zcߗ��C]h�I4zD�8sy�:�ȯ�06m	h
���?՜eA��8�d5����-LV�+UA#i�|�q���w��fZe+P���h�/_��w;`d?���a9P9�!aY�6��-�#aչ�6�� ��<w�z9��IrT�Z�µ:�Z�Z(NkK�i���^��A�#�oh'��nW��!��W��W��i#�k�f��у��۞*P�󪒔CH���ʺ��!z�׀�z�o�}1T$e��D_����K���g�F�8����Qo��a�E�-�B\ ��5lmN����>o"9��7.�T*�,e� �,�U����'˺:4����IB�i���n��}ebе�2W��y��Sמ�����&y
أ��|:���@�x?=���i�� ��n�n�fO�Z��+�V���{�m��!`y��W4�G/;��<��%�=��Rx�DZ�5�R�V?�>ܙʹ� ̜���d�P̊����Q�Wpsբ!a˄��m��J+ka%��ô_#x�3����5��-Y:�&�*L�}��� �� ��K|a(�?$�U����(&���{�5!fL�.�_��!e��%��pk2a�]��o���X�N�������C��Gt�I)ӻ�6DĢ2^4�[]�>��r��yj�#��@��2���\w�=���: �(t��U��sE���2�_��?����PT��	\n8k͢˵�6GO@ᰭ��c�_K]�^,��0+�_�%���8f�z���C���U"(�%�N��j�52δ9P��Z��Kf�t����sye�o����6{򋈴�p��"�$fm��:��a4�b5��K���M�{���y'�Y��W�O�%۰B��h�ٌ�nX$B����&s_�Prc�:E�]��{b��q��w�� �:�����F��"랲�%-L�"-e��(:�<��1S�)�� ��j<�P�t��=Ǵ�<��ahJ��q a[뾥Ѹ�q�|�$
����2p&&(F��N3��y���<%-�`c>�H�F�b>��u)��6���L"��nG��M����)�"NS�����j���4ޭA=�����,γ��@5���EQ����p[���ڡ<��06\,XN������7ˬ!겝���E	Ŭ�W�5���v�����H�Ls�L�[��U��.�M�f]�z>C�FWw������A��;L��6z#�������+oɅ舻4��J�WtC���Pl���>Hwa̹H\���f����L�P�{�� v�F�4���8�C��;��Wy�,H�E�Cw�X�K���"9-�t𮩼ƴ|F����*�	JpRf?��D�e�ml�c'߁�� {��v��VJ١�T��,��:�<�̽��aA>���ݍu���A��0����8��ζ9%r�y�'ݕ4z�#G�fBy�Hi:�U�]�C*���n��W)F�WlĜ����Ù��9�X���������{k�H˗��h+W̋�E`��)��ƷZcD�	�_�?��Dyd4]H��NGԢ�ᾈ��m��S�w/+�Aכ�@�T�Wwn뗶���i�t��d�#�*ͣ*
��{�:]�I��'> ��$<!��[O�|`�G�|�y6�n��I+Ě������?*��m�~��\d:��-�\�T��'�6��'(e�<�����Fc��39,��i���.�/����7����z�`��ȥ��^������μUsÊ���l(���+XW��T�A!�3��U�<"6�~r���;6�G9cUlV�҄p��G���`|�٠��
�v��@�Ap75�M�
̡���cQ��Q����o+�2�����N����?�(a��woD�z+�1a���OF]�%kړx�G��/VN~=�ЦցV�>hO��K�G���_���/^��2�3	��HN˕Ȍ��$75��h�%�Ȍ)&����+�dP���%Q�<P�T��:w�&$<�Z�kr��e`A��?�R
.���^(p�;�	�S�b�h�y�ӂ=#�j�cB�.�Љ�h���t�y�^k���Op��Rf-L���D�m.:\�L����8 O��g8e���*� �)���fԐ��$�.9ހ���$>�����=�ml&����'�18��i��>��ZaBh3������^iMU\���p��r�le��w��M��j����-6P�U��������L<$
_�찰#%��P�Y�&;��X����&�����4d�l�;4�<��������%eX[ӡ�*��Y���܏Ũ����Xj�i˟@��o��Vc�W�넖P��A'�,�z2�E��i䦝^�k�Z*�2F�2�O٥��Im:Ut���+�JO�r�ȥ{'�cu��h��X������'O�a�e�s�T����`�R�T:�q��!Ё�O�;k�Jk�_�
��f��a ���w�*�ԟ���������č�N�,�Yq��ٟ~�*���9���'����^!����Yr���NR�B/���jT\L��A�<��Y��ۍR��d��s�e��D;"݀���*N�p�Qp�dƮ�����Mwa$���@� �������6W"��K��Q�����ɯ�"�����i#I��T���V�I_9�������͛�fs����ފ�v�p��g"#��2�6����J=�o�ָݳr��>�l��q�@Y.5�o�w�%m�>^��Vi����k%�*!�9:�p�T`�|ѥ�iq5��so&A�:��F���hY���ǝ��^A8��N& ��%M�?�F�[u�!��S��R'`qVY�>�25��eCR
�έW(�����u �eq�f�5����]���M�S�2���Zԛ���<�����`���l%_��	���S*�xq�������O�a|	 �ͬ�3�-�1�Q�@M'��}��L�ID��$m^�ۡ�����R��S{ԇ]N�,�ku���/f0�U�šoD!覬�c5��*2_ |��
�_o�m�i`�Q��-��*�-��0�L�֒!*�LY��0f���|��9T[�>��ΤS�ʥڤ�R��h�׸��Y�QNǋpܮ��֔��}���[�9�������>Fz0�u�92��`by�%����jt��ȁ��%=TՕE���N��Bu�O�n1>2�HW/.���ʐ};�z�֯�l����OO�����Qſ�\9�ow����qp�j:��,UnH�+wf[�ʯ�z�U����s=Z�Dԅm�$�aZ��I��faV�[Ƶ���LE�9�C��1��!�ώ�_X�,���̩\�}����Ai�<k��f�SW7�i��b׺O�����mB���A�3�'�y���2�*�~�eN�j� 54M�B���
s�qԻ�����5K<G�� b˲_�J��/>8/���r2|d^m9B�Iל�$aP|�.�������/79�Vt(q���6�:�w�$�K�|r��=�Ș�ei��1{&,�j�.�4c���,#J?-xb�/J��!*�[K���6�; �e+(�1#{���]&�tF=3�̪�����~c4�7x�J��<9�{�媳�T�V�q4C�@d؏1���=�����9��ml��>3�	��=�����{�#�wBhz�{H����G���!	S�8�]4.ԙ����<��q?(���Q�็gFΕ%2�����ϓt���Mr9 ��S�T�_��ɫ�0���)��(�Q�˾%�s�SY�Yn�˘�	(^&C-O�cEPK�[[�-A\�K0�t�X=�a�J�E4dA�&fI4[pK(F��ΦJ,��v�f����'y�c�p�nCY�Gr����֐.��ȷjr�W+�˅.�p��*��/�+�*�D�	�g���%�:��2�����
	o�a(�h��m��X��ӊ��nfP��H?�����w���zG&ν8�zX&�J���EL�v�1G�I���i\Q,#��+��H��O���<U峃-����; �� �M�9��ς>�;�#zM���,>g&L����sUM��P+���3��]˘�BfqX�sg��^.C�Z���B|����{�YtH�`��Id�8���Qǵ.��
�a-�,1�?�l�g#��;�b�%wc'��ɛ,��ֵ��n�-�v&گbA��G/������az��-���4�x^�ޚU�V�F �F�7p�Wd�"��Z�y�yا0�mY�EOM
m8H��o��Si�����mc�����"�;a�:�ddܙ:s���E������{R��լ�~�����O#81zS�/ጞ6�@����Z��l"�T��8�����n4�Q1>̋UZ-�!� %��SPB�e9����6)C����]υ�-���$S��d�.�)�u��eI�����Eh����i�b�#�Mt�K�-��`vכͣ3,��w5%��<=�qץ_���P��B/�� ^�+���xR�:�?HN�%��~�����i�=�PҹNZ!����0�d!v�N���԰���i��@��j�Z|���"z��(GPxσ)\Ҹ+?�W+�����!2����s��|����PPyl��o�
�0V-aC��Ub��u�VST�~���6�k�@�T�gg�� 4����a�M&�������+z���LI��u��M�+UPK�`wpX뫊8�G���T�9�3�Z�A�\�͐�X�f��~�Z��a,���1fo$��8��?�K�Gt�q4"����>��,��r7EY�m�`�0x� �VI�#��2�z�0Y(�ߐ�6dd)�^� ���c��@�ӭ��ϓ�I �������`��Ҳ|�؜m[�
��ldeϲ#��~_!��@�(�?��6�����Ɏa�ߑ�WP+�Pc0Ŋ��e!�5ӥx'�Z`�#�J��}�:���A�
 |��S.7���#`:@����_��H~�[�숫��hv����Qmz��֘�[�j\բ�����2~{�{W���=w�a��4����,�߳AI��5���`2��*h�xb��pG3%�~û��װ�����~���7�M�|;��� �s�k/�7q�5l.�ś`Z[Y�,E����{2����^�8@��u�e�ܕ�8;sH�a��)�Y�İb�U}���o����و���m���8^~BE<n�w��{L^�)�^���;�ZEn��F�LH\;��*!R��8!�.�_���f[��V�!����Tq�,��B�c���#�sh1���{o�<_؃����O-�� �8=,f��j�4�96�XvY0�W$�w�¡`P�t�l:����+�h��6S�%n�I0�-饕�U��