��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>,M�Kߤ��S��#f;�E&�o��X-��MQ���a�1�̧�^�"��0GO����IS�#8Q���+�%��i�︡���1�ڞ�<}g?�֨����1p�u?�%��ؼX}B@��{)�z���Az;S0r�V6��^)�Gbs r�z�E���ft�$&<�A�ƍ�7 T3� 5TX˦�'#�j�1Cþ�����{1^��}�D�_2�$�8Mg�x��O�S)�J2tDf�#��L?$�ǫ.�0��G�)�3��T�?Zc�H~� (>�T�Bqe�5��8�w-~�T��3M��/�U.G�iR�I��Bx�H�h;[�4�?�Ǆ|�s�
���39�=�$��`W8~���U�w<��w���p�ʗs�֕8J���ⲵ���w2�el߿GƵ^C�ki�j�/���I���is�Ͻ�\\_rF)�j2̳�ܯmQʢ.��:x�UzW�:И8����	mEW�k���mHeI�Ux]c�5\!~�$�����ݶ!=`�X^����z����Z�n�3_�o��b}�ۊ�ҍ������^[�f�p�N���*�S�%y�F�rQM�?v���� ��0��ɰ^�OQ �VbǢ�wj��S���y�C�1C�R���RUd��,g����oH��`��e��6V�����|B�R��E���e0^7Fc&LT�2�)4^���|s�D%�C�@u�߯�f�����������RDb�K��F�T|���l+�87t��/��M��SA�(K)�B�q�m���"�(z��7��nZ����5;_�Y"�Os�=���e,��җN7Y����6'�����&�\���ɴ����`��p�I�
�(�]Y��Ԉ&4��/A���L�P�-\ �VZ�g`k��#�)��5xB.�F���P�_Y�z\�������3�`	��/��i��y2)Qa
��-����7l�f�b�	ؒL7�퀙*��������Y.YR�A���x Y0�
��ixmCk��0�^Ђ3���E�F(�5��)�s*��������gYr�f�5�"_�ԃs�{{��ټϚ��C���v�����Oq���0�^z����������<�n�7�{Oυ/��#�2��ʤ��<��|��և}�ܾ�W�� ��^���ӜM��(Q�ET}�؜�ƅ!7�}c�gpr.G�[���)��%�8��K�V���"�E��<����"8N�P�:P{�lw��O�ȹ4rd�|���+w̒UV�� ]��0�5��{C��ܯv=Sg3�ѓP*V��ho"݅���ܖF �6^�o�����
1۫���ke��G�ڈ�3U�T-�taw�Dz�	��P?�c�/zE�c��)7叭]ve����(6��fK�%�s#$Ȕ����J?��~���1�ݻi�g؄�����	�4����	�o虋S�pk�J��0�*�ܢ���Qi�<pQ�lW��M[b���yŠ�v�o�<����4�wL�p%>ž$���79$�ğh��+�`�.�.�Nŕ9��������g��h��w���c��o��/'p
�;��!=�ڐC���c!�퉨k"�S��T��s�;��1�̨��H]����r��1<F��ZS�)s���rE��NP�Dwx'�{0��!I4� P����xNQ�>���'�>�!93���$����新�+ ����SU�U���	���"zҬ�&�o���Z��-�rZ�t�<�����@9u����
1|��ʻg�p�;��E*�<p�ܵ����O���W����Ej�J����#T�w��g��=��j�u 1^�&���~�g\
��v�J"'Ȼv/�Rm%�p~�z�԰�f����Et$o�ױ-5m�x�~(�K8��[��ʭЀRoHprmw�Nt-N;����r�/�(�̓��R5�iw�0k��̐��0f�>�T̥h�0+,����b��J`6e
7�ƴ�����V#0,��9�i���JP7�����5���3�p'g��G�ȝ�N��,f��#K%�u�PK������ɛ�Gp�>l���Ȅ��͎E!��Ou��6LD���M�=V~�ʠK}�SѮ�X��N?��|1N�c�,>��a� 
;�[��<����W�F̸p�κ}\ݕ܋��l�a�����<4�M�ǈ��ݚJ��C��n,�M�"����0��e8h-���ʯ(��ńKl�ǐ�Ŝ���ú�����mB��z@!$���F/4Y�ǁ�;�hza_��*��0�Y� GS+]t�?[����4�4�L>\�~�o��o
�rl�J(����}F��~�3WC]��e�Z�,�Z&��N��8�C��|�pR��ߑZMbn����ecuzx������U�Ve��N�n��?nۀNVR����3�\����ڼ`��`Wt�v}���c��~�(w��[��sF)�K<����;�K��љ�ę%�~�0��@`�o�M}#�]в�3m���ܶL����W��h3(?�P��,ֹKQ�Qz�Mb.����h�<|[�B�:��,Z�17Uẜ/Nfe;fѦ7�u�uT��Cw�	�+�
;-a��X���=u����&{�<�� �*Zr�zIMlu\�83�%ŵ$�-�T�epN�%Hm��SvMnGs�BVI8!s$&t�t$��ۺӫ���t���ID9G\B2
L�F~76�SԦ��p�>��:���z�'�nج5�Ϙ�+ҡ˻�� ���):�{ܨ�
�tB����SH�KF�1f�8AI�ݨ.2��@��y#���+E����������ʚ�Uڜ~�<R$Ш<��A"X�������A�Y�W�U;�pQz�:ڬjl;��vd�!�?2� �-*9t+j��M�FK\�+ؑ7��jW����|�y����}�*��]L"Hd��p�+fGRc�Lk�y�#� ���8mr���8�q)Y[g`��+^q��;�y����lV�{�-��XR�%J���g�݀J�~$� ����5[��cg����W�ϝ�D�Jр\Z��)_徂AD����H�&{{ͣ����@]�;C�y��s|�W�p%d��E?����K'�ӝ���,�� �T�}�����7���S��-����������Ô|��Ȏ�&,�G�j����0[�pt3l䆱8�Jl��6S0H�s��1���}�,/�t�Ž�E*Z���R�>�w���q�P-!H19��A)�����ǋ�6��~I�.E�]��3��,,K	I��㽮��)�(t��f�P��]���΍�$����%q�[��[)�5,��96��c�ˍ'�i>�i��O�T��:$r���,�30z,.&y�3%��݄�ֱ@fa�-ʄ�ӏZ��쯬z�5	[鱺�P g�)
�Y��d�"����Ո_D�[wޙ�Y�����UIú8ɉt����+ޅ�>���_���k�/o�>`�k9����¡;���e�;������S-07��I!�(��ġY�\EIVs���q�W8gB�����(���ӱ#U�J�Lm/�?��c��=H�2,��f| ��![a��N�ك����X�/��Q@��ѕK�/|�CX[#tl�7:H��Yk���2�!�lA��-�:�ꍼ �[r��n��6�[�z.�ou��l���iDsJ����P� ]R��h]����1��JM!T�"W�i�i<���R�b�J��T��S>k�.;��j�@kVP��Tf�?ܕ����ZQ�e�j�����C�tx�X<�G���Ŭ�ZrCX��P��ӕs�t�+�M�_���Y�������G�)�v�f �Ql�G���c��哀�>��)����4���8�7	��c'o�|i̭���� |QAjFJf���*���@��G�_`-��V��s ʨ��w��rG�!��k[�,B�La����6�y��'���1�}���P6�l��攝���)���e%�Q_@��S)I1��(�	�X��njuύ�W#��u|�(�N'�T1���e�&P-Y]�:v��2�E�%���-��ٟ{1�NB{a���2#c%Qi��`�=?�e$a�Aۨs��fh�Fs��ܾ��u��#� ���+W$�s~�o(��:>��g��/�Q��_��d
��i����rZT����w{�Ɖ}�5F5�-8^iC�$�D�e���=�K�=��.��X;FoX���G�9Ǥ���i]�E �+���r`�}K��b=�F M6Xܘ�U���Y���	>�.AYJě�>��D�40"ƾ[Ww�%B����3ߦ)�����Ǹ�!kp{��j��εy4׿��H=��D�>\ڭ.0"����V7^|�^�V yگ�!ب}āu��9�����[�s��|���5�)�t-+��mJ��o���;3��LqF�cz/C��ہ$X��E?��	b�YV)i���b�/�R�bwCt��6�rc��$!�&d�==m�Pؑ������fƓf���
���&νV(��<������`���ǭ�B��q�� x��Ȧ�P����	�a�u��w{��lDAfU�>�K��"Igm�(���Q�|V��|̨� w�@�`#s���P�o�*����C�{4LUE��E����v~��lx-�wG3�>F=5���*���<�֞��c����
���h�;ϾV��x���{}֕��*C�:�YGr䓸��	t���`������akY��ۚ�9�V�d2�4�t�cnM���;�|zw4�(���jaOy��R�����S��gJJJ!cL�Rds`�B=�9倮��+���?Y�F��Ϧ��f���4�����ĻL��֌�a�<(B�����4&)�T؇W��X�2�I��UV1F�+,kT�y��ҕ����H��谩˷�	�:�i(T�/�ѽ��up�e�2��Z�gH~6��mU�O�g|�D���u�{ x~ؙ�Jͻυ&�Pp\�CVį	]��J���p��&EY�~rh���(���.C3F�qdk&G�9���ξK��Pӆ^�ǂԚ��\�0��1��Sb�4�m�e�����.�j�NR���C_��	����E]}u�;�ܒ�[�+2�������"hڔG�.�����׽hotqƜ/�̣�d_(���fc��#z��bO�663�� ,4�9��"p� \b���m/�1�]ot��Yf�&CĬe�Q�$�L�z6)�qTs�驜�"	{]�6N�k�ʌ�M�؈��Z7753�t0U ��p2��;�OB�/��$������)x��7�&z�`���27�ͮ����qߊEb%G)��U'���h��^��%�$�<>I�i}���Q��O�t������J4��E�u�`��1���f�n�����HM�93��J����D��}D�4��ԁ+Y�%�0k%6�*#r���M��MX���E��U����!ҷ�#o��:+�&m�cg9����?�$����@��G%�����)ϟ�e�P�-{>U�3���X�(���+ȍ���-��N�۠��/X� �i���GYtu@��+�Y����|�Ҽ-�De�ܐ� ؄��3�Єr�c�r`b��R J^�}#Fu71����z����V¹�22��&
ھ��K�E����8�H�r,��J-�=,��Y� n��Y@x�0�@$���#
��P�p`'Mۆ���e��`��α�����n����e���޹����B^��2P����.�B��v�p�[�a�-�o�I^����O��4ItŖjtYnc���e���?Y�M��p��v��'�+;���דy�IZ���i���`��%u ��	K/ѕ��*��5nt��"�ص;҄ eBc�:�����Yb���^B���w�A�`�"^&�y�3}��UA��c��gN>K����
W�w���J����+1 ]����a.���!ٵ���+e��p�쬙\۴d'�n��a�~�;&JQ��+"�&M��n_l)����<�g�_�v��9r� ���-�2�����n�E��| �f�-����İ%�$�N������_��Yڀ^ܥd�ʥ45�����X&��
�/�n���ҿ�J>�R�� ������
�+�w��+T��ls �<�[��6�"�3�tŁ��9T�	�(��(��?ǆ>��g�#W`��m!�hz�I�Z�]�9��j�hZqd��8��q>��Pq'C��?tN(���6蘙���zX<�dZ|������kLt[�.�%��AJie��7=��"#u_�?�@Ӧ@�O�啳aQʕ7|\PM�JϘf3@w@�-;Cf�j���U���$k�~��'� E.�������GF�%dL�Vn��\��R��k H�0��x$�+�_�7nV�=^IK�N �=n��zw����顛��T|=�X�`PEE��bW�EM�1�P�I�̶},~��sq�Z��Q.��� w��J��*��;I�K.�D�&���%LS�A� :b�ۣ��>�I͛2u�P�G�gŦɐ,��F��VL��&[�</���@�n���_�.=%��-�^)\�%�~7���rH�����Qu��Ǵ�V���l�箐��!i �V
Ӛ�P_���Y�ԓ �`OY���8վ��5�o�Yf��ǡ�S������|W�H�~e$;����h�|�c����r3-3��B^	��my���_��j5�$}w	3�έCe�vJ΀	�*޸y��$o�;����/����T|�QZ��au���φ�U�1���4�}��n�<?��A��/G֫��<CŹ�:�,���B����&`߈�Q��{a�������	޴�����Rw)��:k���!�,ox9�m���� ���JB::���=7[v�� �or���B8iG��O|�v���ENH��Rgm5h:����U���������pFG.�9�#IR�M��.fΩ�� ށdi�n� �+J)`�K�f�še�U(uq�T}��U�^>K��{]#�r��;#O�R�Du�g������>�i�le�0��zC�$�Ų0Ƨ
S�%E�p��=�k�0���*\3!�3�b���j�S3��.�y�l;����d�ȶM���m`a]��[6���|X�2��¹�S�J��Y���šKu��/�׮������٧mG�=��I�{n�^���	�z8ˠ�����s���n�#An�+���XJ`�i���pI<�;O'c��}��Sg�T~�t:]��T|�н>��=�t���1a?X���yr&y/sShґGL�15�M���"}��70�c���L��f��^���y,7g�x�6J
f�k�e�z���<yH(��L�Z��u�!3O-[KItfGek$�����"�	����3��&&�PɆ�u�A-ؓ�V��"�e׫� �GS:&3{>Kh�^�9��7z`� ��ȉ��f�O{�B$Pk6����]�FJ�^P���,7Ҧt���&�	m�q���������e����j�e�.r�X{YkE�7�Z����l�X����`;����W���M�E�%~t�ԓ���9r��[ C���+������7Q��<.��)�����G�]ƺF'>z���Ȁ���ڲ��^s��x"���מ�-��I'l:TA"�(K&��/��t����O�d��Hᠫ'�p���7�L�_�fPUET^��;q���.�$�/`��r�����^��e�ޱ�s��,�Pj�v���^d=r�<�,Pʏf=L�7��^�x��ӫ��A��D<Ld���p���aJ�Bs���9�I�V�Ώ
3�#�\�>֍L���$D�j�(>q	#cζ&I�\�+�J咪����z?AG�H�e�/B��L��k�vb�Xt^f((�,�2��
U����d(R+h�n�K�rٰפjQSNC{����Ԑ_~����&��F�5W?3
+���ϼ��n?�h�ԯ�-���^�S�r4:����u�$��h��כ�el�r���Dq�'k4�������?W^�9IH6<�^���&d� /R���H{�c	�`���O%���i��@"�d2�Q��W�Пi$�3�i��S3P�K�2"����: 2����w�t���H�b�M	���	:���usW�ך��T�U�*3L��X��ܡ�wry�I0������^8��Hr��($�(!"d��GuGM���7z���Q[��	w<�m�6���L�a\�G3O�itʖ�=�,�_�#U���%�����_���wd
16`	J��Q�6:�D
)"4��B&�GR�	^\�_ z~�
�h�A�����d�SDj��X^N��F�%<��j�a|33��eݽX���hr}�d�pT�'X|�KsEB:@pTn);�X��A��uI茦I��L5�ĿB+��!���<o|�Yks�������}�$$ܗ�\��_�;/�M��fWY��Y�q�quO'����X���#��M����&�;�֏b���������s��I�z��}'���4�ݧ���e�����Иv�}_�U9fRBn��jB	_������d-�j�:���|⑦��?��Iȳ.]�6�d~6��~��!��I�ٺ���\ـ5ώ)��Z��+v}�r�;�.c��X։Nf}IY?SB='�V�E5��!Rjý9���(s�Q�]3�x�]���Dz,R���^��Δm�(X��[�Fi������Ŧ۩$D�3�S����s���������3���Z9�A��|�Z��$�����X6�Oq�sA��oO����0��E�[+��1U�E�RMh����RO�I����Y�&�#!뗝����!1
;.2Њٕ�����ϗ/V�	C��\��L,R���ٟ�&����ʥ��b��=�������D���DQ�;��=uQ��˵��v�Tf��q�"#v�����D)�@M_q�X�iR���#yEU�q[\��X��K/ğ���R`a�� [�.�]ҵ�M{��5	r�:2-�3��4mk�y����>�Sl�l�!_�F���4'�>���D*��k����|s�d_��Nd;�]Ј��>�?�o��FQ���C�u�#��H �`�QЈ\�`�d�$
��3V#9Fe;A�n�F�&UJH�B�����5"��Q~x�Y7�k��K���?�Qts�
"�g9''<_�B�؟m>�XT8��"���@����h��dv?ovT6܂��AaJӺ0s��u"%�= ����W���'q3ds��B@Pg�2{��T<�$<FQ��^�����AF�0��e|J���5:�[)�P�D."m�`�Ԃu?�HL�g������n����zǙDM3g�"{i[�Dߞ����<lzd I��������ģ��%�0��� :$�y�'�3�xlѰ�;9RZ)<��"a(y�sN�Z��
5�8�r�:���[���L{�AwXsjqK^%����0A��麩h"��u^�;�̂zS�2H�w+gזF����a;7�x��uN��S�9�`g���!�����i�5���>��0zO;W�A�W��H���l�"�=��D��h�<D-���-�UP��&��k}BB��u��ʉ����e���.�*�1��Z[�t�I�u��3�1r��g�Jk�u��n�f���KVSX�jj2�_���E�_:0K�.�.v�&�C{�PwduPo5K������6G��F|��&s7�'��ZM���a��>����-�D�.ZT��s-��x&�D3\�1O���0�?��,9��YG��E{x�L�Ji�?���0�N!�����8��ael����m���4S�-%aF=�[��>O�����2j,ￌ����t@Z㌶A[��C���w֜�� ��<��(���r��]�.8|/��:߽@!�/ں�&�j�\�ϼ���{�M����ew�(��hܘ�uw�&���o�р����R�.^��,�=��oa���?g&�Yu���?w�mt���u�3|A�lo�I߆`����5�  �`W��GeU�v�����\{��}۬P/7'5�%�{�B�ƻ�ȅ�FCULU�ߛ�|�w�՗$�i�5�e�:׬�NǑOn����Vf��{��\�`T� X��-�D�~=vZ-M:�=�/]0\�I�Yb�0^���Z�0=]V�g1��(��_�2a�6hAڋ�v5�4�(��;X�֮&��i�_T����K���K��.>������)z*�^��Œ˛z�&����+�?�=Ӗ�z	���Ci�?u��k/�|U�=�p��[u'm�ߒ/V�ӻ���UIpS��Kˍ��]��6����sN�.��ZK�%3�y���!����T>ȟ:I�F���+�q5чEVr\�r�N}_1����G�p��IM�+���f.�-L��o{n���f��2���%B��_�)���9�w�d�g<�q|����R�P�A)�kL 7%E��C�Hqt3t����c.+8���+�%3�[�0yì�j��|ށt>k��ܿ��E%�Sn��X�n:�!�^�V3/�����Αd��:x�D��bM���)C�b��H�e~�F[�wK��qL����А��
r��V�����̢��L�j�pg���%�#��'f�wc�1Z�,���B@���@��]�=s�_Qy4x�	>)�>|ᠮG7����
�d�{?f�۳�xY��#�V
���ܺ$�["~�RV8�8�:)��0ܵ�F�[�����ݑ��)~a�[�VI������"�vR��MsA��T������)��ȁ�1֬�7��3��:Ni���K��V�h3b�ً�}����_t�b�\Le���J�gzuN�C���{, ���%.�v޿ʖc�9�g�8�������Iه|��Sg��S5#�]s�Y[C�$�g�̡��N�&S��B����W�
R�X�w7%�-B�7�4Wu�8�
k�u�9��B)� �٩&Ikh/v�/���:(EE'����˜yj��N�?4�U���F���g�é?- �mR�/0���Vz#\4�i�$���,K9��Ӄm �u�-�K���!�G���Oi�w�B[��T�c�<���E�cށ�ib�ou@��'صbO&��5��ajk-i�n���\j.
�v��p�P��B���lnwB��5`�T&/R���ЈdgW�i�|���I��b�Y����/��.k����