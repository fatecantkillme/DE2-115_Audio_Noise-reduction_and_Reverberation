��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv �|�
����Tӂ���^�2����+t2v�g�VU�r�H$�\%8/�!8�1���1,c���'���c l	�� ʁ����h���z%����\�?�;�=�6����w͸>/Q'\p�~����|��k﯃�`d�C\br��a��D�z)*�&fV��X�v��H�F���i$�MJDK6$�����a����S���ŋ<jN�q��r	-��?��4��✑�j9č�O�r�_���4�l��`���l�M@7���Xf0�����5�㼬��[f>�Zu�*"C���Q-�`��d��E����Pk���Bb�3B_�����PV���f���l��4?U[D07G^�������7v�2qZE4��R�g�3\ĺ2�H��h=q�2*��*K��1�ԗM�=��JZ��cрw�du�)K<*�ٛf+}<����Tkf��!}�ߙ�"���#q'6�KT�r�%�~��}�`"	�q�'���~4�:Sk�c��,>�{P�w�@�PG��aK��0b�����7g���h ���ˑ�W�U���a������������v�>��\��'�Y�D��u�P@��A�uw��
�b�+�?��*�܅Y�~��;� �ԅ�����:{Շ6j�P	������À�w9G�HY�	��x�޿��72�f�m�,���P#�{4(FJ��Ә���f�M��㛗�?�-7p��,���`��ɽ�GQ�ؖ0�V�й�`��؜��_)a[�)��+r��Mr�ܐ��K~�B�N���j�*|�CS����.��'�KY8J�u�,���/�Pa��n��M��λ��
��!?4*��T!4�2�&G�t����|;.���Yt���2}�k����s����"z��9vTd5"��3#��������uf�y���a��F]��|%z!�7/�'���l4���מN�������ǘ0v��c6���0����n9��-GpC!<�m��5�	��MqXV��a���,�
���w��N�#��rN~߆��!�[n�>��R´������)��9��k�L\ƜC�aj�,<�����2#�]Be�
��y�z�37=(�zI����'ݖn����a*�xp�o���G�Pz:J�l�! ����质]w�}�e\��H%�����Kx¼��ћ|Lq�ӽ�6��1�T���DK��k1�JP>�Za��z@cK���\�I��5UX
�Ze��%K���06E1�'[Vi]WU �j͐~�;0P�l7��	-"7��S.e�2"��c���iLilċ1�C:��i��ހx��t\^�[���2Ш�	6J����c(+:̞��� C%�0͘yuOR��V�5]<�*4��Y����r��I��!��lx��Uԝ3��ޓ�I9|�؆H��+ʘ8��6А`�߸U�6|싘���Y��_ty�K�qdE��	�������}�X�f�<�ǯ<c~���5�y덣����ob˗:�B��
X��P�SOh�b:P���(���QH�}e�k�@�Gs�Nt��a�K&a3�k[�v<�pI9���J�}.4X������y�l�^��EJң���x9�s�����.譝X�6��]q���4�����e �� <{����P#�D�*.��2>�bdI�� yr��m]��� �&�����c^�oZzmw�%���J��
M�s�ڕ6^9��;�� H�a;��	��?'�U�rf������b�\a �3�u|�O�&F�d�58ҁ}�{��͐�{u�dĽ����[�>c���3E��Ŗ��͚w�\_Y&s���gLi昇CI�x!����g���'^RbJpO[�k��欺uz9���mx�zzG�4���m�u������5�C��@��;a�"[�&O��	ūP5�cW	�\����� &�;�%<�bB�,)#�� �!p�~����}d�"k8�:sa���i�}�H���Z���^�������5@�(H6���RS 	�K�>n�N��(�u׊(���TL�� j���3�_���Cy��h#q-��96#R=��4V����O6t�4M�Y�]ĎVQb�����.
u�5��Mt��ϭ�p3.�ư��� ����懀ء� ��F�&2u�h�0�K���Q��v���f�A!��?�uyhC����F���߫�F�"�AM�A�0�H�HU J�glx���sth��NvC�ܑ�?G���mqSJR�3�j���3sj����u��i��ש�}�.-�lZ��h��"�
>l��O�0!@o�t)�\��R"C��<�㹴�������1���T4�^>w����,o�*!W���DċT;B}��%SmK(mr��6M�m��{f�"���O�!���h)�c��[Ж��4���|彞Ț�^T���T�?�l�y�������)F%�cGȸ�ް���Z���i뱏H��1���D�<���]�M-S���1�����{1ђ������/0+�)����}_:�7%�RȢƾ��MB?��Ļ[�16R��P]��"^w<��@B��M��6�������v���C�ݯ�i�KIھ���R?������b�ry�h��T���F-%�Aw�����[+�ohF�ܨ3��Ok�Co5�[�S�90�+���"܊hݾ�=ט^�&�^\��3�`-��zbQz\|��C7J�e	qd�!�����q��*�VՈ�T��S���߇�U��q[�m���/�	C���*M����A0x�������8�ʃ������Y�\�qZd��Q�3d�S�Bx�ܥ�����0Y�W��RlJc�2�����O�a{8�(�$�_o�@�N�T�;D�,�^]��"��1�V�:�er��ǜ���M��M�:��GT��.;���$Zc��'�%I\l��k�@Sd��d,�%گAݱ.�q�~��]�4}�U:�
�YM��
�B0�/�pR�� �Q��:�@�J@��{���Z<E�8��xS.�1�4D�Պ��VR޺J>�P�"��Z#�p2H���9a|��aG%�k;e����f�q���E�-^��B��y�03i���a8����x��2拖J�f��:!��G.����z:�����7̘4�ח&��^��q��B:*h�7���b��&H�1��'�b2%��	��*W�w2~��*L���T=�-{�ud��1����=�q��`5��س��y#0;��P������%�ϵX�>H�k�$�SB�o�V�5{�)�Jhh�VV��
�Q�(�g������5 ���Ppч���ŷ�����j/;�U�n����ѫ�P��*�V�?̐�_�9w�P#jr|ҙYl(�~�H{��#H5iѫh4h�PVR�*��{�ʮ�D�c~<�o����crtN{�UnI��D#��)j�4�#HOV��w����r������I�Bk�4����6��7a���#��qZ?}�"4e�>��؇�ה�죱Ru@>�����W�K������N�eu�ܧ���<qT��]L�i�~�@ �z/TD�$���@W�)WPA�!��r�5�|�q��,D���C���)�,�����:���,�y�K���v@BƟr��جkdY%}[��1F�MB��ow�'iY�y���]HE�dlb�'X.5l*.�A�:�����i�@b��}�4�-%{�((��_����[d����S*ɥG�a�)�?_I��Q�W�X�Ț�W>sE�o�-�\!��Xѣ�X�����%�#�u �"�a���
��ꆐ�e&����@9څ+7�9��l��T?.]�Y]��4T�+�_� �|���XQ�;�&TM���(qO�#���6���إ���<Z[���/�u���߻M>rs�r�T�nSHy�`I�uw[���6�d$���<�^�O��x��A؝ѝE�2����,C�}��U��,���f<�W�w�8nf�l�6r�M���J90K�hL��	)�D�n�*������I�@s'.�?2���5>�����7yDWP"�'�8�a��T#1z�Y�sd�����
H��?�� ���G�I��4[��F����8eC3��-��MyD�i¶�٠x�8ـ#h��L�����A�>g�y���+Jt8�Y(�#�TLŻ��yz�G�q���qop8�[�v�6|�hK�d���!;{J��=&BFkF�_��DtF߲�� Z�A(��[F��M� ��ci��,���MC�,�\��s�����s5_}80��<4�c(�pe��6Bw��U���3���2�&����&6YsG~�*:ݷa�K�7�gQWbK�ȭ�w��^�q�Qu;�+���E��iF����Uxje=kV�m�'>����uR��h�BE._4l��.��s��k��P��E�}8@�<���&ǔaI�T���q��M^G���NiPM"�V}�`7� �h�n���-�bdBz��	J>ENy�#��yFHvEl_X�虵b�`��	�TB�mz��h)r&��G�3t\F݅c�랟;��pH��r����v��[�u�����g�6Y��g�N����	�,$E�$��3��6�,^��V*�����鸲�y��7c�������0fQL>�������R�Ϳ�<h�ȡ ��ǣ��ߞ߃�֩H�>2��'|�,�Z�o˕��X�,	��(��9f߳3e�_�}�m[�!O�ZCi����>	�n��\Z?k��Y����y����2O:`P=��.KW�u������p���Rhu��t����ct�N񯒟�T��d\Ii�f��8�xjs�N�f��-5�p)�yM��6H�&���4Qp|8��tSE+�Y��jq)�zn�u�u:�1=��I�@����\ .5[�������wuӍ�:�ü�F�M˦G���\e�Dh
��q��}���An��6L��U�����`�$֒��8��t{2�|"Q��_�B�;���&y6O��[vSQ�3����>'�P/�Ͱ������
	uv{��XN\��
��������ۄ�u��z;RJ�wۇ��Y�=���ӓ�}z	pm��T{(
�o�ҹC��jv<��f)�=q��J��Б� D��%�{���hf�O�M3����6U���e��GB�|V�^6��|^��:n��7h�b}�&�ő6��i�8+�^���?|�V�3�eY��Hd։^����끂�sd��U����9d��k�ņ��E���[����#:k�8o���
��:0̝��k{[.��d��Si���N�]�u����yA������kC���e��*حCa�(��'�˻��(�%6�X�|�̗�E�y���K��f"�Ls�o���&ye�;uJ8�@�t~&z* @�[s�|�T#kW3�N��c<��i�2*����p%qn� �#c)wC��n���I?	zG��q�JmL {�|��Y�ǥ����,�N�u�=��|������	����K���L�&���n��+9h��Ȼ�J��y܃-��V֎�P�%�M	��?����/e+�nv����'}�b�.u�"�w�'J��{��Qp3sj���p��/���b�P�A�I$)�TW&b�_!�y�e7y?.#a���/�B���5h�T�C���m�+F
�!Z�Wؘ��_���C ?FZ����e.���\�L�˴���ƪ����>Z��b�{#`i���'e� R��N)0��?���Z���i��f���A�� x�80�]����\|]�Kw� C���ց⤊[�W�Y���>�z(Z��B���wDxd��Fl,�MiV�^R�|	1�7aw����Y�ʋ�l��(��~)������Z��q�ϝF�u|��-�G �* �:���6e�p�~[s4��H  K���	�Y��@I7�VB���F��w,��5E�/�62o�dA:YID�v���M0�6���%��{��e�7��ѵge��9�o3�`�˱�n��<c��ᒿ�W�aݥ9\"���xv�E|-Uď��m�Iۯ�xL�A���������NDXU��d�}<�)+t�����9Qhȼm������hٍ�fɞ8�s��H^�K����ho��Mw�2�r����W��@��O�1>� U{IV�g���'7��]�y��[�q?�8`�g��a�>��>s�
�T�J\��m�oc?1�Q�B��. L�(�y���ʾ�a���{a����2�
]�7\��&�s��WZ��P �-�n�"�~(R�-�-NՍ�S4�f}XI�c�D(�(A�Ҟ�zq���ĺ�QL6�Ӑ����D�vY�FC�b��T���<
{|)�T�4O�݂XY
d�;��2Σd�߈��f|E�o�-Lg|�"|IbA�T��H1
���+h���cfX���WJv��VP�W�q:��Lpf���)QыҚ�����;8y��jsϾ#>�\��#�F>��h���k�� ���Bo}^�vC8je�e��D��36�`ѾYU�x�[/H��Py.�xts�\��"��
O^`Lm�o%%��W,�?��%2�;.*J� @��$`��S`x�殮��d����Z��?Q9[-��7�nunB_\�檃4��x���L��m�b��B�3��d��*y��e�.�
s�"Y�T�e�FZ(����nT?�n��,N��\d�X����>Uc�X��@�{Я�+�'�2�C�[�~��c�O���1���g���	���wj�	0��]4�Ŏ�F��©���-�$*�t�鐝J�OT[yoˬ��A�N\��m�-W{�l� km.&A}?����a��穎��?�=/���G-��i!��Z{���4�� q��F���?F�Z(�ӓ��v���R偺�>��r��6���lJX%8Ns4�X�k��]j e{r�^�? ���8
�{)��V/Wވ��ųC��OЬ_i�C\d�
k��x����qjv�#̄��J��䡊ư'�5�qr��Ү}m!9�!����Ŗw�cZ�'�P��~����3�ؗ���F�!A�x*?n4�[&�k����WN����tt��r2vLT��P�FB�gD�+}��3|q��?B�j��X����Zc�Yd���g�@��U���R��g���4�^v�|?�^��u�L�����T���r�z��2h���w����H$�2�bv�v���sP�}��J�!���jB�5��{�|1�����
:Nk��������uTg5�-� ��"�~:k�� I2�ԑ@B1���4���w�9yZ�|�T���a�c˳�ϳU�~|���g&tZBmҮe<=�A������w	W�P���{N~n��]��h���}�Oa3m���U����]�!֭�	{/@���2��P�Z��6i��ѭ$�]��Gn��r�i<M��J8� ��qr�2J]c�k��/]	�4.������kt� ��	�W0������1a6�%қ���42L��p�~'����Xw8�H��c�jq��@�ʊ��
�ڢ �?��a=�/1x���[.]Li���I��<Չ�� �[")��-:BpqE���d��������l�r���B��l��C@��W�K�jM����&�����+��,<5#*�e�@�0�О'��?����0;���q��6��h��"�kJ��s����:k+��#�UMK�q�!��t�����U[}����C�w��8R�,I�>�q �3�v씆�ٹ:��1��o�o&��29 l���^��T��{�r�Į�~�w������J���dd�_z��I���� 89���͟�F�q�1�H������T	z9��]�r�|5S��� �]"e�'�򃎫�f����U.���ʅ�8��+�� ���i��#F���9��@+��1!�C(��GA��$p��Tؿ%G�����Gb�>[�'C]a��X�uD���Y�l3^k9���{��\v-�ğ��������CIΔr���ZNiX�󝙉l�N��$������~M���p�U����Mܼ{!���#c���m�RW͢��z..�0��jX�� ��m�<��+��pZb�R�Ԭ���V���S��H:~��O����E����;Y8��{^Ts��_��z��=�/ؽ�����=��"i����.�k�ɂ)�g���s�ɝ��`)x:=�`ĀU�=u��H�R���{��,�#E�(��c��,�Gs�<�0&qD+���ëː��}�Sz��ɂ�R���3��+7��J�Q���GCc��N#E,+✚�C��js�qD�Y�z?�^3���O��@�*7f��1_�2+���O+MB�2G�������?�*���Ki��`�X�y{'=7�l>T��#���y�	����iT�;��;�c�T�6�H�A���X��n����#������E2^Z�M&���r����c��#�\��d�"ZsV����<(Ƃe��p@O����j_����hn�M$mc-O��Ws���yeQ�v��j���'i�o�'r���w�BU�g���L5'�f��l�[W�X��B[ա�t;ZP�x��
� �!)��1�[��F��=����Wm�`��k��8��1�||+�P�g�gL_`������4�52�Q͉�A�K=��׼L���G���
ɘ��3�����h"c�iV�@<�l��S���y��W��qu;�}���4�V��1\����l��=ʞ��U[���f+=��*Nk�ڽAC	�<�I�1�����m!�z�wZ`��5-��Yh����܃��(��� V'uyىv�����G�I�q��%i��^�n/B�+M���x�%��>��Ia���>���X��f(�Lm-'�͡�kߧ�w�u��f��moI����!K+�A��c�����]p�pɭ�vkF%w�?����b��:��	~�&�A� ���K4P�J3��@��(����Y��0�[�s�e�����ͱ+4��3�ȝ5�I��?��g�E��cz�h�����1�)]��"�Qg���m)8!!�h����=9����1E9<':���Ν���[��{W��D�v��A3�A�������0�V�-�Ub(�shlZ����
9��ǎ�hM���O�39��m����5�"L��B��{cN}JЁ=��o������(�QAΞ�7g�F�������+r;��܍�EP����U-��d��?����+(Px	�zMeTɒ��|��,�4|�r��کZYт��2���A�.YS�9a���$�@���VXs(��*��s��V"�^�U�w����G�|�'~9'n�	 l�!�rj�;zF���&x%o�mi�Ľ��{e��I��Mvk�4�f�?d�gEcF���yM�S�����JV
��g���+^*_h��/U�g)�>*ӄIW�Z�*�ٰ�<�A@�2|��k��sxӀ�V��2�jߏۛ�����\N�ȭDS���j\[�� g �݇>��Ҧ��4L���F�Z��V�_֓��IQ8KS��$EE]�����3�h]��-�x�Y�,���K��"�x6��CA������Ñ
O�� v����3��݁#���7�����X�
`9��U2ʻ=ɡ'��ɗ�L=�(��U��Ы�e3�r�y��CO���m�
.<uak�i�EI�zl�j�"8�(����bP��R��4�z��l��ǰ�E�����p�.O\	��1vH_M�5r����Y��(�>�Ф���=t.61��x	�8���n�m��~���V�D])(��D�N�������T�Kwv�iF�}/	Z�/"G���W��W.@�]�Ǉ�,,�W�q���r�'
ga%�-`U�d{��:F^s3�$`@}�s��e/���dן�Ve踡�S'���"�wHR؎�|�C&����U���F)�����>��~O!]'T�Ǵ�n���8���(N�����<��w�O*O�]�nN��~��K�h��'A�߯���o�����=��Y.x���H�-�+̇��mK��,ݹ�_���ov�������ܤ�/�]��K����q���K�B�@���/��u��*D���� /�a�被�D���iKͰz��-��Y���#pԡ�q���:+Q9H�9��P��,��զ��:H�����y���J��7"gTM3L`y�C[���l-M�����*�o��ʕ��0�R�^���&DY�V��H>��������OĮ'&H�gu�7��29 �̻^-���LY�>+Q֯��f�&�����ܙ�)�*��t�l׸��g���j(Z�S�z�pUÝ�=���g1o���?�L���ҮɄ$� ��[���*.c3� ����6�L"��\��C�R��d��9z�[�s��]���AX��*����'��$����h
�s�2x-dPN�6�Q�?ep�E���Ya$��AxWj�DrA�����Ǻ�7��_� 	��ɪM-[�wo��d��7���n�)w;��i�r>���Uk���^�X��4��ym~l�m�,�c:|�m��: n:6��i��7��+;>R�2�	�p�F=���4F�"���6;ps�@°�1�0�Tx	��`t�N�Oj��Ʈ^�L� 2(�v�x$(�U��|��s�~���a%�xT�e