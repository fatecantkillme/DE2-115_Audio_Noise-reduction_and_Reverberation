��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<���=a�bm� |��O��r�5ɧ5�q����� �ni�5��<4�11���u߻������U���[5����uX���Lnt���{��[r��f�����K,��K�#Q��"÷���i)��1�O��*q�WLgR�R,N�՜bE��|X�vʁ4`t���k�+�dhE}�+KBx<�������¸h���K$��tN)=�K��7�jEqWL
����~�����'�NM��ц���ABnH�@�tWF�,ur�Tq��9x�%nK�K�h[ ��w�'�a{*�$�g��n9&J{�,_��>�Oˌ�5x�.�C�ӆ5� Δi�	ޏdߪA�7;��=��Hw�M��/zٲ�&�jH���)R�e)�T:j����o�� m���1E�G*{��=�z��\�`ނ%F#�C�Ե�7i����Mh���L�Aܷ{�d�����`Jf5�a~2�J�Ym���H�ӬTi����"��8�&�~KG����'

�g:vM���O���W,��1Z�:G �/��̧�\	�ᕕ��"u	���r&{�C�"R�~,��L$$.7�����[�V���u�3�@�T'�A�晙-�{��:��5(Yt�ֺ�1�/�K�u��M)L�s�TĸHP��%
��w*{_i2ݝPr�e��H����E��L~a������
�O��lw�|����ߚܼ(C���j�� ����k�|�L*��u{�|i�ݮ:�-�Dc��A��5I(6�����Oz��3>�e_RP��i�_к���WM�T\i��;��C)�����+	�U�!)	���&"�L̊�UgYp�u�BK����T���q 	[���
���!�1$��=�ƙ����>M������i�rY9~�V�P~��� ɳ��0aL�`o)7�	�����W�Z�X��'0�g񻠧sb����s�;��S�]�.�Z^�ӗ���.��������Q<la�����p-�y^��J乻���l��!L��U��&"���7��f~�yjN�MY-6 ����\=%ݗ*s�qW:�sƛ�BCY��G'�3{�vd�U~Y��Z����9
F�БU ������Ϥ�&�j�Yw8��Ǆ�e�k�$"q}���d�TjDӑT�c~&;u����s,�|�n���T��SY3(*�R�+��9��s�R;�K�3
�ȡ��2�Q��Ժ ����{��?��ӒW�^O/�$81��T/+C$���SNH|��M-�,�Hr��,
]��fi]&X^|��z�}��<�i���$�"J_t�L�c��y�PL���{U�ُ��c��)�M�-lw�������� Bq}9P��j:�	��ˍ�{�:UK��K�7U�s�/!ݲ1��������t�z\���܉}0��y�4�!Ԭ�	^Qh�0t��j��/�P@*��)��Y���$"�^.����3��9�oe��܈������A�פ�������0������D�����mR׻��F��S�hL�%_���a�r8�=	��&��,sR#�s���0qBR�������7MF��j�b�,#e�sox�!�EG�T�?>���酇���#���,�|�����ۆTl⃊����S��oݒ��פ��+O���oM��XX������X��T*@�
�;��2ʸȇ���6��t����[a���xg_+l�8^��y�S=�B�*�DO�	MPE+�Kl(k�ѵB�	�e�`//2�c+�Y���= �.-޳%�h?V=�%VbLS�!����҉�a�c�.�Y~(�R;︑��H��P�iz�S���8Ga��y��t��E<(�Ц7˷�6�����ހ��Q�RȈ}����fQ�"���wj~�}�������$�U��M`tg�
�_l�5@^J�ǲϣ+Z�/�F9j�W��C�<�M=�=�#ڄ�H_��Y]p*��Z���Y/�ba����d;B?K�z\r�m�����3���p���P�2	�򵜳F�S/�5�d}�?�U�����;�DWSx�)�R�
���rf�lH�����sd�KT��O�3pI����J����J'�(��j�EN��ӗw�@56���8�Np�'e�y��E|�@�6�sK�"&?�����*��^�r+�Z�h��w�f��Sk_�Чܨr��ɤ�B�Z�$��r�{	�U8c�iV5QЍ+8*i�=+H���V �/2���gFkm��l��y�Po$�#_����I�� h���@M/��p>(	NP�?l���%���%�pA�G�B[���Z�p�n�D9?�/�æC\*�6=��އ˗���GBP�?����?���1��~X2��Pڽ����!1l��o��"v�!M��3VG[c�׆g�o�
0a��Š,�㍠��ێ{��}㵓�6w�JJ˽�җ4npf���8#	�=r�}>g�~�E���Ӕ4�	G�90x�u,Qm���OpٱKUQ���g7��J�z��r�N�#\��o��Ӷb�\����}�=s:�ɍ>Q^��1�hft9�y��b�ƞ����TNK�߂�x��Ώ�	�MM3��*ST�4��?����5LHތ#ԩkw�� �wAϑt�����d�.H�dU�H�+%������d��|/&hE��r�L"V������ ����De���VP�+�2lϏ����`=Y�i���_�Q��z�Q{t��&V�Y���DZ����jt����'Z�Og�cw!x�����:E�`��u����F�_,��G�V_D/�c�����r��W��FN��m����$#8	�*tUC*=)e죨�����o��nI}��M���ZB|s�b)��/�Sү��S�r�&�>Mt�,B[Ͼ��h.��	0�#��핫���	�u�������B̞�G6�M5ƾr����NgX���Ư(��GR���6A�xa�O@|T\�@�[_�E!��D��A���:��/�ﳧm�:��]�����_�A�p�Ա�f6�#����Ц�7�K��<P��2��l#z�<?��LoX5;/�B�s�}�W��/(OC��]+/���tg2��/2���.Ξ4/��+��:���L�`�_��f��ߧP�&�����O(�:
PA"w^�o�e��_���~AY�� �t���a'S3�ګ?�J�\$Cw! ��(#T,է8�\��ť��be�ԟ��@#)�5�H��L��#����l��a�ΫÖw3I�)z��ޣ�K��J�=���Q{�.�yL��u�� �pɤ��#IT�Yg�U�X'DQ��21O����W.v�s�n;s��b�DR�bI��~�W×d�(�8yF�s�ү�d5b�����>|�����b�<ҙM"�N�|�<^��>Qe���P}u�=1/���=������	P�`�"�	�g-��^�{dY`��I_jGt��w7���w����#�Y4
[����JY��E��s�	�j�;,ż�R���+�I6����K����V��.�o�ԕ�Id]��HEV��uC�w8uC� �(h�`�A/1��Vi��鬼P�|��F��#~�j�镙4������i�#�5b츁�m"V����~���C��\��v#sF�
ϺS]�HOA��3��.�?��+ ؟������+�}�r��-dXd���[�_�/ �x,oP��h�"���*�Jpz�gSE�Y|�l��x��g��js�}Ij�ݐ�.��;��+�n��~�^��j��E
04A��]�۸/0���q���=�%�b藲��s$��C	Z�J6d��s{W[s��8�p��i,%�6����}$&y��.a�-i��R"�W�#I|+^��D�P_��F��Ϲ[<��������������a�К��D���p�qBtltִ�6x�#�
e<£�OcMiZ!6/j� _8�ZpP_v�@|��Z�i�}�@����)�����[w��FU�� 2�}�F����\b����P�m���w���r\~{����<#�X��o.����GfȔ{��3���RT��04�����2���S��Ǵn'MU���WBx���/d^������J��+?��i�@p���r=����gs��I��&'ܾ��d�6��!}�%�����B�A�T!%�r�d\b���RT��|�y�bZ�S�\]�H����3q���2��J�>'W���?�[��]�c�kk���ۼَ�
�^}�
7�·T�@-��>1����	=EY?!L=>����/~�x ��
g�8��FD�q|=3�$�~U�5t�6}�Ϛ</�~�?-PN�k�ҽ�N�e����N0I�so�"���b�,ܿ���qs6Tå]��	�4e5���[S�7�3�IP�b�����s�I�l�7�	�ףe��H�-�oۣ�m�n�2�o�� r$�,��j��z�5ֿ������@2�r�%r�D|�e�Έf����q��F�}i�,�����
����CL'��WG�F�)1pp�~��ANb�;?㓢L3�s�� &��z�['�?%KL���Ρ�Y�? B�"o��^W��`�s��^<�?�����#�fc��NGS�q�k�F�J'�C��M]%�zlB��T�CG$��0'e���q����h�b��V�V��@3+�"zTGu�[u��KaS��%��t��	(��H\O2p�O�OA��}'�^������G���[yg�O�í�M��^���>�0�;���sR��9;��m�5�M�;�L\��cAB׈������iw�N7�s�-,��R*�}�KM��"��?�8�Y~��!����b�{[���.������z
<���"+�/2p�t�ۖ��a���1k��z[/V��"��q�V���ƎWE��#��^�T��/T,��g��P��Jm����l��S��V$�p��RX���*M��Z)�������_�k�cv�W�&��9Dy���B;�]S�s���*�J��c�l���\mX�K�ўa�����.ep�u��ũO�V�¡;�s�g5��l[L�x�in��Z1I9�q7p�ůU�{t.x_0�؈�դ�xu]�6�o��L�q�w^��8L�م�B ���,vf�BRjEٽW���kM�Y�b�D�c�ú�a���>NO��'�C'Y�!�A�z; �dt�[ˈ�ܦ�`��4Q�P�5��Z�8�]I��"�%Uc�B��	Δ����N{fѝC�q�fw�IF��g��E羇ӽ�+w����;������X�gn�#o�B�jwh�eԇؑ��M�d&����븻"!zfU+������ú�Pt�1ٯ������"�3:�*� �$1si��^���^i�W��~�J^m���n�%�%+B��<J#Lg����5X�m��c�L��9̜>u��*��)�����w���@��b� ��KP58ԎR����4�&�1g�m{Ѓ��A]��0H�Х�B����:����B!��;�L�S������\�\Ȧ5`W��}y{�� ���8I���<��k�o�SUj�9Kv��#�T@���l%mf�8���OCD�� 矲�cׇ�:���ko������['���O�i$x�o���J��JIv�"u��2q���74����[��S���P�!��P^�vAl�5�_-��)g5-��nl� �CL�zH;_D�D��M/���"�vN�������W�֯Zرm�<�Q<�/�z��D�Ꮦ���4b�Gy1�7q	���q��m4e�A*E�{@� j��L�N\D��©�У��rc*�T��Hd-���!�?{�y��]���#Y��ܥ�5;4_g�6v��Y��y�H����1m$���N}��ϼ죺\�PBc��rp�u?Ʌ�"��ᧂ������ԏ�N�^��"_߈(�\�
�&�˛7(��2���~���7��k�4�:���+s�[x+~K�Q���M<��G�����)([+��m-��*��)#�dN�tTQOb�u5
>L���O�ڸ����Zj����(� �S��=w�vZ��#��cY0j�dpi/��������Аt�p�U�0��D��N.m�cњ�8�0��<��8��:��������>��\<�p�%~��\��p�������Y���?a�#��f��D�>���H���Puŋ�����
T���w�����5��v�O��^�l-�����.��n�Eب�Y�+L���=���T��i�;�	/����u�zz�e1ӑ--2���D6�''5�E�F�>�3^sP����HB3�5�j��1gN$��ή�z�=�|	�*Zu���� ka`�
����?��/�1:�l��w3��η��p�L�R���L����X�Pҙ�/k�M��;8tKݻ�'�RXL���eh́y�1�Y�O�#�����p�Q�e+��Q�F*�p��wٮ7����fʴ	%%��t�)��Q.4|`�2�t-��qJ��.$}�˲6"�w@#B�LӨ�����(q�B�ڽ�S�fA�m'Aq\�;&_��é�ed�-�nҚ=��5�~��b�oD��"r���m�t��!���O�b$j�|����.�_$2@o~��ðS钐|b��@�.�Ɛ�\$�if<���
 몸(�):�����)���i�E>�����/��s~�so$JQ�­�/�+�/c�R^Z8��!�yS<�V�E:�XF��,�[o�x�خ�(^��)���Sp�^iN�������ڸ0w7ƩLdV�A��q����/ݗAr���{ճ�`Z��P�����;ɖ��e9��)7u�N �����q��g�{��/�M����j]!-btP�>���Nw�}W�t[OO�� :[C+� ;\���|@�ieX�AM#��b���b�A�hp�ͭ<{�