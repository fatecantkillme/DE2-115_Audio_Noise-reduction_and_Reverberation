��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<S��!O �&㴎��#�t����:�V��4G/�)Q(J�?���n&LL|t�z�im���4�f8��2�T_��t����KEph�U@��{cDTg�@�	�x�)vϘ����:<���F�e�d	� �Ĕ�ޜ��(�E����
ٰ�BK벎�j���E�$��`@�P��-��7�o��?a��2 �? MN1h1Ht�|�|�P]���/�&#�� 8<��o�����MG�)�;tx�Ә8�EN⥛����N������L6�I�\�֫��o�{Dʾ3b���o
�fS[��$����Z��8zZ�P^�'��BM�8#�;�_�=͟�`DmC�42��䯔NΌ��7K
���^�ѩ貣(%�O�?�I�����2��S(�{��0'�����5���G_�Ӆ�}�Ws�Q텑)��z��#���{؈]>�=+��l'¦��}@zC�x�-,����K��-�����V����F��n�,�b�{5����8gF����@Z�'.<���nKД_̣�_K`0V�ߺ|�G��P�ު��(�ξ�mc���b���SL��"l,k�:��M)Ʋ�_����e��n���1T"�朝��P�4Q�j�_���hn=_p��@R������S������H8��t�ڥJu1�K����+ޑޏN�d��i�&���]I�ZD}Zzvb]A���h��E]�(��4�$�#��Ʀ�_���VX�a�$�B�A@83�2���s�����6H((8Ó�lm�=D�	�O�q� ���@�nG��|zQ�s�uG�D���C�:LL4�m�ᦌ_ZA:eS���]�-��˾r�L7��L����F�qJI�|�+�O�>��ޚx�	٤��1���%�&�wH��)���f_�Z�p,*��Ub:��?m��ܓ@���TbTUs�]���ᘮ򧉺`A�cN�TQL��i�w�bu��H������h�09���7�-���|�/B]�����ȌgL������<,`]�S��� ��,C���������ễ�RӼY�FT��w�}^�Q;a%6�lN��`�F'X�X�}�4��t��C������ 
Y�����N�ޮ��z �;�1	����3��zG��sٽG�Hq��a�)vIA��y� x�ꃠ���D��/̾�,��o����Y���ڲmq=ZhO�M:K�����G�
_��
B�[F���H]o�v���tiE��O&���0R�?���?��������%���E�}��	,��qr�y���}m(���~�놨:3��Ø,q� P.�8�(M!֖�0�X&hh�W�8����dD�����]� N���(�I �\te����FA��" `{�Q�EQ!w�O���cA�M�JϜ���p�1��T�8�픥�r�ϣ�j�􆐗��W�ѕ<6�I��_����Of_�{�+�8��id�!�-�~Sח]�����)��۔L�Aұ�1f͏���� iv��^�Ô�0d�j�k�"��.*BQ�kEv����Vg�u�޻�.>L���.+î�̌�w���o�'��n
��1p��>���@�w��yq`��s&�u#D���%(|���X��IE Y��!"���������e���6�e ߓ�Ι���H�a�����<&K��l���V�b����L2���Wv_�|ALP����?J�L�3C�q\�.��/�i�Ӱm&�����W{?�4�<�e����8�{��ٌ�G�#�W ��Ë;�� 4)e��!��!��
HjG�@�,�5��YLw
%�[�Y��^�7�����H���V��d�?9��nv=���(�tV����э�D"I�8O���D$L�����afX��>+g�y\���<��:�	}�𹕢���A�xM ��h�\+���D�r�G�A���
���s�`	��: hm80~� ��3��E�U��-�n@�~C7D�ҫ��l@��^,|���9�����Yy���Od�k<�#6J=���M�O�q�7N"F��W�=���v�����U>��2�2i;���{��Idl�p�>!$��Y�՟�'��H���RPz!�4ɂ���'�z��Vۼ�XX�=joI��+B�pL��@�:�ʷA�jW� ��"��Ik����5�r���ژ�~8˱a|�/��ly�@��k3�bc���?��%��;�.)���@mho�_�I�(�C��c���&	Nm��x�5�1��!M��	+��
��V?	}���H��f�O�8�=h�����y���rX�G�z�@o�V�x�P��O7�>�]<��춒��:�*�}x�B�G�� 4�z�o�3��Յ����l��,������~W� E8S����~#�.4��D�	��e�~�+���fD��ݔY/ԡT��wO�B��7[]���A�ߎ���%5�rW0
�&,�.� �[o�L:zд�!0�6~��nj��� �r5>���TY�k����x�[SQ&6�@��o��퍊�Y�0VR�l��z�f=:��d��N@o�a�W�
������
x;\g�f�-�r���͐/g���ؓ��e-���#46��X�Q�hJAFY؟nu�Jt&�UD^�,��3��,�1�p���5���ö��ü��I���ϩ+hu���!�n� � �W{��M��+�HVC���FY9�XY��\ޥao��-���ltdD���g	_':B>n�6����T؉��XI���y0CE��,Q��"I쫴?'�
���:�{xM0Cu�F��)�˩�غW��'���|�fJƥ��@h���+���H�E�DY8ʠ���S ���IȔ��%�n�R�D���w;8Z�P'�l�|PT�4n/)���ɢ����������Aʂx�V��=��%"��w���&��ïG�>��sv\��� JfZO�K}Fç ��Nq�m��幰"�v_kL���.SG�=hPKl�BS`ծm�L�ٓ]˲���iW.�y�R�,���S�W6�fY�*(�<]��-H�[K�����A�x�N%��z"F�Q�
;U��H2R�4�A�XubϏ�zk��2�_E���R�}&%�����^r�Ko�V��I���D&��ۚ:�c4̙��O��9�����/��+��?����}��_�|.�k�yr��@��]�o*�L�{�f�n�	5���|Vk  kd�����q���ۚ�d�Rf<�sNҷ^��"�:%
����s�Ga��$I�xn��W��a&�KTq��?�f?82Tᅯ��}�bh��O%U�1��㿶4�E�ݘ�k-����D ��dR��Sdwu���_hMF�9�غ|�ʬ�+�C��~B+"`޳��/T�����}+ަ����G���9-6�ˢ��kn��]����um�B��.]sZ�|�o=�y�m.̲^�R(�\~�uw�Z2z�C��Rm�Y �L���R6v�NYC:��y�j�����~��lV���r;��[��[�i.���AP�xfSk6!�Xd5C������4��� �����3�i�"��Ш��p$�ⱳ�|���R�fqO�q��#J�X��f�Q�0�=��ۺ�]�޽�F�s+�#�^2R��MJh5�w�
��(��J�ۘ$)k�v*th�A~�ؾ��X���E�f5{^�Z��+�/<r15���M��BL#��33���<>|�&�Q6p�jť�>X��J�x&ʨ�\2^�!��8���
���s�v��4⦋��5�}!:�}� �����ɻ�-lH�0�y���\P��air�".���@�r��[5��y��;�xJ8��ﰍ�?������F�U+ � s���OR;�sT��ՈS���������>���
^'<�o1���͒-��k�MO��@)6¼Pc�7�x�207�<���f��J,t��"<�����w2����L�G�jz;۟�_$���d����h��*f��I����4A�# �8]a����䐩�8'#}f�.KXY�һR|��C�#�+S2�ژK�u�hq;�VZ�{�UsV�Z�azK���,�����W�ť�\�[�Ŧ@Gld�������g��n_C�y���Rt���:�5�!�I;��-N'��*�T}{��o�0wG��n0T�����"�x*�ǈ*D���6���%�4�v�y�<�c�	6<���a���'�	7�6ߊ�[�����s\����7Z�HM5�c���.�ɽp�$מv*y�����O�#�k���Oj�J��3���ޡ�_�~�t��o$ޢ�æ��v�k_W�C����@��ဟ��߲��bQ�Z,?��R��@�ln3��n^x�}^aE�8�.���G�@��1�v-(޿u#LE�����e��Ib�>�kqw��SR&f�n�E)�b��8�?4�Q�v��V�1��^���p��K�<c�cy�E����-��?�n��&�*�}఻$0�D��!�].L(}7��ڟAO!/��+7Sa�k�ǥ7xb,[�������"x��D�d������N�� �Mc�{Z����Y������@�Lޛ�~׶s�=-�̘��v2Z��q9J�����U}R<B�ՍP6�0!�����3��������<l撓ޙCB������|1�	����F?a��RF��~�*� �`�	�=����Ɨ�/[�Oe'���N���D��+z��Y��[�eE�ߥ��'��})�#U�K!ի ��I�r��n�����J�)���gQ-i<���y� T\oT�E����)!9`]'y���c����5y�0��;e��C�:8X�J^�w�����| ��o	ɕ�OY��T����2J�a�TͿ礮s,�o9*bC��7��U�k� ���)P<���5̉����l�8��H����!��@��dau��EI�ު��8~�Nu6��3�G�Xp����WIP�F�Lg(�ω��H�1�B0E�9(S��`�U��t��c�H��]���TI����C��421���x'`��.D@cst�A����YJ���`
��j�MQo��`�dTv����z��������i�3��")��G@i���&k���-f���sĲ�HX��:�u�ܔ+�<hny�1��93��J��sH�_�R�u�2���1���X,�i�y�!����-��,C�������{}:#qCp|�z)��\�=)��;���ʣ�q��݌ڻj"��i������a�a9�+�:�v��R��Z�{��2��:\��ߚ�5Ր6[�t��vK�g8� ���^�]���7�Y8]E"����m�����=�H�$-��û�@v�jA'C>�*7=�e��u�5@B�O�@�"�x��Ͽb'�{2�����$WL?����kP}���y��Ky/��?C[�f�l1 B�>�Dt3�H٘��G`WE+<P�����Xڈ}���}Yh�)U�)sx~��eUdL9gY�5��ވ��71�<j�Rh��F�8�
)�?�Y���z�<c�H7�6�\/(tP�'M��CG�#���e��9OaT���܆�˥/gݱ�x؃��o8��k���Y��S���]kʕu��0;��������!�f*:�}��SJ��Z����~��z��Y\���H+�%��Zy��b��s�iV�K8e�ƴ,ׄ�{*#MN�:���xu*�^řU
�g�kj\�^F�!;��]���D�K�:NI��'��A�InT��]���8�!z�����S��0=�|੸�f�t�i��X��B��O�7z 4 �n,�u�g�@N&X���Ìq��0�*���f��!ڬ�r87��}����~�ץy��{f<���&FL����	$�P�cvV�\������r�;���c(�(v�ړz�}�N,7�i�U���.]��@3YҦ��z{R\��."ɯ�_:��a�Ǆ�7��l����(8�u��<\c�jK�{����LPp�m<�y�_,���<��N���H�DM��,���k�h8�2���v���mZ�3�vh��^Pm�<��75����5��3	Hȑ�p�P.�t��ʯ��K��T0G70�Tw@.���;��χ�VF2�؅�	y�W�7��(�O�w�ӝ����b�J{ۉ��ڨ�F��,�4ePo޳����U�@r�̪�L�����Q�㮅��5a�`6���_��_�>T��,D�	��"�w�Ÿ=N��`j]L�@lkN���d�'����ܘ{A��)��h�.�W���(�Ӭx��:>11�G{ЌF��\�����ʡz(^z�bK�
�v)�igyB6�����s�)�<�o1���A��ټ�K���)�k/[�@*Oe��X�䪸�8h_����tu�C�^4X�nrq��b��ϿC������&	>��JlJg�q�9p���.�)+��u*��b�CwJ��M��T[=˦AO1��-o{�>�UL�z��/f^�v
0���؅�a=S���;����t���(|�������r�)�{WF�9����E��@�\��L���0��$=�CU%��5�t�5��HA�������ڭ2��it�����8(���3l�˓RG�#�ˏs�HH��Wz�1�س�m5+����%�ۇ�z?>(��XK�jű_����MA
4;��R+f��M�6�#�˛טX����d{��V�ʝ�&Z�ф@���K}� m�4ޕk 7�Z+|����8�|�e%��
�ΠWhb�q	^6h7z��8vSG��Fwe��jL�[v	��ߟ�
շw�k�˭��k�|�F�L����7P1̼�]<�����T+����6fKG�#�N�h��.��>V(��0�ʅTԫ��M`�P�]����JZ�ْ�!��K��`�-'��"Ss��q��T�Gj�b��̩B�}R��u���x{�u�ѫ��F+:u��O�
s�X������j��E�:=E��CUᳬxw׾��Ug���w�G�_�}���t��4 -_di��u^���Kd�J D���O���/z�;�ʀ�}�g~���G�jf�~x�=���X��9����x����.[VC��yI�Xh��Lv�o�MzEZ�� Cz�k���d�[۽S�hxkm'����,�9�>��Z���Ӎ�0y�l�w�����7����ė�FuRu:)��Rh�������H�+5�v�c`�ζ�aF��ֹ[��I� �5[s�4�F�y0��g<�f'�cw�� �]����cE_E3.��v#������C���F_�١c5py.'{�*J�F� ����5�ήM���	�Շ�ۇ��1����FCN@��6��9�p�����$ם�l��S$���f*�XE���@���I�ޯg�Ξ��E�i��s��	D*�wprl%^W���v�����Ť���y�g���ſ��w�phD\���� 

axҟ�0�m/�i��T�Wt��楱�!��VGd�`{m�P�/����D��Qf�� (�N�e&� ��~��G���I������{����h�!��_�um�=��v	�Ʒ�}�*�ɡ>�)��4h�����w(��4ka����~>wB�"�]����p��M(�0��@v>��?cz�e"���ٹ|�*}د):�O�����UlH��\O����=�ڷ�fA�S.|
b��y�0M*T��w�8w��6'��vX���<�\�9+�-�wr�n�Kє�hZ/5$�����k8\RQ��6lB��`P�9���&V'���~�2t&�ʮ(��1���h�� 2�T� 7kl4Q�h\��Ϸ��}�Eٍ�]	`~�3v�����E�y{� �=���։L!�����zT�ļ[�F��d��߾4�c�r-G�����˚n�w���s�7�s6�4�5
�ۛ/����x�!'
�z,��$�_�#t�ؗ��p�:�3����N���$�����h����wR/03uCsL��;�ת����-�x=�`�j�������������I���^v�o�d%G��Z��D�Ղ��b�ڮ~�H\k?�}���|�?��O��$W�^�d]z���Z�A6/b�d��=���n*���Z��[�rҬ
�	{����9
W���G~?S_	�m�Cc{��vl�%l��?�FT
����;5��_K����T��%�Ji�"#p0w�.a��:8dZ�oO��\��	c�Y{%��$e�3gQ�ràIv�:��!]D	ʂg�:������'#�J��j"�;���C�e���U��>9��x(B;8M1 Ax:����k�L�O�i �(�s3�����Q�4髗`���u�N1���@!Bò�2�6��Ǻ��Y����Ӣ�#�j���:�
ݜ���Xw���������H��ʢx��~މ/릌�Lꡠ/�Fʳ���߅��c���6�.�:�? ��U�-�^e�*�PLi#5w/�ۖ�w��S(G�j���a�Lxj��¯[�W�2 /�%�dLP�aTt;:���(,HB���Nd������4$%rV��X��#^}Q���'�X'-��1�Oe��wB'�\+m��l��� ��qilǆ}2lJ(aO���!v���j���3�s�`�u���:�¾5n������$���������O�]�`�]�����=�0�����':�Z�d)	��a�C �qQ�0��da$)JW�z�+/�@g��Դ>7KE|-
Ol�����zJ��Fn&��Y�.s\��h��<�ͮ{N���>Os|$#��l8�����-���A�VJՁ(XT����M#��I�=�oή4��^]�!@���UO{�)�ڀ�QVzϭ�������� Mq^�tX�"8 ��.����|\�	-1�u$�jf񡶭!jR�����ٿ��.���yg+�D���O�>R���T�55��*�&'Pr{	�~���<�g� ^�1')�����hl��{�Y�B=g�(��_�d-WH��T�$�D�A9flJ��*��X�'b�kXk����3�va�
��b����y]�J�J�N~�V�����sx�I��[���(Fyp�z*����F�V��}�е�uy�G����:��0yB���*���>��t����Y� #�W��� �d|�t$��8��g�.Jn�g���v���m}�"���yf�M���]��U���T/צ�>�M�\i��� =��b���>���@�`��ұ��v��2�sQ��ER�ʨ�A��w�4�&�3��r����C�%��?\ DY�^�9mHܜٿ?D��D9�bf���=
%3VG��:�94x6����
���Y�5*Y����b�ӄ������Fd���\=�w�Xx2������3���`������21�M�U����������Ӯ>��$�� 5�?{E��)�_�66�F�J�4��'s���=��t-�qT$7�>����F�uD�
����v�\$���,������h�A��1A����-E:9��D*����$=H������/P��W�)�3纙%�Q˱2�e `���J�ku�*U;�$��Hod���u�78��?��iک��5��ќK��� ��i Y�H�K�N�QJ�2v��q�D� �Tg��oz�+v		py'�:j0�(�\2) `�����Yg�0��h4k��<��iVezʰ����\��G��Q۶n\�ɫ�T�Aؠ������G�|"}�ؠe�
������3��b���KU��s���`�毹Ze��^hkp�6�� 6�;����e���ò��{��+C���u߅;��1u�9�T*�EM&���k>g�q`7��U㥹��ll? f���������Z=W�K����/^-�.�cTa�ՙ�����F�{���|7� �F���!,8ߘf�R�M�Y,s�?�ߊ�ԧ����M��ॏ����:P;�S�P��Nm���v�C:B�`S9j��>��ֱ��1C<��Y����ô='41]K��N#���.��+.NyS��K�č�9�)V�	>/k�?vw_i'���Y�K{��L
v���D ��+qΖ����� [>��ͨ.�8�ɳ4o	�����_i�gr�;3SA%�T>�
�eƿ
����빊H[�) ;���K����j�� 	$m��r�I�����K*
 �=�K�@@6�6�#;�_v.F��7݅�
늯q謢�Y(�e��f�%�����7E�3R�i�!���ZHToɃ{�^\����Y[��藒d,���h�(�XI�/�Š���l��t"����i�d�-C��&�'��l�4>���+ yӼ�C*�K��@���fD�ܴ�v���^�rPMj������o�IN�T���������izS'ٲd!�a���K-��7|[IL�2���B�:	�5����n��A�F1�>*�=�����YW�����
��m�c����m|v�=a��Zh�k}���/�/���$�ͦ����c�N���QU3X�r�h��m��?��'h�ڴ	,��(tu~ԇґX��K�`�ҏl�c�^�2Q�#��V��Q���Z/;�´����0cq����+>�g?�ל����cUp�O"2:>��a�����^��:��ݎqx��A�.���eT;R	�%�P�M$-e��>��B�5�����\WN���0�7�.�*�{�3�䂺o���\�[P�y��7�`<�(Vi i�"V�]��PtZ��װ��t����]T-+8�'vʅ�~�öai���n:�S��N78�#�� �C�7���34y�*�djFڒ��v;�4�YDHx����~�Ռ+�jgɤ|(�G�Kk�Ô�V�~rQL��Z�E��I��t.��\4��80U�+�@�Q��j�o�/_rn��h���b9�H�#dΞK6y� ��S�-}�&%qs8�W#NE^������[V��]��Aڂ��è�?��+x����$����zoU�+��z����)	/|��K��Y�F������Z �%?(�E���ڳ��2���J.ʾ؉A���|!X�Ɂ�&�6gq�%��"�̉�\l&�6i%�i8U	ۋ5��9#w�K�>k���)��p;����דd=Fc�Hu�k?�p��,���\�Fo�<(�|��$D�E��M��(����Ջ�|����O-r��3���u��y�~IA�+���;X����>�/������(�ȟʌ�:�6���;&���7�f�r�XP1IHǻ�H�{��	�rw�Y	jmޝ1��af@���L��_-�����}!��>;��+;�N�%[�C�xxh$�sN���K��f���0b]]o�5����6�zX�q����R�U�A�a�����+��۳I����� ���'�o�yy	�8bK4z�?�!G�t�W2t�E�����W�pV�3�����w�7���r���ض�N
����뽲�U΄��c�`�9AƮ� HͰ�i%q�����c��Wٷe�r���7 ����`�X??�홍*J�y,��B�@�A��X�F�͠��r�b���ud��}xc#<2���Rܶ���|��'[9����^�+���( _V��y�QO��lJ5B�� �O�2�Ş`NTN✯2&� o�����|��ad��WAX��V�S�� y��̣�gu9)��F��U~sv�H�oI��"y�1h�p"����.φXP�ă�v��)J��sA��y �p"j! C�%�Q�Qo��rH3���mc-��Mp�4��n��@dƭ�cv���i�fЄ�4E���2ɀ��4�GەF�?���<�KDv͌ �iO,�k���x2��P����&�<*>e"�g��w���A�;��/�e2z-�x��3I�v��3�6�f�oa	LV2j	Ptc+�z���=3��2���%T�:����.E>R�Ā��������:o&ج���1�'g���l5���L�"3���5���Q�����Ӓă�
����_"�%�9I=����o�)��"8��B������Ꭓ���Ҩς@�6q���J��)U3�/��X�H��'����6LH�w�ב+�oM�0�~�5d���vf����2m����L~�M��D���+k��e���h�����h�/��&Us*D�"i�У2X%.�"�ۻ�Sy�����?y|���X��@V] �Kh���W�����;Eq;��^=|����|�Q�<��>)�x����C�OKsd�`;�l�c�8�2>�'(Ĳf�R��ذ�ي��{i?��v~ݐ`�s�����0�\�#�o�*�4Ѩ�f5yy��h�շ�m���_�q�����in�_&�"����J*�Si)j]	����gۼ��QjBʄwR���M��P���<j��ڎt2Ώ6���An�5w�z;�-��`'3{��ڶH�8z���uLM�f-[���1���}���ȧԗ
�~�֪��϶��W��$�߬���_�x�,O4^�Z�3�	��܍*h�M�ӯ�֌�4lX��hۛ��6�Fy��e*gdm��|�C��տ� l2�̎�t\��@��E"���<g����?���-�:�&�C�����@V��˥�!�.�L�Ɛ��
&�`��i���N����r� �!�O�(�b}�ܒ�b &�f�/x�M�eq0H�S��YQH�Ϙ�&�"�r����2�v(���/���	@n'��!D��q;��\��`"	��x�����Ɲ�Ns<R#��̣Б�G�H��a���Z-q���
�gi��YZ���T�r�H0ݮ���������j��X"�|��|$2=���55R;n!�;~wF��;��ü0��ct)��� C�?j�~�#&}��4�]î��ڈ��2�����Ɵ9���9�@�K��5�i���|&�K�&�>�QG���D7h]^}Mq�dӫ��c��g�C.;�����8����>�P9`(+�gY�a<��@�A9��T%���Ʀ?� ! nW�JBW��W��S���0e�3��c��Y0��h?��/����q���4��aO�2U���@b^k@�ռb�$�Ż=i���{Fz	"ǋ"�����r�t��R Gnv�ӕ�����'��@}��}~�a��Φ�؊�b^^I�>HV	mՀ�J�>"�<�L�E̸&H:M�Ǎ��i�9�]y��
�;�Gd��޼��ފ��J��6#���h4S�uX��`�����)f��F�^�ν2+�Pr���f@"ޮ�<��ښ"h)�G|W����Sԅ=D���sn��D�:�Z�T������A���cꤊl���UR+7�N/�X6����Tr����N70*AmO�0C4R��.�K�v	�1@�ځ
W���Q1��_=G(�c�?y��4��-R9�A��xʿ?�Vp2�Yk��q�~�U|�͏��J��	�Ⱥ�=�:������Gx���� �`��e����4#�L�J�#��q�����l��i�T�0Q��Je*��Y)�%�J�8�q�W�ىG`ݥ#4����x9C\Z���-���ɼ��*o$�T�w��]����jTX�Zě+����q	����:]禔Ҝ�Sa1�n$��{a��K�3����B�2���]K���*\�E.��g] ��9\GiS���*A�A�;"�F�"��p��0E����_o����~J;�~�,�L$��P�=N4��{~�>���T�mz3��h,���9W�n)^�8S�^�o�XA8痒�s�#�|:�y٤���c�)
���|�o�{o�Xѐ^�N�ۖ?�[.*J4�i	be�b=��U"���P�@�?���{x��>P���6��SC"�D��p���M�����x/(��+u����u�7�������;2j/�I�y�&�tnE@����M�{�J���+X%p"��iǘ�,�&	��r��8�2p�)�V�^t���?v�ŀ�T�UR��`]Ě"�)'�B��zr�+�Cu�U�6(���l���억�6����Z��a�ZÃ:��Bx�a��h�� qX�ߩ;O��D��KQJ$���ע:�r�X'j��">�/_�1)��"�B��Ke0b���Mz��A�T�~��g\P��\/,��Ef	|�N��cE��r���[�2T��u~�V�׺��n���h ���}������U��k����P��k��f4Z�?�z�:��J�{w{�U^?��\����!����a����?u�c)`9)�����#�p�v��nKs�����o��R�KB��\��>�D��k�p,���Z��]63�R/���k�Ú(5����o�W�fs�o��z��`�ߡpFkf �U^6��}���)��1�?���Hli�K�Zkd���G�Z[���R��w��m:�h���U�@�YG�gT/�	��FN��:�����Mo����z���mu����[��|~x������z��?K�>f@9U��]�
�g�l!|�I�������H�	d�S��Ժ �j�7u"�:,b0V�*�4-e�^�'*�J�$5�D�)���_,���X����E��0���κﬃh�����(�xk�ۃ�Z�U��Bz��ɼan1АT��c�<#xh�>s����������ӎ~��W���x��.t�a��垿v<��{?��C=�ÖāA���Ƴ�PbW���m�\����$��>L��ыE&\S�J�3�W��)�:#�Y�����c���#� #'���b�+�+�g�c_:����&u�s�e��,����YJ���-�3țU�t�!�ur�y�Qƽ��I��k�M��46ԁ�q&��.�t3���_�ǋ��3W⊩z�т��-�q2���XF����bp� ��f�-�����v���d�VO���O�1�	XT����ʬ�*~��b6y��.ۢ�t' �����y�{��*ꆭۍ����+��Cu�=N�Q�~��_��s#�%Ց�-i9�b>0�-A��	�	��n��j��U׏������^)�_�z�6��sC�g�Ci��B�-䉇�;�I5�Oa@��t�H� t�L��=c�}�^+c���W���_X�����<N�[}
r��!h��� �-: ڈY�ǃ�zq�de�[�q�̗g^�۔G�I�ؙ�#[YǾ#8[=y�g�2:9t�6��H6���Ū�g�����5ҥ�nB4�Uv��Ɲb�C7*�Y pL��9�����>ƽ6C�S?�?��������4tC��i˴Ck��'J�I���9�x`�춾�0�e�9E*io	~�1m�W9�wj���D���~�E�(�6���F��f��d�#OYl��f�;��]��Z����k������}����t�a��ۻ��S�W��O���Z�/��}t�a��S�*bvw��b������+g��	3,L�Sf���":��Q�,�P	�.�Rk�
��b@:6�tc���V���~%�>�6��c�g�x�Jas8 ���ENu\�?��aYZ||Jj��,cŦ˾@}/��l��ⵢ�L���5O�ޠ��my���w���HV)�0�R��-	����ȝ�� c�)^����o��9�Lת�\ϘC�y�~�3�5����l'U"G�LzeU&����߾��s`�'Zx �����w����{6x��PÈ�\_}2�Ŝ�������V������$Q��"�����cq�h�U%��ؚu��1��r`��a(��>.�_���e�r���7�����#˼����k?��T#�8DK�I#
��������UybW,)*�0�j�3to�߰YpC憥�h��b�T �S�.��'v�Ԋ�n�יݝ��I!�,Ug�7�n�L��쑬fksk_%\I��g� pݍ��n
�68��CZ/8��,�� �yx���#aI���z,$����/����t�@D���lkpC�%��d0���Q�ɯ5A��F����֘�y��"�H���»F~M�d �f���^o<8��~������z�5§=�v���g�hq�+̹���q郡��gi2�`?����{L�m���4���L5����ӷ�'����R;��ι�0� �OÓ�PA�WpO���=3*_��r\�+a�e)C��������ј8��`��Gl���%�|�hp���eCr����x��,�W�3�İ���n�,��#��3^~D� �W����BEz�I�̩�F�M���Y����je+�%De��]z�x����{�i�{v-���Xk�� a̾���a8�5��_��>,ɮ5r�ֱO��(���
�$�2*ʭ����l����2�ȼ� �l����Z��f*���4�U�ś�ڟ�z�Y�IAg#ɦ�h+%o[�c�JPm=��b�)��ਈ���t��Q��!ڝC�r4%��C9��ǃ)��w�
YNi(1 s�ظ��oe��]�"�$
V�P�eD�����a��/�c��.��t��Aw,�* ��o�r�[y�.S�5��Zfm*!���zC%�H6�ɽ#h*�X&����E���y�\Q�@˒{i����~{M�c&�MB����Eȳ+�`�+�9�:JtE��m#�g���[�;��b��s.�Pxj�^.��PO&�έxe�=ݨ@|1�>jك0y�Q�*Tk\�8b=�I�K�=���D�����+���q��!\��Qh� 1P����Ut�r��v��n��^oa<7�Z�Hx^�;��Xh�w�:v)�>"�K��m��Ǳ�W�\� }/�J�h��+�p �
2�V�����\��׎��=v51f0J�_1qQ�q�����PP�W׷�UYK��R$���џ�S*��}%��>�Y��{�Zm��_ ï��;V=���ڲ�>Ɉ��Kȏa���翚��=�[3��Z|�<�N��Y"Ŭ�W�%\p�b��{F�O��j��7#;3��z���pV)@C'|E�ǿ_R����*
��c�)����W��Q���̬2��yv�4��3fY�W���?G ���)߫�6��u�]��ɿl&�d�~ڀ%�('-���ƚ��5#0� 3�&��I�C/������?�����^�s�'�R��+��xc����S,L:������)��ݠ��I�u�BE_R�����6��O��Nt]?1U���Ϊ�7z�i��M�m�qI�h�G�~L�Ѷ���C�O<�jUJ�k0���Y ��W�O��2��L
��{���dzh0����e�E�\�KM`��D��%��e{	tv3����Zi� ,j�M9�*F��ޫ�6
	�������3`�9�t��x�ڷ0�t�>��3��V���i=�
��^�9��]7�����Et�oF���ۊ{Vq����{t�FQ�7��,��?(C���oq{���?#�n(A��BC$ZA���IO��ʊ3-C�%:�XΠ|���=�~!4��ePrD����l%�9-E4�vh�m�q$)�_b��sjC}Y�e����R{A@p���\�����u��ο� .U��A���A�XB\w�Ȕ�&��>c*T����bed�������e�`'�{�zy՘�;mc�ՐԵ��!S������]����EB��z�hL��d���L/�L�_�v��(��(5��p��4����x�:a����L3}IcB�W���
����[L��p����:��>.���i\���ݗ��K(lCx,�5�1��'���O��6.�˽���ͤe4�<�}ϓ�<zU��Z<��t����X9��4Y�����W�|�� ��� �����q�H�ˣ�)N�zyd�"��7���N_u�����|�F����3	�X[Tǉ��V���VR�����7��]��j�%�wB_w`�N�R�0J�$�vsD)
������H���q����e�m9���{P��ɜ���{�PH���0��U�1�eF�����qb��g���?������풵���� 4KYŞ�^��]��#�_'%�{D΄�;��T�V ~78�k���V�1��s�y|��]ґ	��x\5��k�W=�=������G@��k9Wm�m�Kp5#� C�s��q��<���?")!΍�������5'��ϳ􍱯a̴���A~��́�8f�ϖ �a �B.g6�a���!��
[�C ���L����\=��u��L-�W�+E	�:�����O�X���&O��hQ�W�=��Q$���q�I+�	H����r����%�e���pI-�	t��ÿS<4�5���z��6^�+��#9��^�yv�6��j��7]8�L�G�I�Ќ�V�Msg#�kNW��Wx�@0JG�9�'���[�M�?Ҡ3z)Do��9����Ƙ~� w�X!�x����Be��#ɽ�5)�V��x!���1�m���G�-:oX���$� ���`��h���WBG3�g��Q׽ْ���T����.�hoPJ��}�z�k'Mq (����X�����o|�W�KG�����X��i�"�0[�̰_�z:&���p|���,�{�Rė[�3{5�֤��^�9��f[LP�M��CV��-9��M56�aT�>�=�g}�\u�ӳ���z��:Y\�{�RM�bHX��n��46�c��'J�f����7x
�]'���,u}�[L���8��V��y��7�9�QU�'��6y�EX�U�I��19�B�ܱp�cػ>�ޅ����ƿ��xl�m70�Ⱥ���;�x�����2��u�]��CY�J k��f��*v�I�Ĕ��q|�ݙF]Ҟ(����L�dq���sG�*3o�4C�ʿ�s�<���HpO��y�������V�B`��[5g�l�=hiW�ɾ(�	�����$	���ԆcS2�¾-
��b��EK3ĕ��*�}��A3'z�Pg�2W�f`wp��)۪cQ��*�}��X{6�a�_�y���Y����<��95b2C�i]W)e-�ዚ��Ú\���Q-f-�g[����!{A�!��G�����ω�0��H��K�\�+M���pp���d�HG�ܠ��-���n	Av����y*0#��._�뎠�����N&��o�����' �������Kg�_s� �b7RBx��c}�x�=����݀�r�	-��#s`�ʌ���F,��(b|�����\��d�y/;*��u �'`GP>����S=�-'��`j7�j�܍��E�-)� <	�j�h�b�yg��O�].�Z��k���L���cTL�	��#��h,{nPKy˲�Y�)gӡ���oO$X0����w::T�� ɑ����6�<X�u�|�١�q�R��DM���~t��{��0�L���~��_8k�N�	Q�S�H�y}�� NFl��q��<	Pvy��)1r�R�Yb��ђ�FC��4x�����d���,|Un*���>��}#qw,�$�u�"�!&ʃtba�{�~�=?1G?���bY�m`������3�"���G�&���+l�{�%�J�X_�����̤�@+�CAD�n9��ϲ`}��(��󊩱X�22*g��IC����Ű��C9.U�G��}~�5��%�o&��O�q��a&/4� E6l�� $H�R���vm")�4�(����nݟ�MZ�$3q2�HOnx��� -Gu�_̐���B
f�V�S{��y>^ϰ����ۍ�Ik��3�UAOH�vX839O�`��#e�EX|�T}�~�Q廙�,W�[+b��\I����?��&���ǧ[f�!�~	��G��B�z}V�3� ��Dk�-�>(Y${��:����>��-�m��b�.؊P]�z�-��j)�� ��9{W��mU��7ʃ�5|Qt�`
<m����v�})������қ� ��u$)ٶ�C�?O9,�lڇ�����1J|�C���m�_�/��5$6�e-N�!���9E��(���l�ĚO56���$y�j�zvv/���r�)M�|��i!\�I��0,��Cs#���>W���Ƌ�\61�������\��<����o��-��M>�
����<O�����r�M�c:��m��oJ^��4-�\M�WHNB{H4���@@XWk�B��p�c�''Vd��I���`]�i-��ך�E��� 8Y#��,_����C�H4��b�yyE��rH��aLEr�:`s��:�������FpB"аlx��T<���hn��6���Vgv'V�r���v�<HRL�U'��w���/P�Fבk�^!όG#ir��F�>��Eᦎ�X�i��rk?��U�/*�uM�Y:��C.����Z���D��c��y8t-�~2�b��D�"�E�т�X�O�V�x��2$���+�FT�[�C�	�^}%��g牙�S��HA������8�����D3�|W4����F�M�n�eYZ�bicH3�^M�,:������U���T�]�����x��8�z'<�[w��Y�C�Lp"_n�r �I��0�|>N6�{PmkM���ڢ�̅��C�@�~=���{Ie�<_�:�#�D�%��t���i��Eu
���zK�ƳA���8���R�g��U֫��V����9=y�aRh!|*�p�A��mg{��s<��v�0�L<����W A-нU��ɴ�
Eg.��6�ʡ�_lՐx�<����3TdѸ����K�ySν�����t�������8m�:r��e���Y�#|`�
/{��E 	b�]�?0as�����/���i�[i���e�6KpǨo^g��]NGq0-�`�c��,�Ig'��lPf���	�N�뻙��A��Yl�ވ��F@&���>c|pW`R�bp S!�ܴPWX��C$�	qޙ�.'���2�T�PO�|!�Y�N���g�B�X��O!�+1��ԑ�!N�%;���$��! dd���je�=�K��}���b�q���U�'1E����fpM�J�%l��T�-hӦ,m�0-iœ��{^G���@�C%A��I��ܿ����
� �(�q�I0�� �kJ��8��j|y �� 5$����o�~~�Q��җ����L8q���n�w"\p�ҵ��$/�H߶`� �[��_��N����d6�����*_§�˷%�S��>��f���q6-�<�⮞n7|Z�Bg�$�}O���P�-�)�2����"�L����+�/��[@)���� իN���c�Jb?_F޴rU�c�B4���h���0|S<rv��S�[	m��?�wPכ��R�"��ڿ��V̀2�\������+b���o�4��x�I��� %�.�L)JJ쾎yD#�$��"k@��"��ӳ��1LL��1�{ܖm���sER$����@�88q�QX���� 2l�|�}�p���l(���b$��RJU�p����q��ʱ�5�
F!�AJz�څ*��9����s�Z�Mwb(�n�����t��@z0��f�L�D�֫xm:�}eڇ�]YL�����&2�{�d�D�a���@�js��`�)��ǐ�����t�Vc�'�Ɣ^��Pg3t�����s�~���Y㛲����>wi��� ۧ���=����/v`T�I����΍�,����&���q�l���H����a�F�gg�ǰ���u�K~�N �ܗ0�"���8���������M]�>�1u&�N�.4^�נ���\z�?N��΄Y�K!B��FzaQ�\�B�/Ƹ~g��ݭ46[=�՞1f0�������6�I��&5�q_���I�g�r`V���Б�X���}Q	�U�'A�_�����&Oz��e���f���npT*���U/�+r��~�֬0G�:�ά'�)(O�Ns�R�`�nKc�5�������o�q	ꝴ�*j�&t�מ�_1o����@KV��-z�t�Ă���&�[rx�|ck�=�v��mU{h��-�*^oʶ�D�0�o߄B,��ByPk��Y�Eb�ME-�㎿�%S��+eɂ�ou⯨	5�_��c��nd���n����$�O�3��H����j�vP/�:�(BH �����7��Fq,;sG<};P�u~:���3h5��sW�?����Ҝs�\�W���:ɯYR�j3 ��ke�`�;����5��M-٬�0�o콻���eW ���-&�B�n#��W��Bڟ� U\��1�T��cr���B��psπ��7�Xv�oh����I��I%&l�m�(K�1[ˑ��03��\���0��G4b��Ǝ����Z����vӋX8�8���E喳W��9M�ˏK�i[?�k�������9p����p��'�M����Uܦ�>*p�v�Pe�����Į�߲mU*z,`_�.y�ϯ3�8Z���S�*;�`�̇����GP*ŸI�O�u�kPPs+��*�t6O�ei�>w���'/٣���F�n�Ҙ.dv��r���K�|o��H��r��H"=�}��cO����5�����<MI�W����J�'�w?�N���h�s��u�y;��vO��_�,�ĹMn�,��[Q�C���i>��h��M��d�ƺE���c���
U�z�Y��#�SW�����z���1(�S���Yø���I@s��^�T���î�I��s�~���((��=��
*7M_��H��I�����%Qr�9���DW$�+�X����J!NYZ���;0�k�
�v����e�.�o�u�[=�[j�17Nm�Ϗ'A��Cm%����MKq|�����6���mq�4+s�5Z��Jq�.X��|3e�,U��������Q�xz���˘�d1y/e�jf���	+.��+�UPR)�Dg}���3 Ln����mȜĸ0��7���+��K2m_�ܠ���Z������ F*���fS���B�Ln˨�������=�sɻJF}y��
��q��*�q��J{'SP�� V�,�8��{���!ƴ�gN6�=\,q�_ȓ�7>��H�-"l8��<�7|�lk�%�N@���-�6��J�۲A� А��ʊpFwM��2���C%Ǐ~!��|�t^Mx��ۦ�9�:^PKJR��x���4��&	rݗ(�`]*��Ba\�gg=Cu&��G%;�1{����%Q�#.��ڜ떴}���1]A��e�ْ��̻)�k�ʔ�?I{�
��k��[8�1��n�Gv�{1)��t���������
�h�yM�u����9L?D�sS�i�|�.`���}#���=���Ҋ&oԹ��/��F�;&d�����I!�����<c�� ��4�a���`��&����lX,�
���d4�}r���[�}ѝ���j@2��!:�|�ܿ��Q�0�1�w���x�`��5�]30u��ɼ����Z]��7+97�ns�����ˑ��ˤP����.=	�qv�UK����2XD���
�d��^��n5�ۍM�'Q>�D0�0mC�$\~˕F�(�h�y)(�OT�C,b��)���+]�q�$v�<�tL����Y�������f�vg�!�ݢ��ݓo�n&׳��G����|W��%	3�3<�&e����r�w�?�Ai@?�y�2��I��n�.|�F��Hr7>�)�!\�/��m������l�4�ƨ��O5����6�8���0�0���%ěSZʲ��=��I�L�2^u�YRR�WfCp��6����t�L*�cA7ի+<Ow����;�b8��(��a=��<@]���"�v���}XY!P���_?sg!p���e#�JC��r�˙��ӝ��x�Du$�+zL.U�UYR3��9X����9�;���\�WjD�+�X\~�Vn�(:ځv��&�F�٬c����J�fH��9�
j�X��g��w���⧆���308'�|�� b�5���"����v;��d�L�f��}��W�XO�������D�o��`�?�kl��ۍ"� O��$ K��Q^>�8^�, 6(� P�j�7صJu�=����� �g���P4x�����"X.���?j~�WE|\Ch|22�7��^�c�U�R�ܧ����_�{p*p��\�L%)`�&����;�~��%�.f���5rU0��+�0�����)Hjl�h(/t�S�5��!����ݔ���ċkg�͝H��#����r�W[��X=I��d����a�;��Rb~�i �u��ɁҦ���ڠ����.���}����Dr���~隉O��';�8�\��at�܁�8���߷��\%sc�[��Ƭ��8�9�k�6�]	�K��M��������MģCc	}���W04��0����,V{�5;��@w��m٠���_�y"�`7Vȅ�;�o,�}��p�=�u��Z��e�y	;�V3�$q�p�֝Ë�⧬.�/�>P�L
�8 b��a$��Q����k���=�=MQ}� hD%��&F�@��/��
��MM���~&YX��w���H�W�`Т���Ş���F��� '� ���8��G9O�'�8U���}���� ���v���)���Jʳs`�[���_z1��-q;{�{��Ω��t��8�#p��ӱT�i��$LO��/��]/��H0��ቲd8�"��(�K��6}�ʷ�xg$=�� �S�CN����!��$K�e����պ�,���^���������A�y��r�V�@��,���c