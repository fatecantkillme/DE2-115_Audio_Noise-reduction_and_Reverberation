��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|����z=+���v������P!��:%G:�FiC�T��zn��K7x��8������pR7�F�'2�L�=����X�m��88��!��DP�X�˴�ELQO��]���״ܶ�d�{�,N8	"����8\Հ��M�42nzm�D��ˌ��2�*I��j��{�̀�1�y��9f۟�
���*��*�P�˯�����ʎ�Xc�۽���h�'l;�=��#G����o��5|O2�����&.�>�5y	S��p�g�E���@�m.4�N`f�`��]a�g3�j�d!:3�I��� �[�����X��Q��K�ev�t{����|��LSԺ������<s�x"��2�*�P�����IMK�� ���Č�Y�քCɥ+;m̳������I2oZ���9�C"O;�L�hm���9�������aۼ�ao��ø��λ�!4-��^K��
�3hވ[� �D�F�@�U�6��^I}��$�Y�ˍd@� pDի:(��VR�K0��!��um]��_ֆ ��m,����+1�Z# �&ҙ�cƄ�`��=Kbo�x��o���\J�w��K���ޏ*jв�Z�'��� q1ܼJ��Q����N���@tR�㉋�#�����KQ�Pk�O�=;:k���ssθ���:�w���k5�*_Me���	�Q�5�睒�^����xS�U���#��*�%_���� �KtG�l5�6?�ߜ��\!�`�*�$5����^Hܣ�K&�w>�E�!`>Y@a�!M+�0'*�TZK<'�G2�S����KB���R�zla��w^�i���bN@�o�;4.�>�F���>|>w�m�$���l�f/��Yl�:�ƟC馬��5�����
Ҳ��;eJ|y9�#�C����QN���WtiI�·D�u��2Bd�,���8�-��j�GEaa��KzZ���Q׭��
>:��>��O��5�W���|��IYT��~}kKa�a{�{I�����l	c�I
\�aF�&�>���n{�Q<:c+��G�ȥ
Xw���<+�+l�ݚG��rV��]&ҳ���e3rW����W���Z�����Z��L~	��[��z�/߰����u�7��y�`�,L�3�Vk=$��-ψ���9��!b��%hHqȇ��R�����!��_7����? @�̢���y��8���\Ȋ�ys.IH5
h�|��r�'��ؒIZǰ�56�w<d6�ԾxB������3tK��,d�������G �A�T?N4�=���:A�|��10
A�"è`oQ�9�-x@���COD_Y�F�
�p������g�<��uXm��r�s^+٩���D���]Nm����y�Ƈ���T#-V������c�}�f�{�����:�S�Ǘ�q��3?[���Z�]��mʣA�,�1q�d�[��ܤ$D���B1a�t���������A�`wA�;�[wkg �۟��q��H"���.P�s1�����^o .�=�kl����鞮N��s������wL����O��e��>~����Z�)>r�c�Mk���x����9d����z�p�y�;Q_�b�6-Oqz� ����ǐ�fv���J#+�.�"0d�{�l��x[���Aݱ����t쵅y[���B�(���&�ۑ��C�޺�ӟ����|���]2���<L�b <Ē
/�ۺ���2��:@�4q���Nt��u ��s��M��uR�V�B��&��vA=��Da�~#�n��Lo�ֳl)��u�u�����t�#:��J���GS��J�M��ړ�5�����i�#�=@��=���jX� 1�z*��k�*4
��J�'�����?�o(?p�rK�	?_���E���q����<��H��v�H�d��HAa1鷷���|Nq�X����8	:�B��B����?�`7����X|\u�CB��ࣻ�����4�pɶ�̈��8*�ز\�!1���� �_�;gO�mz��F�)���`jB�ߤ��V��(��Fe�Ui�~`?jw��"��u�������xT[ŧ|�~�����4�\�0��6�1UVr�l1d#�[�q'S��F1�dt���nv�',��pK��p��M��`��gw���K�qG0ͺ�gl+�5�j����!w�y?��*����6�}͇k��F�a�G���?ک��/�]�~��E�gC0?q[�.b�|��2{����F؏v���򿝱��5�|{ZK��=
st)0_�w�}MQT�z�Uxsމ���yxu�yGK��j��#���V�����Dz��@pld�
��S�a�Ӕ0�6;�u�d|�XMn ��*�g!Jz��?jL����<��^�ǌ��.О��Ղ��q^4�jhE�
#�e!h �v>�"lz��͒@��xX���4��3��a>n�A����s�[�J�4ºy����1��i�^�YPĀ��<����|T�-C/A�ObxJ֟���q��͆'�h#J�I��k� �T�l�I�������lUz�A��A��u)SN�q���Q�JFO�B�����tG�\^U�P��	_�����?7�&I}���O��mp��) ��v�n��؋��RMnFq&�
$�o��Z���й��v�7�й��׳ӌ�P 7�{'l}�!I[��3f�h־�I����kˣܹ�X�w@���KI����ѧ}��|���] )H�9�����G�e�����
�S��Z��ᆔ��R1'.a1n��'���kkY3���L�}��T��U��x��6��03c�p<���w�9���:8R69)���D"����%ω�AcEΑU���^eb���;R�_�@ 4<gy��)�i���'���C=ď�h�.2�t�Rr��KOؚ�C�W#l¢��� Ʒ��k���,��{�[w$�����	\EVٹ��;L�H�@j	Yl���4��o��Ą�rh�Eh@E���g�v�*�������4;���g�<�{h'��)���k��]��v�~]�R�Y������^�ַ��-��L��N�ר��q?�z�py�5����hY�Ĩ�]�>פ!���B���(������Ag	3�u������T�3�� 5��}��$]�hY��7<��=�Òju�)�i´���<�~�� '$�Ay�u����$q���T�?��<9��*�fc��@*Lr�v�apR/u�LG���)�t�VX��}\�����iV�7�%�s7�0�bi��%�8�Rʽ8󲙷�{������e�i�xzD�~�����G���N��M�| ,}�ӹ�����L�+v��O7��T8��K=M�6��L��tұq��ă:�$�D�ً>x��ۤ�n̝�)	��]�:����k;�7�H�G�~��&K�f᪩�@���J�c=R8��!����"�L���j'Fi\���e�F�%wpu+�-~���&��x.9�׵�.�9���R�w�ސ`0ǝ��x댃�5H W�:�fA��p�\G�(��XG�gU��1���{b��.\Z`�@ܞ^j�$�'M�A��6ڸ�