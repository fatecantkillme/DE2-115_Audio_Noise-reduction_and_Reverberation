��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�8k�)9�k���J�f ۘEN�R��>�Ug:�&�1�X�,l�v�u�*U~��+��g9�4��e>ɾ�H6I*.��%������<֡uE!�A��`J_璈!������r0�6�"�X�!�R�p�"�`����a6�;�& Z>�=�$I{�Vdmn~��S�q�0�~�����.V��D�j[lهZ�@��Y�v�i��c�ke����8��AE����*ķ'��-����N�{�����_�z�}$�f�Ǿb$�s���!L}���j�4�:�z�áB#͍�x؃X�{f!���	���R%#&�<�N��w����ӂ��&����b ����+OGh۪Z�=���W|+VJS�L��,fh,�,���p�в~" fu�o?ei�l*�^����|�5�t��jq�2�bd& v=J�>�f��I7~�P��zVk��OoSwS59�0ά�8��v۾~C���7d��-��^�r�A��BV8�Ǵ����R�B����Y�o�T��W܈G(kk�j�`��f��B-e�銜q���u�X&
X��~�J2��mNc�AxS�$P@�"��P0��iM?�����6c�zZ1o���ذ��?DM�����&� ��b�i�m>L��7�CB����g���ړ,><��wE�#�7*�r9�f�q]��4_�оL䛳����{_�2I��`�̟��^x���r0�|/U�	�!p���nW�m��&~�a\9kZ C1�$��y�v��nތ걙�^Qv��h^���9���9:UP:h,S�d4J���N��B�#r��Ec@�T>�������B�_%����i.��{��Q�DAX���Α����3�� �ju�3��ӊ8�5����S�Z/,l�ik��#鈠�Y\Zm�vp�2��a�gH���O��$J���j�ڼ�Zv$)���7��i��p��L	l��?��wG��RPx�}�)s��=�w#���o�oM�S񡞽�'��)6��?2+�\��0Uvp �������ڷ/``?}��q�x�ez��~�k"�V1f
Me���?���.g@�Ďc�>N[֟계�p=>�U�'#���� ��2>�ߨRA��u2⿋���J�%}�U&jzӂ���$�H�/T�^��J�����Զ|�l�e��ɹ�|� h�^3@��w�]?� �R�
Ǯ���/\nT8�X���T5FW�sE���$G|4��)DZ��*���\͎�jn�=�{����O˛\���i���	��5�%|܎b"��R�t��u$	���K�fEX�P	�4��1s�I��;��e"��=&_�&��9�	`�;�Z��v�vڨ\���3c�n������s֭	���r�ś_*y.y���d���]�jQa6��=1W�EѦ<�x���.��([���p5�<v	>#d�7b�J�;�$/�e�u�_���/k�m�͏���Geі��e�~>#�׽(F,��w!��-�%��y��r�ك6�g�B������DΌ���2�u%�Id��ټ�u�|�N�Z?u���G>엣U�܉�S��"7�ث�S(̢��.��G{���N�	��^�щ�'}U=��X� �����M��M��+lꮩ�#.�q�D�F@�[~��:<�A�e��ЮE�t~���)��*g΂�}r��M-d3���B-���0��7t���s%xt�**o�:�@4�(����[Դ-�u��!j�9PIiQײ��������2=�<�������PX�(�.Fl�^q��ظɚ�C[�����=�$\�O�2M8��t��ʳ�K��5�_o��0�,��������"�ϲ��
9o|^k7�cMu5.��!I�CSbש�X㲍-�E�l1ü1�}/0�
=���S4
{cvX�7[��hk�����P} ;{��Q���j\l5��5�SD�<�%��������b��{.p�c9���R��!Tth,����2X ���<�-�+���
�X�J
�V�y���% GK������
,�˜O�:�4����r���s/v����}��$�4tKB-�����8�8�^�_��l^ ��{�n���XsĒ�m��M�s�x�*�"��0�!��YnZ�����YLϳ(}�x֮��W��aK� �{ӆ`w�^P��R���?�
?��֩�ph� Y���D`su�7��W�0	�z٦�g��vT�z}��a�Zw�����@�G�~c��&����]�,ת�P�K�(H�ŽM���jOu�h)&�]�~�=%z�G}+��'L�L�޴�	l����4�U��H�(���8�σm���:���O?�������9L;@z���E,qe�b�����L�K\a1�3ifs�5�����P`��y���'��5#&��[]���~Q@�1Ԣsy��3x=ˣ��@,r��$��A��L��qK���-�,��Ky� 9lk��O;:��Y�6Q�����:oL��d?�W!;y:؂d�CxDK{�y�u)Up�������������!��Kt_�C���HQ����l�z9�]Y�:~Y�Cg|Z�]�l�rK�^3-���9M?��Ō����F46ֆ1��X�e����������myЄ#'M~���l�B�YD���{@,���Q5��}zF��8��iF�!3���>H��W\:2����kz"��z�����3>�(��d�u���!	Wf���-�b�#\��_�X�I�W@Kv����N�>��$O5�YƥVZ����7�q�Ƙr1�`��4�x��fiYR]y���>O\����ɋy�;o�8&�[s���G��Tlɟ{�A$��7��+��u� ��W���S�[�E+�j�2��I� �P��#�ڰȫ��ī�y�J�μ5Y4lb�
Zq3[�7�~(R���[cw4P �*q�R�G��x�W�l���].4_!/����>����i7���C�+�
�uw�!��^+�{ֵn�;L"7�H5i�-��Q'��x �R(�;o�Ym�$���G���B�j�+�f�P0U��v�Z�xin���KW�tt��g����;�F������EE����<�0ׇ\� k5�[H.��ܱ�#��븴K_�\���eR6������fU:�1��)OP>,�z	Ϥ���,D	�j�1�]�9�k$�����l]�+���]�Z�י�5����Pm���;�r����l���
��:�,Q���R޽%�Y�bX��w� �"��hF�$��9v�>���n\�N��Q��Rǌ�=� �8Pm"�����R���:A=�6��1s������<yiF�{���Y�Ǽ��)���AzƝ�U��_��Q��bN�/>�h�f�T��Ƕ+�-�3+���� -7�R``W�%�P4�h�ĕ�K�ITG��dK�OzA��Ho���z;4��B�mE%��W��Y��[�!8Ƶ�P�޽X92�4a�vO��B�7��Դt�AQs�)��#]�cX���ԋ�W:�-WX�����oo	|�xR��%���P|�����]�EN�ۥ3s
M)ܠ��=�U � J�%��BG�`eA�'>?�Տa�	5�g�j`�K�T
=Cs$�2��9Q���\�5�(�/W�9U8��Ƴn<�;��fQlq�����2�Ao�m����7��
htiS�j��������0�L�Ԡ�$ERTt±�ĕ������@�C'�h���ɰ��
�<�����ͯ���I��F��2e��Z�	������L�y�ss��X��i��N����v��ߞF�NOM����x�.M{���zw>$8�m����6�_���^҂Е�Nϐ	^ffL��z~5�2��?S%�G���F?�q%@������N]�T�=�$�`~�O��K>Κ�K�!�m�����{��_�!k���r�	J(XR'T<����w�3N��n�(��z� ֶk�'� k����LX����	��tǆ�AR�_V#��r��PDP�)NDG��86q-cn��ma(��h�|W��am�smZC�j�rX�u����C�wR|���h�P=6�UXca_B?c�\-�m=�P$����!�ق`c����У���6N�� �:T��L�h���U�7�ϋlG��-��6L���\�a�S��Xw11��Q/��$���\^褟u>��i�^q���C�]���\9)<���=��k<��v�Ĵ����E�ޠ�+���a,��$�憐~@ٜR�����p�v��F�pF^#�]���=C���l=E�^�:���y#�o1�K�щt-%�$����+�3A�E�\H��ڭ�zo9I�5>�G�"�o6���ýۯ��$D�]˴�	�@������
\/o�m��Cx���Me���)t�������z-� 9+��u�����!�l��X'ū����F�Pp.��0*��ʎ�&�l|)���F��
�1�)��(�JZZ��PPd�7�D�l��1����ì�Q5�V9�ֹ7p-0��\��>�I��	�c�h��lC��_gJm�{�x�Ԭ1�(���"b�$�1�X2��T].A��f�Yu��l���>�Z�uʊ�0�O�R sz
�2gN��M�i��"�S�R]�4b�鑡��lAq^|w�J�E
JB"0�Q˜�z&K�'�v@!\�כ��B�Ik�2&����a<�l�C�%����o�=cGS��ɪrs��$=��N� ����H���2�u����)��&b�Wcc`����9���2+��V�R��f*��S�,�����������3�(��VduS�k`�,oJH��<h��r�?S�DC��ҕ�D��s+��T2���*��.��s���~��r\��R������Qb�L�uV)\h�9�D��1C$�m$�En�H��\3���&�Q�(���=R���3V���k�u>�<���fh�75�b�����#m�惭�g�q��b֞�����*��䘽Cm�_v�>��b���;��8Mt�<A>�00C�����"G������}�&�%}���٪:Z6إ^ ��A����l������e����?t��q�����>��	R(U�ڕ��2"���!���X�Vկ���}�m� ��b	-��4�׾�&�}�Ԕok۵�Tja2��O�em}�}��d�Ƕ�5�k�ؔ�,��Y�~O#SMw���c����]R6�����7.�2�w��	o��Φ������R ���F,~arI̽x���<͎wN-e�ض��΀}���rV|���~��Ί�G��n�?)� ��� �+cNb63�8q��ōi+�����X�lU$�5�ۘv�<i~��K'�y���*�:�R���"���,���8.x��˚�_T>�B�����q�x��q�Ʈ��i�l�1-�e`�T������Ԁ4yE�,N�ܨ�g�I��A��WЙ�e�>֮JK���8F�+�*:7���#[ȉ�oZR1A%]\mH2c]�;�\/�&���Z=�J����t$Nr��1�
wS\�@��\o�����-��m�8;1d����af[�P��{yg�*Nk�<(��ё��@�	��r��CS�ݽ��<�������BX���CԴ���@{��d#���O�:��來�����"����6��\'�$�Y������E)�'��;�'�\��a,��buqQE|�S�3���,~]��?{F*�Dj '���3b8΂H�uvε�k'�;��E(��R�qT`n+�7 Z�{aаTK�E�0��P�|ѣ����a�	,�hlgiq���/�k'u��c3�!��Ã�d"R~� h����v��S�T�g�%M5\�&���F��ކ��8�n@3�_G���*�c_�E�����5r�=�u�q�6�x��f�ܖ�5O�T{�I��6H�P�q���F)�1n�h�i*����X{�@1� �6�{��p��*{�5�u�Z}���c:E�x���ѕoL=Sd�d���XW<:3՝��[��r��'/�K���tY��y��<T�4�S�T<"
~��qA;���P���GƓB|���Fz�{Ė��/Q�5����'��Z`??�����Z�2_�r���Q*;=�Y �P6�NYrk��VLH>h����_�~���\q�Iso���_�F��g�SѴÝ�^ڈ*��ݮ�(!TG��I�ϝF�aNF���::\(U�.C_:�-�
=}+,�C�K�=��r`䒤���R�JP��d�d+�,sNI400M�r8o���������dy��l�jtӘ7'������[w^Xju�)v�yi�y��,��Tz4�e��ꃨ��Ҳ�]��0�� �%�v�c@��tB>3�eu��6upwGYl�}�)�E�U�Rh�y�5v�jA�i�2./IT�g`�;��5@^��E��?�����w;�&�֘IL�y�:��8M���.�'I@��e��]�f�g?��,�Rc���f�a���ՐS�J�Ak����le>3b����=�w?���;����	_=k�[�/���W�1��
G	غWjw��"��V�|����;�Fht=XY����ӬX�!c��	��+�tr�u�e���p\�N<\w��F�+�j��r���H�8�9k~���$��H)d���X��s���AR?�|E��{ӝ5υ�0:���˾�׺ ������RS02�kqJt���t�8��[�q-�oZea=:R�Yx�y?ɗF`B�H���)F���5�46�yqb�ɯ�h��~B���.[�ў[�D:S��X�ݛ��s5�^[(�H���{pޥ�����.:&�3fa�����R����"Ԯ����`���șwZ�҆lp���j^j6y�l��Z�����t�C��#��O��Uf����E�`H��H�#ǘҪ��i�	�DuG��Q�Dd���%ă0��
�+�>Ґŧ�XMgwš2&�"��Y���L-8��1J��
�ׅ�P-�Ҳ��} �Gm�Y
C��uƎ�,�����b�>����7%��<2uj��YȐ& ����@�œ&�G�e�RWc�{Jݣ2���~�����t�d��_���Ud��_|�G�]7��G�+B@DvR�h;$�_v&������FPc| �B�T�Z�4R���!\�~n�1ϋ<��#g��л�"7�)��n���c(�Yc?��T-}���i���)�C�S�m�9H��[�CY�\�JS�+��y�~@�!�P�H���epI�[~!&jȸQ�EQ'�0�n/��'-���%�