��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<S��!O �&�>z�ْT8�m��mC�4�N�}z�C�q���lΚ��օ�#�I�Dje�S�)���������V�g�m)#a�����Ђdb�e��O��
��uc=å��x��g��$Ѫ���c#;3n	d'~��;W[;�!�]/bO����VX�i�]��^�����x���B���~G;\��l1��g�[R�RgnyK�pK�"W��OXs Emӌo�	K��Ck�u>7��t���E'�R&_�=�(��Z�"�%9v"UdԵA�7cm��xk֘�D�'�d�S/q=�lo�̑u*�b���뗢ިn��;���&~�(.�/�U)B�~p��^	�5�}�Ɏ�)�Ճ�$�a�y�pOJH��wbL�E�m������g���A�F�p�����aAEV��dbl���Ǵ�����s��Y<!T��j��[�p?�j���3�q�Y����z�q�hvYu��/	o�z>�ם����
���h�=ʽ�7m���l�(�=J��ʎ���q��«����\��&�.$`��,�ʄt'x	W`���0����h}Qr�
��5�,�
^�������j���{��#IĤϿ_������Yu82���a�>3}'պ�cȘ�꩙��o~t�[��iݯ������!/�
m���ZE�t�t�����+e"߄����Ŭ.<��̋�&�m8��S,+��Ap!]���p�89�K�Bi�gNG�?u'���Uf�̒_?��*���AF{��+7'{�J�,į��t&���;}8��{�?��(���Ɓ�,���g_�����gp	�g��`Ћ':N�����FO���(�r���N�cE�s�.�A)��Eo��MmS�׏����Y�˷�74e�x�שּ<�9��l#�{`[�b\+�蠱�f�,����9f���H]���*S�l��q�J��?6\��L�t{�@�pF*�2�'9>x�@��8�IhֱS���!�Ք�_I��ͨ�� ��f��j���Ƕ�dO���Ov��Ҡ�ߕ�E�����\�Nz�E�q��ɗ:���'��\"߭�N�V�z��5�"��7X� ��߻�s�!u���u��F�����ᓗeY������J���;��qz~1��{Yb[]��`T2}�DWyċ�.��e��,�{]l�%���1�R���`�V䡎0�*J/�Q���U���tӿ ���.z��_Mݣ��=1�ي�'+k?���jƜ۬KO�{&*�dcaY�A-���\�/�*�1#�y�	W9Z�{��4r=�0{��,9��Ed���&rD"Grx5nI����X-�I��D��"��چy�̓9乥�V�&SÖ������uƄ���,�S��E#��W��`�\��%�|{�ss���N6���7tzR���u�ԅ��D)���Q�7y!�*����ܦ�7c`�� @�\#TwC��:'M4�qx�[��x��h�B�� z�B@`�[6�N����zt��SWε8����b,�F�Ϻ\)�?mM��M�-_!�<p��v���D&V=G��m��=�xB��e����3n#NS:� ��c&t	}��^��=E���uKx1���na� �M;Yt� (�_��b���}��.N;���H�ΥW���H�m��ކ�f&��&&6x�Ҷ~�l��'tQtK#�bE�����&�N���l"yg�7j�t �<��r��O7b����!��.�NW��$�(���hQŻv�0V��yԦ4E=�Ho�b���:'�#�ݝ�����]��I;���w
��W���P��N�Q	�sW��`����3�������hڈ�ޮg�	Vߊ*���E|}��V�R����]��s0�RQ�!ΐ����C}��َ�OO*��#ޫ���+�%-TX����-)�6����D�D��#=�K+#ש�cT���1+�T���c�ȍY��r')!?i��Pb(	i��`A���+���b�⼾"q��7/�H�~�{�U���kO�F��郛�9�Ҫ��b��k�Z��S��^���Aom~l�I*d���m���6�m� tt*i��j�A>��F�qx[�i��}be�CR�m'םċ[<��F�����5���x�L����r��]@��f��$��A��)�&���-���?_�6Iz�S��Wi�G�E�}aP� ����PzF�v<}�}�yRz&�iұ�b1�Sij�u�`�郹�g��2�,*����Qß� r\O�s9�Vø��H8�����D�ߣ���?Q��T����p���3�Wi^L����٭�z��٦�q!�[��dM݉HGqLt�L���ν#:�tQ=�->f8Ѱj�DC6�I�X�eguI�������٧�r�
v��8�Ҫ�D\A2�J6���zP~=ۘH��{;�ONE�Ҕ��T�u�5��0E�Օ�k�$�59o>��
kS��~n��G۟�hu��AJ�GX�J�v�������[�����'�>�]���4����3=p�lv��%���a���ٶ�;�kW��ɗHD���C�Y��4eR�I�֪�o*V��W�A��}^Y�I���e����Z��&�f�S�Q�xh�������2}g�O��L�;p9/�8�8�A�2�����J�9�7R�/�u@�s���(S���}�:ODiq�Ȏ��ځ�/�al�.�В���@\7���Ő8��	V��p����|0���V`�BW��jt{s�0Hr����g^�CU\ǐ�/�z0&�����Goz�zz'$@i̐��X��m��nI�/�b�T"�(n�W��Ufݦ^9�s8W�����m�+o	R���t�)9`��5S��y!&����o,�Fή��V�;����~&Ƙ*�',Qn�a@��;qç%�IC�>5=Y�����)4�U*�{2-��6�e����L�[�2�7���/�8B���A�|v���ߝ�,��UX�Q�"�Y�bNc�j�`�NY�)���0K�+�v �!f�����^R�l�-J!��B��krk>Mj��EB�kwx�~S=�) �.��8id��S�sf��i�����"t 4! j&��.d߲]�?�F|��yY��Y{KC󗰼D�H^��M��D��x�)�i����b�g��2$�4��|lw�{���{�k8�����5{qm��-����?)!�$�i����d�2�M����b�^�D�,�9��Uߓ���X��v�Mǫu6~�3ÓnҪc����3͡�ڼ)���>y��K�ڿ�]��L'A��Ś���B��30`��La����^���r�SD�!���[q�C�M꿳 Ɯz�&1�^(<�K1�A�<#l}�̃�`���x�2���l5�j����%k5��G�X<���>A�������d�`��ɓ~ȵ��� �o� ���[�b���-�؇:N:�b��S# �i��
�Fc��]I�3�?�>�G{ܥ���X��1�p.��Z��bHixx��:��]�XMt����@w��0���p@��~%!;%�f�!"t:Ε���e��
����m�,;�Bm֬���n5�� D��(΁�����(S��A"3�����su�W��L�lK�kf� ���D�[��E��9�VЖt���ë)>��D~w���ryη��SKТO��@��|-����X����޽�Z��]�4H~O�{,j���������9��M�k%`\��p̸JOъCx�$k��T.tkO�Z>�k��rn�*�a��I6T}\�YB�'F=�Wba�@�p]W�����4�]����h��P���h��G�򋴫z$�4�fH6��
>	��s�)iU����/�F���4�O-�6��i�vuCS�pe�q�g8͝�|�,����؝�V���&�H���2۞���EI�4q��M#��.M�����''��Q�)ǲ!�߄P*�4�r�o��Ā?����߇����^�'�{���T��A�_m$z ��.muq�}��@�C��xB��Gk��ZX��ɕ�7�d��i�ED&�E�Ժ�
.�hK�Xz�a��ڠzI�y?�	��u47�z1EV�������90�d�S^>�P];Bcf�������J��9��p!��&0>�;�D�p�9=K���c��cx	��h����Ҋ������o+7�\��b#�����7���k�½�%��!�I�a����d�ٺ�E��꯼�@Y����Pm��<-b�|#:�̍��]b���X��1��}S��GE����ə�Z"��/$j0���E"x�w�jd��v�"N��LG�!���|Ssa ��cQ�V���)��D� AON��`��>pXbS^��6�7�T�Xc�ܹٓ)��=��|'xg�!���Q?ᩀ��u�~��|i5�`V\� �qN������x��ظ�jrP�rKZ��U����<��Pՠ�O��36��L�:9���F��PM����KS��\����~��_�(��O�|'G���O�t�I'g�;jbL�,�hӊ(5	 ��e��%=I�[�<�
�5�7�� jQ�r)0��0��
��%�#y5��x\�Ƀq����cKA�,��㧲��ȃj&�I�@W�N��������Ԕ�Uݥk;�<��JN(`�}d@/D����*�Ηң
ZڊQ�V��qLe4�e���_XI�8�3{1��I5W<�¢�=���s-�io��;�8�m���W��_Գ�MG�u��J|E���ӯwQ�dD�ٽ�b�L�j8�Yf�K�
����#% �5o֊���^��	�~M�ߺ-��Uqg.?����2��U܍���-_>��[�-gm@1��_N@L�T F��϶*��P��iRV+��%MD�F�C[���Y%[Z�%��Γhe�ң�y_DW���,��B}�gXz�53�S�σn+���z'�C!s�rF��آ�S�\�1� �=�癳�p�N2�$�_0V }�θ�|�E�A��^���r���ĶZ�U�Q�z.| �B�L{�G_��q�5����-��FU��X}8L����S�(�WB��H����e�C���~�Y��u
�o�l���Fx�,L��G4��J��1?��%�Z+t����OI+��:l"'D��:���g-� ���p��ZO�0�~Il4�yD1-
(q�Cz��"�t�'`�O{(Kl:?���q�Ǯ�����V_FFY;�ki�G�VKUX>ey��P��3�O�3�4a��s-�ey¹F�a�]c���\]��L���@����^x�MJW8Z��A/9{�qk����M�7P�С�+޻0J��|N�FRm��EKr�z���S^Q4ߢ�ip ����]��'p�d8`�7�8�3���tU����;$�ZL�C�@�m�GG1����7���0���aR�L����[2a�z�D��s�W�a&$���*c"�H,�se��Dجu���}�U��%��g������"�;l�ھ>�������a�7�4��D��y����M�A<�CG���6�Z�W��)9�\��b���q��ו���D���1�<��y8��5D��?��q�N��XNt���v�Lv�nGzjl�K�#�3�K'w2��SK`���*�H�=�)[k]�Y�b���j��B�F�����z{�cu�y�_��
�O*�_�ߡ`�?�#L�d�uhIQ��B�A�ܮW���΄��p���ksK������_c�"/9�4�M��5����o7H��hgф���[j�3��������F�C�H�{Eq�ں�L�{:�Kű �]�����g@::q*R�ZȲ	�Ph���mFF?��ߐ4�	*���aպY7c�����(o��|�u��@k�qx�n� �4�}�)���_�~�n�%����w?��p%�,��>�����<g�O� ��;ı�#*NRSxh�j�=U�Z*(Q.���]���b�F�6�s[��8K_&6���.�"t�du�.����ɆJ�)��������ȅ^��tR�F~s�<����x�tS�������?(��c2E��7��
󔴮g9\m��	��f���Ⱥ$.����2��zT�C.�hh�5,$Y~�v*w%)�͊�0Õh��Kɬ�%�:��!�F��1a�T7�iͷL��������?b����C~����T�����ln&�n㶞��H�ǧ�x���]hz�gL�ș�yϽ��Wo�O�w=�������̣z^��m��E� �Z�� ���b˛��hx/J����E@�ʩ=5ZfG1�4�P�mx��ebل�ejS��L��F���:��r���ízZ�q�+I��4n��c=NS\�)�.���voB�T�Խ�z��h���*{yv��R\����p�Y���
�xJ����7�~�p.��6)��c������=.WѮm��˭�0Zܜ���V*~�?-�*�O�:��-���`���E��+w[d�����>X�	�:N��͚0S�ϙpW�#�ܻ���@j_I��c8��Bb�(l�[��<� ��]����O<�S��[쾔:`}/k�6T�6��nns��
)Z��x'm��vR��es��P?v��T(|�g;�F��w��9�M�7�,uh�������n��@ʟ���9�`$;���[Nckd',V�q��S�%�9�W�
Z��{ٴXZ~$�Gx!�z[m��A67�ւUde�!�3&~�!2��@o1���6�~G���2�����3�=,�Ց版�]*[�u+�:��� ӄd{��'��
TC�ы4�M�����K�g"VaX����l�h�(&!F�:ak�wL���NE����#�#ѽ�(�ccV��	]3��f��<�F9Wx� �	vY���A�6{�<��R��w��DB�ģ[�,q G�6��cβ�7�rԐp�܎�$niӋK��X�bGS���P\���} E�J����%�����٥z��I��t+,�v�j�����4�d��[+�Hȅ	Mh!�I��� �TTū'9%{���W��`E�DJ��X݀/4�ۤQC�Q��/x�4*����2#9Eؔ-_4�!p<�&;�t�1t����d �=݀�N8��3��M�~�oc�!\1�̋�dR~��0:1�1iP�����+�I��lϊ��Oi�T��Ji���]m�&9#��ـ6&6d�&��׈٠:N������8�S�mk4��-UR`�cYW���r )���G�.�_m�=o���*�)*1�~��>�v(Б����#��F��u���)9Z�H�̦}df܉$�/En;9߼F��M���>??��j�UN��e�T�.>EU^��ؙ�嬎��߮bu�d���:��L��ؤ� [� �RI�A��#��d��{|��`H+���H�>�N��`F�t3l�:!�;D 	H����>JdƬ|�c֥�{y�He�A;ھ/6��p�^웱]��eq�*;�a����8�W�B�8�.�X$�J��{�`P����Yw��4�=
6�4jL��+�$�<���"m�����8�jB���u�T�ҞPH�P����AՌ�D�N"��b���A��V��ڹ�m�s���<�*��L{�<S�H�cI��,�����I�îak�𦓐5�!+V�`�R������z��Y�M������x4��h;�ӛ�R��S��L,V���ı�Z�4Pk)�d��XR���F��#��1y�;��!«�p���Lv�u�LV��L�&*q�s��O?����q$�3��T�M�����q�>��4�8Ag����#
F�]��Ŗ����_~X��<BͨU�\��W�����X������S����O{#���H�a�'.���s����{�����Px���s��y��)�>!a6n�}#��\!�>�>>��������e-7��I�� |���V��6����	����l�K�[����j�`^O��� X{�c����}cH�G�����0���y��`s>t�"�����(0����'A��Y���w��@Ͷ���������t;������aD��Z\�_�`��*���{��$��jU���EK��|7�����[®�c	�d�U�׿j��hW���	�)��;6u�w3!4�b�K�Q��x�:b�^c����
�K��X"�]� �Ky0e���ݗ���1ZZ�Бd�=�B�2 k�i0�5�y�鑪�3kҩ����M��hZB�rn�a+]Y �,���d��1�茍0M���k�ȸwE�`"��z�_ɚ$�!~ 	��h��0%58��1	%����;�c�i�۬�s&.�;��VI=1�)�q}��E~5�*["�c�X~�v��40Tn�7�rD	I�(�Ύ��or�7��+��
_�>I�O���78q#nC��4-��ӈB�w��6`cm$x&e�����R�u�/�LX7b��,L���ل�0��A��I��[�lځô���I0���7���F���wv��7j�ڮZ�1gT��}z���M�lW"�2��j��n
���ׄ�B������,�	0L�d�tQh;c�Ǻ���"!�MAd�;�ԇU1�8T�������Vz�#������֜p���W��Zx���z���?v�p�1-�]\V�u�N�A�Ab�4�H�μ�x�:~-R+�_��f��_��
�	)�� ;�� ���Ւ�L�sI\���ZBH?�{e%��6~���� I�($�줈��<<ZGP�v��OɌ204ZlD�oƷ~h�����Q��kv�l�%%E�fpK3ȿ�o�}r �p��M�ٵ��UwR�tX�>�- ���DA�u͌�EO�.3��(�t���Ɇ?����t�q�V�_��q��_6nD�G��<����7���ن3�5�Rv� �����#��j���b������*�;���%n��o[.��A[��.$�j���a�okKaI��ȵM���D|[�k�� u0���[�:��E�Yĳ����s:�$O	oj�lΝ�ϣ�]�e��w�,J��홀�f�n�-m
�j����;�<:��qj��S�
��\Tl׼6p�pcȸ��6������ڶ�jxhM\g��ܓ��e����-Eҡ;���˯��%u K������c��T`��:����8������i{�����J��P�8�k{v��c���̗y��,���W�s��Y��y� �A������7{.}�O,���oz�W�}�%	�;���)�s�[8#,T�Nqo���@�?�9
�-+�b��!B4�Il}�	 X�ń����y6��R�&���b���<�T�c��+Q��U�d�je;7�7�W��`���} #^S�t^0�r�^�艒h���%J����57 �#r���6ָ<���{�
�`IpC�Dx�>T�����vA�=���r&�T�(-� ڌP3K���+�﫫uH��v���Raz
�tb�@��Q����*[�����~�H�<�Dz�፬޷}�@�\_Y��Pꟊ|�	u����a�'�XB�+�|<2���C���R.3��W���}_�2h��\��ژ�M1�i7����A��W'�7�uo�E$�Mw<%�J7� �%�����3��k�5�yu�D�dΪ�m�y �7Vqs�z���Y�ODT݇:�G���,r�{e��A���礼�։7<Ji�/�2Uރjt+et,̽;�Q��'��`��*�;3��181r#g�B�E2�v
���>et� L�F�H ǿG���r��<D;��|D���c�C����2x�]⨇�e���gw�|������vW�{Q�ZfR��~m�
b��?�I��b��ĝ�A�Č}�Z`�*��I#�Q�XQ �/�4�[�c��u�R��V6���*�l�u�߻@�����w$���2�k�ͻ�Պ��@�|V/[Ri�������twB�4�(Y��SK?����@1�������5-��6�\������t:�HJ�ȷ�e�]Q.�����B�����Y�'e���K�r�%�pșm/����/i]���9�l���R���1H�@t'�d��g��xd�8qs�[�w�s�C�i60���P-n��!de�צuC���G�b�X5��b�ݷ�d���b3l���N���1��<���
���ܒ�V�������ؿw�p�RF��M�"%���:����b��}�cاG�+�ʸ�
����o�o�v�=�B�5�S"�Ƹ��6��%Ѝ���[���'�ູ�yF�Tp�[�)�������y&����}�fD���`�P���Az���}�0�:a�a�э|b�O����מ�\�V�Dr�a�79;�i�F�Q�)�U�����������:aF�����ToV���Zd�a����^]%��6xc����%Y����o��^�(B
/gsk��eKaQQ�>z�����~�_�EX��A%�&Sʃ�m��q���(���o�W�BK� �[�U��敊΅�[N���l��P8��r��TZ d:���/, ��q{��lK�T�|	7ap�u2�1�T:P��,o+�����~TK#h�C�C0f�[L�vIs���'٫:3� ��Uc� �Ym�X8��T<M:�]��_H[�-�S���1/*��3�,��Ƶ(�xj�Xf�|��� wTR�������6}9�;���:�//��� +X/!�^=<��'NS֐Av��K>�4�0?JQ���tZ(P�gҾ�MF���U�����koBb��c��tm�cJ��=���i���8�G�+��	p�wV�׫^ǌ�Mę���׹����9�a�bB��t����Hƨ{@-]��Wê|G\'2$�`��*�����^g�~�u>���*T�C���a�);���`�n��6�{6��G�~+czS��U#����g;����X�Z����l'ING����uY�xAwF?O��W
�:��w>0b8	lGi�Q�U&�x!�;�)�Ӝ��]
Y��;���<~����:�����
���	n9�MD��9RK �w����oO2�:r&wt"̥c��R����*,~�����]_3ҢB�K���|�~��l*t�U�뿔�糷������1�)�Ҹj ��H�r����4�n��L{]�Ѳ�������o[�.̨���7��N�;L�>G[k�x��a��&�|Q�&�I�C�A��$-�c��&	R�J��؊��Ղ��F���dö90ʚ�c��埡�=�U�f�j�<��O��Fsp�`�p�j^.����dR��s�̧�Ν�}Yϰ<�����.pa_�
�k(��}u�`�Fy�M@��tw����I��]8�Q��XU���ll��}�HvIPom俒���ydp1�~�1B�+�d��w�
��������#��A��Þ���$�/_�FKǗ��6N�z�D���t8��k�)����.X���n�F��,�Եv������Dǲ��
L�l�3�u�QU"�ZU����"�� �S�Ma�eո��k�T��;l8��n�-}0C�vlg�uY��ǖ��&z���Z
��O��&c4@�A�1�U~:��(Mg�
�щ�P��=n����ųn7n�2����VV�ݙ�_��c:}�N�YhH�)W'yp�?��8��q��_��{�t�����m�q��H͑:�<��{g�0O��V�����{.�x6�B���mg�����{C����4���\�t��ўz2��b-$�&��*�tAR�|ʋ8G�Ū�n��aH���n�G
�JU���j@���%)����ŃVp�Jӗ{����s�u���C`G��כh��r<ADG�}ލ*$N&�6`�q�|yO�.��B�5��I�2Ɖ���y�Ȫ�Ց�>�c��;���i/�گ�Me!�޻��W���$Υ
�[�l��zc��f%�_=�R��5I���(������S�l��]S�j ^������#׍F��߉̩7F�a���~҂O�pJ��ռ���k첱ԧ��������@aL�)
�I�����xr�k��ø�Ui>��ѩ+�^�׀Q���Q`q��B@�Ѕ�:�A�(3L���(��֩ӥ�%(����Bx���F}]�|�,���'����M���k4�E�"(�$�{��_a��&T��?r��0�B"M6�&��.�x15��:s�{] "pNp.��`�/�J/�s�~ob���c��WP{���܅0�	R��)���A"�ma�[
�[��Sr��P^S�.T� ���=�M>��m/Rd�V˘3���_f��J�=�E��P�ͳ@��˺h܁��Ia��U�ۼ�sL��b_}:½Ok
/F"��ì��/��=�\E`�%�`��0�d�\'�bǎUkwHVmK-��:,��~���SE�H��n:i�y�P�Կu&��%E�n��.#kl��(���u-[���|W�۪�k	��Nr;ʓ���%>�~N���)l�T���})�u���0C�5�/u?ńf�%�N70�ם9�oL{�Z~mM�1�y���p�ul)�Ѿ���
ŀ��jx�eK�����x���>�:f���oQq{3mg(f��:�P�T�٨g��%�n	z�6z�����xo/"�Fy�|�"�%ް=5�l|]�?u��6i�F�X��FC����-β���C̩S��|:���	�nK��a�J&�X�7C9�aAۊ��{�>�������=R�J�`��Xм!��uĦ޳9]q�.�1���T%��1�]xw�s� ����'P�g�F��?4��}�[ӷ�_�j��'�4im�{8{�\B�5��X�X��^f}7��a��9�6ۖ����qt��,B3/^��(�<�nW뭟"#�zB�͂3�Y�Ӌ7���!����!��w�O�h�K>���w�Lb0<QSƐ+ R$��ƚ;)H�
A��Ȣ�~���N�l?9Ing�	���F�Xtd;�F͓3Y4��)��e�?�������6��#i����(�A�R#H6�B�3��л�=Y0P!��K^�M*�"� �6mƕIzF�|��%;䮺�-��G2*�w�L:�
�L��oVAj�W/��1�Gf�������MȳuN��ͳ��h�������&]��iRY��	���i�go����|�0����<:1�����D��^���D�^��q���R�~��#��Y\���,G�L����jv�H���&���sE�׉��@i�g�Nu����<�˓ֹ0��0�){�(�z;�q����g���w+��F�V��J#�i� ����8̅N�$jR��֩��Ɓ�W��v�yINߞ���]=o0ՅR�ɦh���MHp���Z�"�4��Ƌ��o�#��ڜ���������4���k`P����_���Ҧϯ��w�	��*@�/��jE�1{��xG��e2�A$����=��/t��%2<w'�D"J�v���v����uЄDE���R�&��Ť����"��U���bE���SLs4j-��a����4�8�8�����w��鍔��������q��H���d7���z7�|n���s#��>��L�<l�b��\}x
�3�9qL���(9�Ǐ�* M��m$���
�C��ʁ�p}�������J8���w����!ʬ��~��G�Y3[q/#�m��<����Z�K�KXU[W�!lU��g�6FrQ�[G���t��iI�w�L�<(V����RI�lM;E���f��k"W���/�xP�c��c�]����z��	$�����y?N�&���_w���$䣪�=m�9����&e���)���K_��.l�1�)���/��_7�/����bN�N��ڀ&7D0�|M�aC�3�ߎ��Mۻ��eȀ0"�G�pDq5�P�}������Cl�ȧ~b�J�WR��>$�6�K�|���a
����!g���"�1{����BY�#�t�l	6[�H�9�u�k r8�1�Dwg)��0�$F�ݤ�$G��A��qe���nf��xX/Y��OS���o�H�]RI��<��q:���� ����V�� e�u���UHWP�n) �fc�Ůp1N�M��rOT��v��"�/�⢘��ém5�4Fl���p!�S#�z'�iy㙄B'H�6�Ҡ@�Ң��K�XX�È'_��x�C>���s���������|9�:o�0pjA'Xi���b�$5�{�.�6'@g	�)�*�Ήm�(�V��}h&% v�La��+�&��P�h	�����o����#�^kA]�Mų�b%��Z�4b���xA4�*{d3.C���n�;�Ek��E������ۅh��>��8�] �c�=럪ةIh��^�sJ+�����º��[�l�Ys]��?��4?��d�4�l�ya�A�dQ�F`�����E& �A����]���-	��Q�'D!P�n�Źm%_��?�d������ �nJ�vȝ��Y��C�צ��`v`l^_����01��=@���&�%��6v2��f6��l<=-WD����\>c�w*�6mr�҆�����܊�z��wp 0��~F��.�:�H+h������\�����3Π&<Vk�9��X�c�@��N�[v�6�C�B���9gm����b�����Q�����w�\�J�[
����9�]c�rLl�����v/L���͇�|���J��j�[=��ۦ�p
F�6�IP�<rqLtL_X�|[B/�^��Bʠ�'�| �#1��n'�]��j ��̃�5M�e��[��D�X,_�;���ba�ԟ�ᗖ�ǳ>�	�0��U����%˳'7F�[�����R�i��0�	.aӀ�]�m�Vp�@�];�HM�WU�'oN}K�[�{~�n��=��)'��Y���Cl�Q��%x�}.BP� O�yp�8�֜k�w9fB��{��^R���z��]��C�(e�:4c� ��5�|��HвA�H�m9�i`�2B�~�,��k1_5�4`C��]��8#�
!�ߞu�Z�$P��T0eyNʔf�LW��``�?�����_�f�~]ARa��^���T26u1e��v�n��Z�Cya
�@_���a�\Ь���KY������CD��|����%&5�"��W�������c�yۆo��LL?�	��g1�R�K2��I �[
�E;���ƥ��6j/�[��
�7��_�>�Cy�3i��7�mK͗Q��tՈ����Sn��sq�M��ZjK�Ah��U���������Ns��v���kq4_U�\��L�GwT�h����9��x�\%e���=f��p%��B����JQ��d�n��I:{li\���)��$���I�<x�*O�a$�ж����Og���+�mB�,��L6�)	�\�;�Ķ����H`�n�"�A a��KY������{�w�ehS�'PA��R��{qcGN��/���*㳇5�O�n�h�f��m�����������BH�$i��@#T��J#��������.���C�W+^5����9�E},�y�*�k�e妡d���0�*�"&E2=��m *�J�vF��_�҅l��C��E������������H����{�g�_�g��+ѷA�C�!+��f�����m��LM'(\��f4���I(q��[jN�=ㇼ?�m ��c���H-˷8k�Q!�����R���!��{�{]���@̽���y��I�F<S1� ��am����̎�g����������H���¶��/�ճ4n��M����K�|��@�Zu�div�ļ���0��Ր]�����`c�).(��54l��O��e:#!I���y������Y�I�@���gP�H�W��|��	�z7�JCk�JY�N�d�*͢Eǔ�Y˴�ҭ���d�U�6���"��a�Ak���>:�RU)���Ko�җk��^��Ոyv���7ߡ7J��5���Z�q�Wв���i	��]n>)��D�h�f���E߾<�z�a��>c6��\�&�m� �Е\BA��W�����[4��ls��W�Y^�x?Jb~wU����H��)J���
>D�� 2	UO9�yX�?��P�b}b<!��p��3,>�&�E�|�d�{��ۋ7��
�SX��av,�l�$��[��pǶg�uY��e�*N,�p�6�u`-�dփ@|��9]P�F<bPRٳ19�ǔ�I�p��61p	,��"�jQ�J����h��O0�7j^f��_V�B��5�ҟ�_tp���6}_p�5���Ĭ4�����8i�����ꮸ�`�[�(�u��/Ǚ\pB�ò����1��Ӿ�;�	ؖ�w&��kO{�j�FXA��L�H������9b8ބ��@�!z&`.�OE�s�.~�2��YO�8#�Î��I<��$4�.WvT�.x;��Y����1/"3ow�!���nt,��EE�n}�je�'+��\mD��s��(A�-�3/��K��3�aE�OA��hX&�������P������,1bF8ҵ���L	��:�����ysƓ��Y��Sלu�q��9��Ƥ����.(�f��>H[
��Ɂ�7d3�;i��:��=8��lY���/|"�l�������z�$�u��񍋊�{�>>n�]���,�>o+?S�
T5��5���)�+Q�������\r����+�]��'[�8�^���\���(�`��D��{C@�"�����<z�?=I��E�l�K���Me7��n��`*	�.��D�9g���p��]<�r0�OA��G��YHqY:�"�;ɹ����3\����֚V�I;��V��T��M�1�x�e<��+o�bE�Cb�bG��r�t
3ڦ�2���c4�e�Q���Y7�~�p�S�`[1q��
��}n�%�-�����1��N8�JQ���H���� �7g���Z�M��X�E`��G���
[M.h<B�S|��?�[��2)l�W	]����L�\E0������F@Ίhb���]�Gyq�WH	��y ��2�w�})Z�6{��>�HLM��s5�L�4�M[��dW��C(�Yϵ q���]�]d�TN4/�Yv�s�O㟳���N �ڦ�Dձ
�����ӜR:"�k�sQ]����$��;�W �� �i!��/ʇw_�%�g�ح�S���H��.b=B�m7昬� Ⳑ��j�i��Qgh2Jie�#
r�]a�@�Q%���#�ݶ i�*t�,z�(���ut�&�J���03��_p簸M߆w�� ���h���{▴T��''�0���јx�71J�ޙ�DO��<�Qx)y"����Q�[�o�]7�{HA�����g{b�z���=���w��hi�1�]a�{�o�Ax�n�R��k���O6��}.#C~�"oҒ�1�0��ܥye�J�yt����	.��!���>��7?�wvs�o%�6,�4��s������L�u��Ͳ��+%�$�x9<�-��F�Ǉ[��g�d���SgZvňFgĕ�p7� �*ըݔ�c�Z�����\$�WS��u�Ji&��G�)$a�8u~	һz��m��.m[m�:�p�{"r���/3�v���ǩ����l]�S�Z?v#���-�H7&����k9�^�aFa��I@N��F!�Үc��m#�^�f����s\���I�e�sXF,N}y��!�r�뒋�辖c4�	"r5���ɽ42�ȃG�:�V�����pdp?��q]�?������t�&�9��s���.�W:�c|���ĹI(�gI�J�{1���v^F4���B�_G=�Q	\a�KF!��@��M���>3�=X��a҅02Vx�x�����G��NJi��Yy���Pa��u��jvUR��;��\hB%�c������Ë�9�_���?d������y�k>9cX������H���-'���z����1U}�	�)26 O4�ء�r+4o�^��9�)?���ɳ{��CC ���<U�	9������k�����?�l`$u04b�Y�K/t� �D�7<3�Q�	���fu5�e�Ŀ�z��K�'��ϧ�Ԧk�{)c"$(��g[���r��v"�������R҉cO�@���I`KA�/���f3G�|G僙����}�-��ٻW��H���?Da;��~e٠�Qٕ�\�(�씜 ���V%l�Y`��9��zzدKO�-v��[/�'���`�(Y����[� ����Pzj���$�@���u�qV�m_�jN��?q~)�r��>\{Y��A>�	O��FJ5��?�{6��%d)�|aHO.L����T���J�،�A7�)e��^��TV��qi���,rDs�	�PW�W;Һ�(1�L+�ws�+^�4.�+-���X\�^�bs����َ2��IQ�PD�=�.aht��Z��5y�H�*��յ��s�%/� ����b*j=N��k��W��%>�i�D+�j�KW,=�
,т�?�־d>;~>�7B�d�a%fV�V�g (/:$���Y��@Z�Y�Ҕ�͊t�(]İ�>K��6�'��(��Ẻo������0u�Y�	@��{]��Z�-�e���V�o��ͱ�k=?�������>3$���A:J�%���b�λ���?�I�
 �h�� S����nŇZ`vTk}��F���U~3b�+�4y-Ac��t�K�B�/{�D"� ����R�Q�e�I��s��1`�0Bj���T���{IH��-�K��iȂ`�zN�+?O�� �o�S��Ց�dJK��C/g��Og����]2�h0rX;(k>ShL�3���=s��0J�Q�FMZ�ô.$:���$#"��M�P �Z�Wܸ�g�|����R�Ӗw4h�6v2�l����]ɵy���8�]���Ґ�!y��n�}$���-��ح�:��
}^�+���%����2k��aP�ܡ˄^:!dY��3�Iy�׎�'T�k�D�FP�����]�h(=�.��W[,��U��u�?���ہ�����_�x�"��]ƀ�Ղ�`�y����.5�L\lEl���!���`	���=��mfv{R^�N��`�\��EHr��y������� FuC�to��}��
$ðA�Y%W�[�L_��7�p�}p�1l�:��WH��N�F��!8ȤD=�[���P�6�'G�U��2\e[�K�t�>���0����2bH�W[-��r��"����?�S�@�R4�7'���Iί=BӒ�7��r� wu�E�5��j������^�� 
�kz:��)�oLY��HSF��n��E��E� ?a��
vrt�K�< �h��m;
z)�v㥕��o�$�*/�#�3��w~���Q��ne�����0�w�jw'�':~?�]�X��-����g�hH�h$.�7Dt+��m��[�0��	]%c�H9�y���=,���Cǹ& �m��$������νΉ"a�_�Ubsl���]I�{��g>�e&.����H�E�Bu�m�f="+�F���&V���i�yl�Tv������vw�؝�-�o��b4��o�y��3���e�v��զ��.G�� ����fu�Q�,^�Ȳ��1}$�ĕ�)�:Z>-����KVol�`�K��>�CO~�$�:."�.O�0�*�8Mq�BY�o��'7jr����C>�s������;�H�O��O�-�d�hA����
f�N3Bvr�����U�>Ot��W�S[ax�V���^��wЦ����/���7���O���6���Z~�kju��+L���!^��䀖y)VK����D��9)ˡ�7�Rz�]��6�@b�4�_wO?�[Z��Dآ�X�@JB�嶂nɅ�6�T��$���<5Q�c���ŢF�l�G�2���y��}����$?�E��ǟ�9�!5����w6 �:Z�k+EL�3��䉟E���;�GEf��ѷ��I>JSd8��Z�5�,ALձ�|dmo����ɚ���� ��eY��١��D��b�]���3DCg�u��<�zߴܶYIp`���gA9�!�t� 2a3:���"9S=�����}of������q�4�?L��$ZRr&��~����˅��Y�P<��ןs� _`�����,��=*�$m��"��?x>�HD��r/r�q����<ĀJ�ձ簃j<�Q�
G2TE��6�aB�R�܆��|��[s�'�̹��s�~�X�/��?�H-�!ЧP8�� �H!J�j�4\{��m�aC�Bw��m~,(�E�3`�ߜ�s��S�3�S��g'��9R �in]����P[��k�n��\J�Vk�'��6л��vF�T�v�o2h:L�ܚ�e�� "&�&���A9Edp����lG��X��塋$M�g��z�4������pD�w���3����)�����4׎��..�U���Ȏ��̅NrP�D=�Kcڛ���]�O�$~�N+�|�-c�oz����$������$��������T�ڃl@��K�:@���Fg?����.^��(��	,6o��W�(��#���!�)�L`>j]2(1��֪��A�~�*� #e~�z7ӑ#=�_�8 0U�螬�Чi=����G�	�C�L�^6M%\*���r\���F�į��}ǘe�5��,aa�xqSQ"�]�ƞ���	5�ä���\[I����/F7�i��~4�:j�F"��'��U��\��/(�{nj�O��!���W@��!���hkN���l�@y���3ZRe�_ ���~���]Q/�|3h�B^/�9��h̔J?ds������{%�HR�V-��7�������� �������}��m����0^��4�2�-K{I0o��x7��%��Uf0H���>yFU|�|�@��jL�{Ŋ�hU��Q~#N��E$5����2*-����$��Iz��IW`��]�j�sD���L�n�����b�w� .S�1C��3,s`�vh(#���֏��R��o����5�E#����G��pɜ)����5P]��^�;I�B�B�� :I�Ul ����������{��OnR+I���J$�A��}�߉��v�9	�d�Bi=�l���6N���8��P��kn�[<Oh�虯 G�p��.�����y�k���"�.��a�Өb����\�Е.7�|?�S��x2��&�ߧ�]/�Rt�[�R�
��!=/�&$��<y0����T���2�`����fZ�U�^�u�F��x�Qh��G�C�H��)f%0n���2|&,r��y���!J�k�t
��Z�j�����	̚���CP*�����YN�� ����3�q@������L����.���,�.�D�qH�읊w����V����Ď
ʵU>�hO��{�ѭr��-_��3�81�b�Cmj8M�5_��b�<[&I��pRט�t  ��w��fܙ�F	#��پ]��t��y�y8���nTox��s���"s�*�hSi�k̍�y����>���os`�U�<�7�pp������~��pqn����C��T�彝@��Q�Ĥy�OșI���(kZ���^H
�{5�Y��y[��V��\��ϐc��o�9ڏ�?P\�g~���r���_B�f�o���숥��S:��;:	o��^&߁��=!�:a�����Y�涖��-vb�#]�/�;�Dg,�&)�͑��Ɨ�i6i�mև]l�Q�.�8{d�k���N�:�]ع� ����Htg�ͣzf���+�;��3�Z����Ąh��Q.�:i3|�Dқ���FVį"m�_��V��~�#������-:j�p��~�;^��E!��7le�u3fl�B16���Ac&[B��O~�N����\,+�Ǆ�f�):qX��{�b˻ZZ�D'�u����=.Ж0Q<?�v��ӢA�\��sǨ�œ�`6*� b=�4��O������`P+� }Yt;��} 
P�^���C)EL������/aB)>��U�}�ՑwO��%R�D����<�����HKmҘ���kX1O�$ %����������(�H%Yt<�>NK�#/�f���O�;[l����Y��뾗�T�Z� ����Qo65Y)����J��*y����{�-UA�״�����Bծ|��6[��w`:�/w�ԍ���|��ǂul%y�>n�c��)�Oq6��q{lQ41��Tyi�2�[ ΦH1j	ȑ�^�����L-jh1��VM�����jUsV���������T���#*y�#��<d�]�|�B�6�%ħp�oi� <�<	�-f*��څ/lN/=���b.�:��d�[0�ay�S	ٮ�9�e׽�T��1d����4r��(��yE�����4���46��/>��fe#���?�]\[)��L޴9<�Z'b�u��	��d�L\��{� �X�^~}F���]�=�PmO��T�-b����
);ݱ�J�߻N?O�:!�睥�� :��<�'�Ea6	)����u
����{�2O��
"�ָ�;L"����縟{
�G��N�g��;}��|
��E�&1" �}���<ǿCJ�R���˸8k�eGC�|�u������!d"�?�_��������z
DGD����Q5R�,8%i.����U�p�מ���Y2�����t.�吿�ſ�� b��N#`lx�̯�Yoקq�"L>�i!�qK/X\띺���3��Y86����lC��L:+��=���}V����ڮ�EH$�9�ɉ\��s�k��&��B��
��S�j���`C��$|dK�>��%���
������*�V��k������͛���	w�bax��^F�tl)���3�R�\��2X]5�����戹`޵ǱfX/E�_�����c8�UVo��%��}s��z�#:���ᭊ���-��"K�~ctH�`�O������&.�8L[�C2A��b��m�ޥ�=3�u�\�w8�?����C�ߢ&�*k9���c�R�z	�V��|q
�In��jX�΍�Srw�´�Ķ���e��)?B(e��7�p1��'P�D({��=wFC����+����O|^�~�U�~��:ޏ|��S��Lj�3u�Bb=A[���8)v�c^$E�d�>�ؒ��v2ZV����?����W�Ӄ����Z�LLEO��?򊮌u���qx4�b!#ߦ��{/���]�xm?Q�g��J�㲔������"��6�ʕ1��!�՘�����0[���	5�k�lq���e�0�3ƪ���]��&+�A�9vqX_>��'�H
|<�Ǭ��M�����,>��	���1`��#oX��$��Pl k���C]EO>Hmۮngۃʃ�����fE�x�7��Sb�6���&�vT⛞�2W�ďc�E��^G������c��.�?���>�a�*���?��k.�zF���AT�c���{=k\��yq	T*o�����+"�3|#�����l�lvGF?�w�Sza���������(�aa��~tB�s� �&4�!�+�@
���$J�i!>��y
��j �sO2��oq8h>�6g��8wz�������-�(N���]
4�p5n��������[�-�{����FC/M%�6U�E�NV���?�W��d�41��K$жo3l��vG�	;z@��,fR��j���-浪���	�����B�B�)wa�c������E���h��U\}��Ő�������܌.�ro�����%��3�'�L6���d����ph�E�eh�!Ѕ-�|z7�E�<����w+WJF0.�Сm�|9�����q�C6oX���O�:T�aV��N�	�*�@�57Q�:8�];��Y���J4�1���k*�4	�	�o�xNmH�Oƿ��l�O흼�܂V��'5��
���>F&�U�"KG��C��_p��͎�*=�k��G�������N�b`~�M��&�E4�K���.oSZ^����h9�h,u����$�g(`,�jn�f��݈H��iؖ�:�q���JJ�%ҏ�fD��t��5t�ʪD��L[��Q|FW�X���ϊU�vWGQ/�x̆��5�K��zL&|�J�Z,�o�/ZZ��M��`���R0D���]�R�e], [0�qs�o��>P�x�FD!vk�6�0��1]lO�xnw]3�����c�Y����\�D����s�9��KT'�؁�dl�*Y�ڇ�E-�Yꆿ�\0�Y�2���/��#:�6�;�u��;P�o{�^�s��ؿ���p���}=��u��뒸q��};�B��8ｶҼ���'�,��*�@��|���p�v�0��5��zs�OP0J�����r�����ZEuՖN��KG���T=���?�+u�HVټ9fz��ƥH[q���3qz`p�����C��F&��gӏ4N=.>"�e>w�l�>�>�u*�s'V��1۲����F�\v��ч[�p�O��k����9E$�(�H��~��>4`iG�>B*"���Rő�.��1���;��� �8�>��;�P�|�
�"�<��|ނ�U��]�����\�L�_H�Ms������D�[]����Cۀ+�����(>Ȫ�Hd�6��.�*�58�M�~�zxogvE�y|l�d�Ѵ���߿�rv���V���=�V?�/����g��]�[��%�i�?i������|�ˣ�ƾ����[�-�-�����[#�����B�� ��#��{���i�V���ϑ7�˔���*h^��m���Q:.�a}��~��
{<k�XM�j��Z�a+סa��w6DJzt.��.����X��^�(���C|��2�Q�����1[���S��k,Ҡ[�OO�WG��$�@pb ������2P��v���{�5�b$��2'h,}�s*��8Fǳ+.� ���"_�Z0@+��ƛ�T��AMz�}�o4�(]gE��B���U#��BdW�a�UVT�]����nWQw&�՛)��+w0��C1Ç���u?J(�m�9ݚc���տ� �?�&M.~���O��Oš(��':�(��~W&g�ƪ!�U�Qt%�>�ܡ�6SS�F��[#����v~|񍇝�A{�;�za�'��,?��Y�������GD�(�o#ǅQ|9Q���j���}dο����LC/��s(�l��Y9}���Wٟ�1r�"��t?	h��^���>^�_�%VӁ\w�S��W�_<ٟ;òӬ�Tt������DF^�H�9����.2:��zFo�2_$? ���o�ɺ�2��%+jN����2.�����2)ZI���eå��E`?���s���_D�tR�
�gKS��I��τiɬ?�5|#|�4)ԇ-��#i�����r� �5�>��U�������>����d���G\֦өu��Lb+�r&��YQ��ϼ�s���/~��KQ�c��|�ΤzT�P�
%�E�ЖvF�HyQ\euA1	o���$��&�e��]U��3R�Ĳ��W��L�}���zG�,2����"�̨��HG�]��n���W�K���0�@����rSu	 �QF��8�=��3��bP�������~6�Z��M��^��7Hrl2�AV}�U_h찙RkVj��MXb]��JW<���+�����x��~�e�����a�_p��IK�d��F6� �F DF������J)N���=Aπd�6�k�.%�X߱���mM ^W���F�pnP��P���_O=9{�x[E�!�H�]����P{Բ��:τ������u�ЄS<��9�4�����
����`�۸Z���{���1n�]T���D ��>Kǧ�$ƻmm�����[��z�tyZ���`��J�I�h	��r�����cr�̑�%��DJ�Ќ���ҳA,�����U"�%(a��<��;zJ���0�f�$�H�� ��8x����`���z���\��G��+�)�NůH[ mCw�+����t�p����;���m'���wwϹ�%*�x��G����ga��78q�d~�j��;�Am��@w���ݭ���[��l������MY뙗LMZ�	�=�S����M���3�,��"�1��$�t��7� ��a���.i���T�R���o�V�������E2ts\��V��0O�gl^��+��';��ѡz�
��	�������\��n_��qb�]��d�i�]}VG�c-�UB���#���z��7`pj�u���k)�|ھ1�� Ɋ5D6 h�-vqׂ�PПj����x�W,����
+=�ǖ�S�>�n�Y:�:�$찾���)c����l�%
"c������;��T���F���p$�:Q�xkR�c1��&w�Zക����S�K���}�f�J��1=g�m�"S�	M��k�"��.�-��7Z��&j��������j6:��&H6qf8|g��0	��E	��wjM��U�),oܕy�'HgU����Jt�^�f��%���W��\l$\�oB\�zv�V dC��)�?��O����<b��7��V_�o�����W\���[�̓/�KC���CD�w��4i ��f�%Y��y�j_~�T�� W�8���ױ�7-�`O�m%}�>.)>�h���>bC e�v�Uu�@���q;u�r$���A��0�����C)�a}zu_���E�Ll
U^���$�y�C� �T_��}?t��0��S���#S���~"b����D����⋱߰ܓ�x���߁H��טgRՙ譟��w�7u��l�#� ���e��rc��P��/m�ɞnd�J���U�;�k��s�Gq�"憊Q�`���m���n����G�-�ɡT���?17�T�e̘��*I��}�Fߓ�}W��yQd�J�'��E)��uP�7��V�dC�P����U8�G�t�'^�J�P�R��m�w��n���V�D ^�r�-(��	Y>�a�f��D��k�:��%Ճ�6�ǗlC�a�o��`쾓o�%�s�Z��޿j���^�5X�Nj�/NʱE�$�C���1�n#�|�k���4��e�yk����Y�T���3�Ʃ\����@暯�ҩ������l�ؘ�I����ra��@|J�[୼�pMa4��6x7�/�s�M�g4�����5ߤt{.��e�I8	���y�%����REZ!#��\��46X�@���'c�ak��6Y[j��
���-�V�g6K'OH����}�-��[��LL��4��wX2��A!�F���`J���\������:�ө��t�)`�9V���*��҇���U��8LJ�zL�>h�K���wG 7�D>�6�8�4�fϣ�֊�P��4�9���T�K�	-�f��m�D������i"3�����m7�������o��l�,�|3H �:31t��S2=�7��iO���
�S�Z*T��"�vP^������CS"��N)��p���/��}�
+��LKgi�B�`�cWW�.�P^m�(¿r��C����#�.�-�U
���^5u6?��r�~wɍ[[�.�]:�:8��u����E7N3+�1��z!��*4`�=��b�kXs�F��)=0)���a�w�i�v���ߗ?Dx��C �--u�k��l�,i`
O�4y��	�P|��#4����]:����"��e��e�A���ڋ
�d�ö1'e8Ta��FѦ�">^�V<O�P�?
��ؒ���m����,�X a}�)c/�>v���� o�@3Sin���bt1�PU���z݀G�T����#��������\͉+�n�����^��-�R��o�@��Z0���(lޮ�xu��cazie�!������v��,�Li�'���	D���0n{�m>O9����bT�B��%��I�w��$�ލ�U&��}���Tf�ӛ�8�����F8�GW�� E]�������s�A�f3� �6X4O�b����C�-:�wk��Hi��~K�~�;���w��п��Oƫ��䝄�����O��5�FO.d#�^2�l���WTzM,��M<��R%��|[1���,l�LF��_����PO�!A�H�_&���+�v�C��a)#{"pE�H.$�BԶ3�ƚ�k���$�q��R�w5�`�3��|ڜZՒ�r�𞪊����߽b�'P0I�eaf�O�շ�T5�����/�Y��D|��y�P%%W�W�kvl
�����ǯ�Yg��d ��f�*�b�1G��&�3�񨿪8��&o� a�4t�i�v����a��W�;i)���r�0�o�d5���l�B]�{���afR\���
�xrݞХ�	&��%�-#x5���uM��P]*���Oϣ+��B�W/hga~�oM^�ǯE`����z�գ��E7�u�6�a�~�*\�)��w�a%�����=�x0�K^K����Ɔ ��)��0�A�4U�L��pap��4�u��itiF9�}L�,�����Rٮh�K��1�_��hX_�_XWzCZ�c�X��m�����0:���,ێs�۰�9�?�ApW�%]�O���_�s;̆*��K�-k�-}r���[pUe�	
Ѥ�\��D2·��5����i4��ߍ�Df�U2��P(�Sjӵ��|�^V��^���k�:�h�:�N�bu��֌Ҁ7c��/FR�y���5A��Yr�m���e�QE�[�K{
���X��v�U�L"�Қ���٭��^s��`
q��@�B����}�cwJ��')����$����>d�[s�e�7	�!���K����(K�C�"�%ت��ǧ��?��L�Ȱ^V6L�igqwd��gNY�$�O�j|�_���8�?c�|R۲��ǈ���k?��C}s9	�G�A��s�l�.��:��^?�\cB�F�c.>�lU}���&30�z�A�v-�q���V���A�(?G�p�ڍvw�Ot�u�C����UX֗���V�e�����|r0J��]��� *2��n��u#(�^TOɳl����-;Kn6�mY���eѰ�0RTX5_�K����rI2�	*߈e�[>����;� �m":�%��ȟ_p�1Ϸc���!WZ�+5���/��*��� VE���̅L?�yvQ��L��'��3�aM��%�@�E���(����Ɍϧ�}ki�8.��,H:ՔZ���"}Vw;���'J��^���,�M���9M����ϹGQQ�}ʁӥ�eit)��񍨜�@&�%A�˅��Ϧ3;��%~4zxg���0�j�d,�ȯ�
w��5=�g%�|�q�@{�Le��.���t9~`��<5;��v&}*rR���4�a�����2�v=�r�d��o�w41��ty��ل�r�*��_����N����D���9GW�`H�h���|����|ræ׸�5x:\��?-&"^���Ou����ض��.�����_ 8��S���l/Pc}=�^(`w��5%�~:X:+��6��~��F���+ꇄ�ӐRQ��MB�&��g�%�W�ο���pq���^��3楏�j���_T�^��m������0�֚���7O�W"�jD;xj��rH�f`�
��7��Q�%��@����y���#�2�f-����D�j��}��j�������6���/kW���fu\���{�.�Vv\�dݣ���w��|<��1�܅b4��ZI�J�磙�K���_a��V�]��	���6�E�0�CO�zt�YU$W��Q�4V�[�PڥY�kmArr��K�ԝ��'U�rV��}F��N�eAS|&�޴oM�.� :q�b~����1��߀�E)*��`FVU�(
���Z��r~A���q�'�]$=W��x��-��BPp��H�*��A�K�=UaH�eK�|�9b��.��]ޅ�/sy�:��T{�W�`�����j^�6���6����D�	�����A7�hm�	�~�MC=0~�Yc-J;�����*L�:8s`���d}��C_5y̓�ҍ��VCw�k4�7r-�}A�j�ގ�請�._�[�u�
�R����hb�TؑG���	�:�ֺ�^_�������W��ŻR�>@�Q=s��_FS��w�����?��0�f5M/���ao|�`+ԛ�Qz����&8}���a��ʟE�`?��s�6TY����Je_��D�۷w~�0����:Ur��pv]F�$sFhh�����xZ�u��#��乵��<�,�������"F�U@�Wf3`� 8��$��ŭ]>l�<o݅*�Oή��Cc�(K{3n�D���Y�9�c)�<24�6��8�f��HD����woP|��h�'c9<+�,�J��;ջ�e|嶤��*�����Ȭ�䴣����Q(�k�`�S�%N|{��G��[��{�`s���	�kn�R;��cߡ�PKݐJ��u�������ŻO�B�{1Ci�
���ͼʐL7�=$������w�{���#%|q	�:t�]Ӣ��+�����V������u}���h�je����5�N��s��+�&cYa��)���(v@���c�]��{] ��� ���d��,����c�9�Γ~+��9����٧_��-�$Q,����R�W��O�TL�#�R	_�|�Pٚ�:�+���g�E0+n"=�m��Gp�P��N7�[��{�����h)���}>tS�f{�պ��S���o�m���6[�y5f�I��k��֤:��K��2]w�Guo�}^k!��Ce�א�����nwC�w�ܣ�l�U�[����і.� X����]�1/�I�ڀ�!�e��6bSЎ�{<��r��ոĳZŸ�ُrH���.�q�xx�c5�h�P?tx{�	Cz\��P`.���]v�U�f�E�_�����|��a˺Jk�y;��Ҕ0FJc��з����xL�@���V�pڳyFL4���e�i�({�x&c�����F;�1�p��T��3��/��*o�Mk3�d�H�6,�LX�,N���g���(:�Y%:�?	��R7�ON����Ԏ��s��D�s�3҇X=^���~ǥ_�@�$����%F��)@7~��B����p�<�U#��U(��D��!�*ik7(m� ��-�����Ӆ#<nc��� �3y8���y�R�J��Qع� cDZ�2������X��m_�
\q?س)R ��� �D�K6�,��}��+��pw�s�O��]5~h����b�ûR�^���)F�>p櫓� !��+=��rx��[��-�v��U=�+����0�Y#�c�q���L~����2j��_.��y�ws'G�o? �a����_<�g ��8M*��e��4B��z�
�,��gN,�Ώ��ˣEʰ��s�>�?V��j�|�/OKT�"D%��Zw��a�ݠ	�#5��P؍.k�xrW�Lv:
�|�t�wv�R���K�]�)����g�N8��lqi�倪�;����>��w?�����X�nO#����8�<f�@:l�4T��K��"�A�<��p�l��GyȏZT{��jC���Ǟ���
2��N4+����i�
�w�4KM�B!|��}�q�9ص�mo
v�J[X�|�I��v�eͪ�t��l�O��$���J�G	��.�����a8+�~�h����ϫ 3�1,Cy�M�e*��]��H��C����wZf���:���C3]��E*%I��,��?��>�D��H�2MO�$�fMD�v�D��mJCF�lE�U��ת�#�S*���g ��$:�9�8dJB42�e��b�m��MQw��$�g��t�m�¸��x](g�c���|?7��3�n�]H��ڲPz+�wA�u�~q�A��6�j�a)k��ʽ��-B68���%d,�<���k9wp�z���ܑ���g�<	�
\�yo����W՗j�y�G�䫿��LF�-#��p34�X��NCa#�;�WWР��+�2'�� �;�q� �]-��v�a��۳;|��^쯾�ջ7`,r~�׼�������D�˝��3՛�hU`2||�8�H�Ƣɼ�A�� ��2 :��87�T�Tn{z�=�1���!� -1��;Y��v�_�� 8O}hCFxp� �oP�ʖ���q�p�����H���m�y�'�� Y$mM"��ys�N��zf;Kk��%9#�9�>�pwPO"�5PO����hA�����#�'^s�x�Z:����f�H�Pf�5&PmmJ��G&D���^M�6Ғ����b��y��xv�i"��"G ��=�O��ʥ4 �3|���d�� 43�܁�[�8q����h�/��@s��=��7!�i�_7B2q���j�C�����e$_�3]�W�f�<���5g�<�9xQ�^�E$|�T�3���ua�+�EO��MJ��Xc�L�q�^�b}*�V�Rܵ��?�#u���8Q>��g����n{c�n-����.���oZC(��7���W�y_�g== |�;������Eg:,1`�j
<���R���� �8����}c�"7`��F: �ߡ3FMĊ�G�GI�4Y}t��q+�i��EM�՜{!s��aoK�c}��Z�I�\�<��D@�%�Z��Tz�r�l�=��5��m��[�YYN�H>p���L�+�D+_��Ȭ?���A>�Ƹ�;���ӱT�ک0p�^ ��53
�\�2���ۊ�X�y������<R%�1��z���V�l���Ha|
��@�O���cu�����A����	QשFh��XaQ	I��z6-���M��
���4Z6�@��:qO�/���Ԥ��;�9d�F�ͫ�� d�[z�$�t�]�Vy�2;��^���!7[��Uj��%��@3�%^	�c��^�@?H�i5�M���$x�H��p�Pý��,��_(�di�nh��@���^�T�Q����V�]���OTKv�V'�K-���ؕ�[N�.�7�g	g�6�rf�,ybw��Q��P���ν�Ղ��*_�! �G�Cg¼����DY=/#'�&� �Ť����tϳ�5E��W�~��u�c"��RgSO�Ȑ�O�6ʴ<LaHr��,~a\��i��n|r���!wY;��J��&�i��X�űR���	z���jU&��.N�`�Ze���*�G0�h�޲�CaaI�F�z�{``��*i9�lT�/��ŴL9��]��6����LϪ��2�Q����z�u4՚y�r�_lv����;���H9EX�V�Aׇp��HAN�ͷ�zIQ�D�������T�M�yJ$�G�K�g�G�D�epS �	�����-F��膰e�*ϭ�݅x�O�{7��[�7$�[^ȧU��h_��r1��� o8;�$��4Z�&��eq���J�$"�� é��!nf9��@p�W�3o�g�e����>�K�ܼ�Ga�I�!S�W��C������Bpkq_���Kcb#:�_d�|�&�>Y�l���p7!�	?�YQ����A���tcJ����7��O����43~�A��R���	o�~�O)�q��%fN �� e����>�^e�����8B�h�G���q�5�Qv~M��s�I�cƌ;�>1�gi��f�LMt����zE|��`�4�� s���usx����9�S���Q ۦ�x�!�]�{&M��y��Ng�j=�@)MD\����M�=p���[\�\��J4����x�0l#�e$h=jn��������G8���[S�
br�6��՝��(qu��02��N����ޟBeW���������Q��Q{��:s&bnJ�cd�k{����x�%�y!|���N�x��`�X?�� B�
9�W��ao����>��)�n_�:C?nn�(f۠�}�	ۙ��|�NF|� \��3�ƻ����̽�s�>�9y�wf�*>�o=C�3-gH����%�c�	��˕8�<��I�����'�(���3�[�6o��A'rUL\?�9����a�"�zi��AB�3���t�&￴;-ݠ��������v�x?v���5+]M$�W�<N�s
�f��g�xzg�f���j
�  ���`7Ga�����/3�QN��!�.����҈�_~O~��z1��>~Q 4!��Jг���#�l��<��ĝ�lB���co�)��f�1�������79����9��b���ر	k�ym�⮚&��8K:9�����s�%���_H���8����̳�\�1-�O�Ao��O1&���?���` �=�L�
t_�E� �ם�[I�Y:�7�wk��6��G��[�APmG�SURa7�-��fUK���?^B4�l�3s<Hv:z���S�Ij� N��7g�������Ç`)���SB�-���tJ5|xϧ�NB;%�`L��h[
��a[�:�x��e��n?��d_	F8+gUCf�ŤD��+����d�m�(o���z���D�![�.i�R��{>���\�5�g�u���~�E+�I�5X���σ�.����TC��|�,?�G͊���5�����g�����!��{ g�)���qQ�"M�L# ӑbhb�;��	@;ፓZ�޷��(�}�W;JO�­�2Tu��_��';�Yo�C�x�� ��WA��kL�bʺ���d� ���N�pn@��[��F��:vw��܈�}���s��\����vb]c6ײ��cБ���4�@��)�t��T<��Ql(,s�F	��[�x�Yz�=4m�� oMk�����rĨv3Tw��y��"��a�
�?��$�7%���&j�I�.&��0�ġ��F�a-A鵍��t�E�m9v��5�9�w���*�^FD�aОR��A��1�k�J�,*�KG&n�!�ʀ}e�L2�E�}ҕ"`��Q,A	n�w3��bT���p�v@o�󒌼�<ay�g�νD���Ԏ��n�!�Z�l6�V�b{�[�Q�b�6���Ok�:���Up�)p�@.	+��/�AG1��?Й��s�`�����y=�>�a?�u�vHZ�"�c���5"�� zR��*H��I��D�Z���	K��2�X���k����5������L��QMq��v����.��lhdȸs���!;X��a�Hc$����}�hN��CdP����0��q����E��q���z`�hz�@�*�T{Ͷ� I&�+,�{�څ�e7���������=wb0�5�����j�L6�*�~�/����5���i���)l��$�%�����]M�|c�Np��"��j���xL�K'��(s<�nɥ!���Qz�����+/_ ���$�������Ac�=6�~��$�߈���6~��4|M8�n��;Z����_�ް�nв�����~g��@�? �G� �o�Z[q�0ϳ֖�0Ww�� 9���|�^�T�s���ƒ%���Q�پ/��e}2���r-}&m�Հ>���s��7@ �ȹ,J�I�Yz2,�h���9�oxb�RnI�"���,�y��cr�����#l3�Lo���Cw�m�֕�k4ܽ��%��@f���]�3l��FK+�bǍ���-?0DY����$ue���6���/dH�v�D��s4kBڈ�#;���2�E9x�����]`u�M��9��;��V�R�(.�L,��#X"�|���k��߮}@C�1�ò?UAW��\
��huԼB��5��I�n�s���}�bȫ��J�p��K���6�w��Q{5n.M �kT��=z�Vg��\{���� �cW��1��ZЗ#�F�2}V?��8rS�w-g�ɪ����ᙜPc��r8�~�`zGQ5vv��{�U��x��Q�1]�q9X8L��j�ޒ媖E�<��:9���ٗ��X����D�ȋ�,�>R�E���K�+XH�X����D]��ߕ4s���ފ��!���q	kުl_3�9k�����+bi�s� ���/��K� ���z\B�immɆ�'Q�mѪ�&^��!|ﶕ�W1��A��斅*�ƜǝJ[� ^tzc�qR壖|�Rh#(�maG�6��g����`�$U�d���9�
����څ���p�o�90�f]l�;:�awD�Z�#���-g���B�������Xbb$0[+�����{�.s4�Q�<��.�;Z5y�K����VCÜ�ӂ{=ų#� �3OK�`O���d�B�� zD�^��"u�i(��Ƒ�	�����3e\:��G�`M��֩�PlTB�v=`�{y��YSD�Gf� �a��,��Z0��q�o���C����֙beW8q�D᷎�	]Y13T�$�����x����#�b��U��RΤo����M��_p����^��3���s^i=�;��Ah��io�=^��(W�Ĥ�Di�����<2bv�~�)3���ޗ}؅Rm���}�s���"Ϯ��(�}�T3B(�k�>c���p/)��a~;_[��� �����QSTR�;�,��Rצ!щ"��2�29
h�V�j����-����7׸J J��]�vw�>*��扖��~B����:�\�4qR����pc�`��p�Y��yf|����L����O�b�!��I��4�3�N�ŭv���l�p��N���H�iT�_�y�wn{/�;4�gQ�`R���P��U�`8��F�T�*�p�EO��9��5� �r3��Ȗ}{���\-��k@�L�tKB �J:�Vɂ�n<Ow������5��QE>	�ݯ���@����/$�Rż�þ�3����q~x�L1�	C!��Nl�Ϳ�kX	� �>�1�]yCK��w�1�f..a<�L�u���8,�T��0���v�r�&�=`\řM,[G�����/���Z�b\��	�Hw�ηә,֘Hy-<��HM�`��	u[!��6pr��SH��v�N��0���Df�<�  d�6���"~�𒢬;~,Q
�ō͖<���^z���n��	%�4��9�3�g!�L���C?q[���T��Ñ����L�$�X�C�򬠿���*�d4�zX�ҟ9�3�Q�V�5茝ܮD�U8�0�����fRF��%0�����6�׾b�UZ<`w�8\��B��a`xrs}����c����E#�y���mԗ+�D�Y7����)&����O�؃N���7�~M���������QxF�^��)���z�4�Qw�ObȈ�J]}��A�M�#�8��	<��4�D�f�)�pr�5��tBx���e���&9�/d�Aɬ�?�ڷ��X#�K�7��i��~)�)-̪[���YT�4�z!�ا��$Ν����������~�S&ɹ7��a;��