��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_����m�e"kxu�Uٲ"#oB2�-g�j��h�p� M T�(�P�+M��&�[���+e�ҿĥ��L�.R�d��HH�~����1^^�]-��s�T;υ_�� g|�H�\��#}J�� ���@���.��P���Mn�;gۧ��@�%�vv��0�*n�� K�ؼ����r
O����*�4Me�,X|�-�cxԤࠥ��H�zݴ5G�ǅZڂ|Q��+;}��ӻ�o��D���n��;@�B=�&��0`��ZR�e��M>N��E�S@׃9�=tvZ���-M�0j�j�"$ɫ d2$�Zn�=W~�����7�߇|5��ݕb�B����������LQ��ɘ�I�v&h��V����#���E~/�-B��A�ެ�h%� �y]7*_Vu=�U��&��=G��NoI�f< @A�����=�!&�u���J�qPb�苙�C�X��t�PDb �܁��˼���z݁v���,g5�J��i>͚xT24�zU���ˀ�9�y��n��������,��<|2���
�_���8���n�CJ���%p3:��A;9��̻"�����fPߥ}�� �U��J�h1�V"
��z�կ��#e�ݏ��P�ߵ�o�݌
$�joL�zE�A���}��XN�\�j�0����O�Ğ׼x���������y��}?H��)㒣���d�Z&i���#	%IӁi	n>h]Y������:��A���i�Rn�Ye">������[u���Ή�t���p��v���e����b����opSQPg���tN�Ҏ�AS�5�ȝZ	���_��4$�4Ɂ�2�Q��qA)~x��4Z��v��'�1��u�V��am�Y�#���텝yݠ���D��~�9�gp���ȍX5C<�������9`T	�?������������8�~J��7�����󰙉N�j�]�7��l#����f���ܡLR�_n�w�ĽZ][$1&�b|�; �8�j3'�%A�A���s��"�CnKI��z�c�x��T�ų5Q�(G�Db�4`��W��Fbc���rg���'�}2btY�u�FUD\ܳ��2Y��p]�P�v���r�?~!�{���y��H��ȟPQҵX=i�E��6ꪈF�+�eb�w���+�3d��Sp"4����#�3vl7>'��8?��"��n�����|�}�����VO���@��^�h0���ٞQ1�X�2'a{ͅG���EJ�?
�a������@tF;�f(-z���k�<^�r��^b���wE&s�Q�c�Z9���ԣ;�W���]�m?��D��BR�R�YJR��j9X�6ՔP ���P+]*&�-�,���I�q'��ߕ2�8 l�\��ԛ<�"xhx�JOd�B�w�.��O�����y���$�� �X[􅝓-]��<!@D)���Zg3�1|t�WB��]��T�]�0+.�0ā_�D�k0R��N�h"�I�=��
LssưG�������r�Fd��i��Vl���̯t� �Pt�u��[AS0���^��tّ{�?7�����@�[5�A�E+����S^|cF'��%=�U�́޿�/9��HI�hn>V�׀S����JL�����Pn���o��!n%|�J 	�Wh�B'�=g'Ò�1PK�znfJX�xC�KY��T/�x^ЭU�Ť�����|^wAC��:��������o�дc�g���U�4o���f��ԛ����Q���S�L y��b@��<�/����RCyd�P�t�'�Ze��T�K����<S�����6>��otx�ڪ�4�:����#/{��ù�5��5�K�f^��x��Bi0�������h��w�z��J��Gh��v�S�AH�	U'�JnVP������vB�����2���44��!�ʌҔ�r
5k/�G�U���|&����H*O����Or=��r�ljʒ�*_����%�r���i'�a���������Q�|��O_��ݓ֦�h��7�w��c[��.��"��x
��tq���E����|Q��@����IEg5��e����A�dۤT��sn<�r��ɊC�9�j����2l�2��j-!.��i�^�>�٧nb�,��T�YZv��������6l&vp�m����X�s�N��A�����Z���YvR�hKs$�q�����y7�=z$��aK�$jS%�m�����G�x�UG���~(S}��#�4���Dc��Xl��(��g�������2�}��1���~9�S�����U2�z����4��3����Ъ���Θ���)�w7tp�g�c�\���>��sX�*aN�P��eCK{�Җ[�8w����t���q~4�Z��sq���h�
��x60'
����8��uZ�;x�וW��Q[��Z)c#;K�L��H�}�h�gp�d��`!��3}WVm������=�A>:�9V3(t�A�#6�>ǢN@�>����I�YC.b�l�؇VE�M�l.�I"qȪ+;ꞇTx � ���^�d0��n�\��������6�����V�����|�eb���?v���MV�a�-�7�J���Y8��̢Ƒ;$㱌Q׷���d������W��8k�򾟍��D,_ڼ�J)f�F�r�1��i�uP-2_H��]֣Z0{�m
)9�\��Y�\��" �t�F	U�~[fＱr�&/���S؂Ss��y�E����5��4{{�P����5Ыk=g��<�xd�������BeFb���T}Y�4C<^�%���c`*:K��u2�9y0��,f����L�~lh9��Z�#�yPࡀ8