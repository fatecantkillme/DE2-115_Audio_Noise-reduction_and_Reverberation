��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<�\5e�)���d{�-N�O�rѰ��t�-�:��}���r� �U��W�uE[��W�:�iN� �O��Ɔ�T%��P����!�-O3��[���D��V���__t���L70�3! $�4���b� ����+�Դ�9�&a�Ýc���<\�Tf��c"Ro#��C9�µ�f�s ;�#�=h�[9��e���:�+�}$�iZ��K0g+�Ϧ�˓�O��I!�����+��l,n&�Y���X�2r.��$�@Q����9�}T?�! p|�HwX�q9�7Q���zÈ'���A�E��;㜥v��m%;b�Ǎ�3�zn�B~β��DP�{�{��B�����g_��O`=ae�UN|��83n���tʚK/�fۨ�'���S+<A� ⹡��ҞhL��'6�@ۀ6=f�`}W{��b=;
�����1��M�6�~0r�8�]��������-&M��ՙ$��>�NQc2�reS5��/}�n�ԁ:/�0v�`,o7��I�w�Qf���0I�!y1%�P��"q���L��dj��N��7S�hD*P$Jd�=�|x� \�����9�H�uc��ho���ﴅ�%B�OU��00�"N�2;D�J�9�CZm�څ�|��qP�Y�E���h�	���,��9�R���o��r���H���aN�����M��*�R�a�}�	M}��Ჿ\Q�.�ZHU�U�v���Xj�s��9.*�b�3s����f�s^|�ɶ�(N��g�n�s=����
d�[�3��4\�M�0�)�9��-���taW �v.�U|O�̥���>ǿ�Uo 
������ aF&�~��X��V�L'���c{�~O��\~��]��P��fqm?u�l�㈬�ʭ���Z�i�����yP%��*D��1��4���Sdq��S�-L]	�z��4�>���%�<��[s��K�T7��G����W<4�r��	�?9��g&��������~�*`�|����6-5f�eN�*V҂�iΥ��{t#�|9>P��s`i��G��A.Q������n+�lڪI�V�-�G�"�$7������2fԷ%#�Tz�'�n�\`������bM߇�ͣ#�AP�l�ץEų�a��u]Wj�
ɼ��X��1�����u�p:�������}���-�hTIP�/-+���5�U�AD˸�[UX�)�ʑ��X�X�p`
��K�G�;����%��n
C1�=L����BK/�0�����Þ^��,���Rر�w֨�<Ӑ�Ì���:J�HK���*z�hD}�k��?зhD�'�c~7LL\�t[!u ���kWp����}I_h��w�]fWjzck�?�� Ij�8�`sɜ�b�/Fȝ�F+o�u�����0lP+��fN�*f.��N�4�x�6�P��n��EBe'w��O����E�L�2
�
�0"�^�IR��L�Y���Usk�U�`�C��T���!������Z� �.��B8�:M����Azg�w�C�UJ5U�u�y� l��y�ͳ{�XM΅�ãd�o���^Y�&@`�ǜ�n��d�>��Mb�Qr��^ ���iF	m����a�:,oǦ�6M�+m�W�m�N-z�#�S���%� �mrec�l�C�hb�����D/���gS�jg'F�,��<��)�����pNY����.
�^Ɂ� 9"�#E!ea(�%&P�{ ����r��Ȃ�.�%]���+�/���aŝ��|�5(�x�p
��C���O�_)�숭!��q���,�W��G�0�"&�?bKG�R@���b~�����U�uGc�U�/`�L�/�P�d���g1S<�Z��'��[Z��u��)�T�n�Q��~]H8�,��9��:��F�MI62�ޒ���ڸ\?�-<�w�X��6��6��IaZ��#�}S�$�EIfl����i����Jv�v&�躗hD?>kT��K���d�>���s���DOͭ�)�8������M��R�1�g�>�~v��f���3#q�*��<Ux��])Zd��^�=�!�:���}��o�8�cs�{��yǼ�D?7E��~{�}ෳ��q��m����KHI�z�u�C}�=��8,N��פb�ʮ�Ѳ�}�6�g�҅|�u��2sĲ��x1�Q����?�]�9 j�Wy�i_fsB(�5�����hETE`�GnE��,�����\��tԖ"���4[��*&�j6����>���ZZ��4̛+�����.tMd[����1<�JZ�t������TF�b�����	<s� �~��>��a�mR�ށ��.A	SGgӯ��AS�]��`^���M��s�L��f��7��a�����;���Å��`nw��)�**��jxP�{��^�����.��@��8쏵�n�؍��j�ˋ���E�o�O\�Dw�,b�L5(ɚn�7����'��l%lBf�:��m�O�Io-j�Ie'ج~�n��M��7�Z(r�vƪᲤ|�.-n�}�g(<ğ���(<t�9a�����TѸ���8Ì���O��L9xiJܽ4�Ty|a�h�Hl�%��É�ٶ�Wn.��*��
�0�GBv����9(�D�I�r�����0�SAY�>�~"�6�"�t�z
sv�iX��ut-tx{�!���ƈ_#A%�S�/m��C`�����x$���7K�ܿ�V�3W@��!`��?��]o�� �B�����伖����3x����Z���,���Bosw3��9�Tx�mΊ��;8bt��L|��7W��X�^����[�R�
|
8���9�ki�^���	�,�Q�S?y5��0;����w���>�S'���?ѯ�n�O	Rj[j�Ȇ��`;�鰹U[*R���& ��*w�:��[��W��І�yvX��6��k�_i�rkC���50v�3��T�#�k�,1�'P�f�-�Gc7�$��ѦJj�3�}=��C���Se����]�|^>���Q�Ⱦs@��{SN{�ᛒ������AԐnqLq]˂֯�6xݎ�8j���y�ƶ^�e����ƫm���%h�Ҫ�Pۨ��H0R��;�$��:�˖��RA	Ad���r�|z$ez�����],t*>��KP�ց-:|
��U�r�����üd�.�A-�S�.}���Z�J�x��f�1)UC5���9��c���Y�\J�п{L��Xv�2@�h�hy�K�w�����IS���.[8�������@�v�2�u����.���07���2?{S��E���V��U�K��BM(�]/'�?9�7��N�ܮ�Ow=�-'æ���rȠl�N�8_�����Z�ci!��U�}r �_9W��0[}��3�(���@		�R�]���%c�^�<��J���	`���g���z~v�`D�qͪ��|LX�֘%���	I���틪_�%5��X
�z�bO��x�j#>,���Nd����%d�S�v��rS� ��,�#!+H4\�L�/��2��j���-�UEœ��PF��z�+��dSH
O�9�[�+X�p�
f8�_�{�y������J«8"�Q�MEt��M�Dp\�$���A�����z|��A�R��Ǌ�j�qh��Q�<���mg.�Nq�ED�Z,�=����*Դ����U�;@�/��5Y�v�i�X�TVBUmyG�n�o��Vc�g�n���j,/-)�>�6��C438�">��o��{��Ҷ�ژ�Z�M��&q��=8u�э�E��)�	���p]N�b�����9���f̿���d�4��,��GQx:}�w���I0��ahwKϓ�W!��4��y(�+�PG+�e!�"����j��	ђ$�E	�[��cvU�\7��(�(A�X��B�T~z:1�7S�W�Dk5U'|�)�mJ?�4u�MJ�����D���T̃�d�~��x�p��7�	x�{a*�,i�K]�d�+A�-g2�&e ��3Ò(���+��}�7l��"��9<΄��lva�o	�>5�s�p�`/n�!1��ִnѳ(��e����4v���������@��6(p�`>Fk�>�4-��is����v|�U*�	ҵ�u��Dc�{�[a������u'� �(f(#n�9w�Q�a(��ϴߎ#\�>x�wD��x��Y���ms�u�B��bs8��Ih���Y�4 �_��1E�?:f�n�Й
XJUP�j� k� wdͩ=$��	�;2˗�jѬ�d��.�l�#J-��kE�/�����/ki���K �Ƽ�F��mO��[�&���Y�Y��|ݻ|�y�����R�Iz�����zv�G�!���Ev���8r�����J�Q�����»�b�S�5q�>؟Uq/�"V��eb�<B�	�.�4.�Z�i�!T�DR|r[8�n���$��}�7;���WX.W�K8"�]2����Vj�E�#]Ĉ��� �;�ЙL�Y�%�J\X���+������bd�C�Pum�=�V��،��h��������t�4ӗ�%�q'"�Vʷ:��E�}����=# �b��4��V�,�oB����(����{/�Y_ƪ���5�?�"h��u�FZ5L�ӏ!�8�<2�5rx��+��{`K�n��/�G8�5J��I�i8�y
U�l#��d(\�O3|?�|������k�����9cW��i��B��c>T���� ���J��ꆌ�︼�܏f�ۦ)0�]���W>������x�&��8�FLiRm~�yN�C΋���\�%����@�xsʕ���`Y�E�����p<6M�A���X�[{,%�W"��2A�IM/�<�ȟ�m�l�gD�!3�3¾l6žX���7�#z���oG	΃.��.�=�@����|����w�Oc#%9f�Y�|s�0xJI�ʢ_�r��+`��y��Lv���R���'O���q�,E�'x-�u�e列�1YmE5� )��;����Q��Qm������m����e���}p�@��ۀ0`�.�u�Гq���:"�L`���wph0wJ��Ae$^ 
�J�}I��5rmIa��,/C
zv+���̍3O��?�Nl֝��ߺ�� �����̯�3��٥9n����`�?�LX��'핺� �O�u��?/��H���8�k1C$�xu����_T �����q٧1�i&L�:�wcH��3���=��$T0Ewf�C�a ۴�n3�֋�qd%��e;�z��'�t��QL������:`�{�oȑ�-����G
X4�k�o�_�(K�'.6̼ý�5(?Kj��
J��ָ".<\�+��,5���� ���A�.��S���Z�gcԣs]�!�@~ȅ����!�#�k�+F�[�kQ���(��I�c.�;0V�����x��r�%�C51�B�6����6���A0W����X���^,��j`�"�_�Y��؎k]`z�gT����@l)��g��V7=�}�rX���nkT���Ǽb�;�i'��L�ݞ��s}����L8w�@nr����Bh�M4�9��w���A��ЌI�br6fXhV�/�<�J��'��Ĳ��2�c/�Q�cW��b�hg��I���>�������\��������qh�lt��W�_c�Z�ţ�R]S~>�h�� ����hSB�m��!��SD���SHpJ,��%� �ZZ�d}&�z�Ɋ�{$H,��ӝ�/�p{���E:�1�$]�yo֬�AX(L�%x0#,VC�7�
]Zn2���$>^�i%mv\�=`W+�r����wp���;��zԢ����B����氩�E��Y������RԸ��{���Dz��k6�"�Nc��iT
xU�{&X�,�jJ��HJ��t���J}#I��H-�ي�g��/�l�V�r9l!+��KH���=���9�|�YLI���뼷1�+�-����M��T&�$D����/ t���i��i�,�U���@Ւ1��'R	z~dS��ێ�|r����NJ^>.�@��=��KM�N��Rek�
���?�0#��
�#,�gS@k5�z�-�u�*r`�)�'o[��sY�xs(	á�'ݑ�)�+6�<h�����Ф��E:Ub_�J<
����"P�Lj��'��S��j�AQ�[9x��ޥ��Ŗ��/�����y�<v/o���s�j(֝w�c�3�* ��5Y��)����:%����1j��
�`���ؖiAB�vlY��6L�"����Qk��a�d�����j>{.�<拘�ֲ���R@j>s�`�>Z>Bn��v�g�
B?<�.�La�Hzލα���N�	��[�NZm�:�vڽ؊�;/5�O�����=s�z�&0�����Dhl&UP���9�;�ޣ��8�N��y���I��p�i���b�8���Jb��� (��H��)�v�^������o���g/6e��A�c5k�R��!�n�`�Q;!����il�03�,-4
�� �n˵^5��'�|#j���]���]����mtj�5N����:�Yūe�o����+�C%:X@_.�Jķɸ�%�~@b���C��g������+��l	}�o3���}���@�WX�����0�7��*���*9�@��]eo��س��-�ظ�[u�!n|P����4���@�t�E^8΍�g��x
�����1Y�J��"�(�������!&o�'�� ����oc�R�ȵq`H�쨇�@G3�Yڔ̥����5k��*��Z{�BuFGԬ�FV�,%�������?r3��[���
�PYC���`�ӜT�	�
\1���DW�
 ��?i�$��݀p0r`R5�g��hv��B��B���Qɣ�Y "Ȋ����~����\ �;!��E;4(�UN��mjk�W�Ͱ�l�`V��9�$ް��=X�V��f���
�̵I��Ј�I*Wf>�;�S�]q���Ȏ���Mv�}�?"���q�6����'�������h��� �����;{G��b�
;��o��;c5��\�:Yyoq�Cg�5Pt��&�g�9<@��@Q^���-�w�2��7����9��]���ѽ�,2+�@k���#PBe��*ʹP��O�Y�_�?�6�Q��
�Z�צ�c��F�
�\�jF]I��6F�ڊQx�.�4��(�P
v�4L�9�����qY)X;�[ӏӤHx2?r�Qc���Zf��㶺,L��y�k�uZ�P�2{P�t�֤n�DK�:��@k�E�~�d���`P��f}���dS��݁	'�S�L��_f�:�<�/�֗H��9CT�,1��53��nQ�K;����銨�^��<Ivh#��Xu��!):�6��B.g��Ĥ�'n/�H�����7�;P��>r<�'Dԏ���ԯ%��`J�R���L�����v$����� �̿����2�qϗ�{�:�.{�52mb�V��邐�1��	�ڭ�%�}&��H�sFv����m��'�Ť!B�4M�}/nQf2,�p����]C @!��Lܸ�h��A(�v�G�%��ߑ/sog�O8�NR��cq��I�}A\9�i@L�l� ٘�/Xf�VI'VS^7g����b�t(N`=�3�I�����]{~��8�
�{�.����m�����RZT��?.�4�"�d[T$��:W��~�#���am-1��&Ӻ[i��~��䥻vѣ��Bh�/x��J�8LBŚ�.o���Y2����1%U�K�M�w�gp���C��!��c�xش�.Z�K�4A��Jr�k?�������gS����x�=[Z��}�6��\$ \eWӌ�����29�?���g��{�>�!Kǿ��on�"�����:<��@Q��-�*��q�H�kmz�nO��o{�9
�������_WE��7|�ժ/--2 B�����r�=l�s f+�ã�^�.����|N�}��U�{�:K0��(�EM��I�O�b���*�����v&���i