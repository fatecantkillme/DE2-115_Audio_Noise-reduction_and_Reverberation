��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�8k�)9�k���J�f ۘEN�R��>�Ug:�&�1��"|ܚ���$��&'A������G%�N˔�6EjA��^̕(��:^
ɶ=� �������du���7��#r�((�*%��+��5���<D`�����	2�I����{֒ym�6h�ݻV�w��E�����[����:h}@� �g�îso�p8FK "r�P�1k���"�͉��C]����I*�%]L�?�v��/,�2��H���H'��4�#ӗU�H���&��m�Fߜ��A����3��~�=����{kg?���C�l�j�qb�Y_Y�!�>(aŠ�g�`����3=m��O.���qmU)��?���P�*-I��Dד�W�^��?�̏��6�yB��*q��w"C�V��OS��R�u�D�R�����D�R���b�q%��@��������"�K��K��$�xV�Ќo𚧾Tƛ�\�gV(����:4UQY�U94���=���J!����	#h����{#����:�^��f[��w������K�Q�XO�y��5G�	�ex�&M��*�s�ʵ.B{�� ���c/��M��qٓ�K.R��;H ��)#dڔħ6�������3�Q�d�xޘEpI�X�x�6��Y�e�U�Q��:�,n�r!,����Q�b��(sM�8.��e���������fO����xg�D$ ��Q��ɬ����MH�R�`����.��>�>��K4��Ω��N���RY������/����`��h99Z�^"y�\~�H�/~W�&N�j�ZT�C����_1n[�*R�ԣ4���Qڅ��ݺ���L��He�^\F\�4��DJ栮K6(���J���}{n[�>T�E�Kj�S�x�|�BLG(����Z*zr~�ESzM��rg�{�k��=�b��3GJ�@�g�Da���zv�V���A`dxlos���z۶��q���!���xj>"%9�� ���2xt00��B�My$��D�@�l�R𰣡�P�E�1��=�0iM�������y[�<AU�B۟.��x��
���5g�,��Uf��On��63�TU�m:���)���kl���U��t���WF�>a2.,�w 	�O��j7ە�����o�P�Q,���Gf�����;""�ak�{�V�FW	*�d0S�����8���g�\��Թ�ޠ�MV�;**%O���3ٗ�/bȶ{Q"���he�`k�����Þ�2��w���O�XF����-�{�͡��(G�u���͡�����o���#�],٩����f��y��F6Xz�P˼��%�&zM*Jp}8#OY_�M�����,8�){H�2�� h����z,���˓J����Y���-թ����Gk�?�L��7������bI륞�lH�_tl�LH�֮����r�g}Uq^9�΅0�*�r��7t�a�D�<��N���=3Z�������i�V5��q3ln��A����f���9PB��y>`(�g��K�5(za��&iiI�Q��$���*z��i�
ܰ���!��@���m�t����A��E�տ8(�����7Ʌ��T=$�3���wLC�^�[��H�r{o�~�����uy"��� �8�����1�i��p�ʄ�>�n�j�֡7��BI�ς�#����}�{����*��wF�+Z���P��R*$�r��ٛ�Y���������j�X�� M<��6�f{���?jT#x�g?�w�0�lMi��\'� �;�㿒����zicu�δ#��Ww��C��qk*V�uzFT����������$���?0�[8�#�ltdl�Wg&Dm�9N��If-ґ����>c��ھZ���l�5��^���'�es#���}�Z��-h�o\\%����D�.�N�$,w�T����v�$��N{mv�w�Z2OHKڸH���6.��O�^�¶Ʌ�G�/6�)g��0�W�����vE�AQ��>@T��Ta�6#�)E�f2�$�傠ՐV���rt:贆�[�I_G}�i��^g�t�	��ϙ�Y���襄L�0cr��mW���l6�t&��͸�s�_GQ;���5QA(U��gθ��M�f�~Rb�Zr�/��d9�	���`��=�HUK�k�;V�N�0�F���p�� ��
�.�d�8��-��]����Y���Kj�G�0zP�/f�V}��#�ʗpǩ����R���!]��VQ㵦�I����T�3P�.�5+E
˙y�OTx="ҥ�.9���3�ʍ��$A��leySD�^�_�� �4=��n�I�]C�)&?��,Q��B!פ7/U�|�k���b����9C��������|T���8ނx4H^��%h�]Зc��5Y�f���H��a���(�ʴ�i?���F�c�t	_�T��Gh?r�i�+oA5��f�P0Ė��N�7ܾ8�W8N�mA^��<�R+x8�����G���2��@�����sW�}����a"$�u'���_��G�p��N7��i��6ϡ��Q�Xs�He�Q'm �y!N�1��ԙ�r�~h �>n(���>����_�õ�}�qK�K ����]�e��v=����e8m���C̵�A%���:'�[��X'K;�KB�V�0�`��ԯP͒�+�fR/>�N$	�[���������H��J��L���q�|���hy�o�������v>�Jc�
eGR͐r�C ���>�x]PE���\�ΟU-�>��%�j:�Ӽ���Wڿ�Z��F[$Ŏr��{��#��EL$��n(k���d�?1�m�|q�H0Z�&�]����C�Ģ�]���=`�8UsR�����y��|ԹHG8�� ќ���vJ�8HX�I�J��Η�zX�:������aV������ai+;�,Λ�`�.�r|�1�g��ͥ0�T����u�Gq��y�_)8!"������U�s�U���������z���P䩸,7��om��(�]d0T[�"�g�ng͌