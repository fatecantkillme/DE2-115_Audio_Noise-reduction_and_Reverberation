��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�8k�)9�k���J�f ۘEN�R��>�Ug:�&�1$�[ZwgOL-�c�&7�^��~s/��@�@aN�#VU��؂�6�f�,j���~���P��)��mbb�T�2�����YOF��&]���\Ck�N�}�匌w�~��L��ڏ�5�}��F��0,}�������3�����\v�I�S��v�i�jw%#y�,z��܇dU��M<�:C��B���|��k��< ��u�S��x@���M�����!K��&���폭�edE�ElGH~�[~�>���Ry�-�i���lo��aĉTp��	�e��g���5��I�Ĩ �?!�)ף�"�
�_��I�ӗ����G�h0N���욪������;��vt��!�����xb�ߕL��?N����(WI�t���c�H�X��}9�R|�2��L�%����_��Il��;@88��U~+֦�>ڦ������
z	��"�MXE����M}�k9	RF�"�Ҳ$`Gs2͒����(��U0��pݞ�.����=�H�&-:<$9�<7 �^��27v��q�VIۗ�	����~�C>MTs̼;�J#��������=⮗�b/�ڴQ9��su9�tn�$�%s���F������s�z�L�m�9u�=�T��Y���W���$f��A �s��[^��m��x$�d�т|<tq��f��O�▩c��6s2��֖�o�䎫ï%������ɇ��År݁"%���ܔ����P��w�S���[�S�E��4w����mIi_�oUxBJA��HW�.^��H���J_����,\�KC�
�_k�uO��p	�Ji5�pv�^\|N[)�T���R�?`U�a��ia��n��Y�U��:pGս�g��J���f�nU��<�'q�c>_Q���qQp�x��8Ai�蔙�}K+���@V�!��ӌQqI��ݴ)^GRɞ���;+�8e�Z8օ-�T�yoؾ�<�Q
b$!{�Z��s0g����<�����<�U0.�f�2�	m�fƩ�q���u�A�|XG�-����P�=#�V X���5�y4�^{q��d���V$� ����\C(%����֘�߽M8�%`�Nٽ$7)%���X
�p����
FW�Nwzw��I���L��Ux�iDFDy4]0����Gp�1F��c�d2����b�9�M_�hQeQ2��+%�;1k.�� ��+��B]�Yv����$�O��ۥО���˃_| ��(RR�t�)_�f��U�d�8 ,��ub�_�&[@���h���a�|�Ylt�6���m��f�##+�PO��qa
�� �_ZQ>8�@*�������6�<=���?�؊6�߾�|�}���GV��c���+��!�e�Ri�͜?�C)��ղ̝nS��
�8R�Ͳq	@����1�-�q��F�~/�6�'�LP��Q�����B�Ĳ�kߋ��.�	q-lm���|*�AvL�Pψe������4uFݴ���x��������J2N�7��L��zT��ri �]LJYt�[I���?�-5ԖmA�n�Zu�tr����3"�]~��Q^,m.^��/Z�ϯh�lJxդ�<9�(ϰ�:��#Wm�� �$l�pS�޺c�V��*jI�'@�I��в�D�:@��U����|�M�K�h=g�*{��V�Q��>��Ī`W��)E�+s����9eV@4"z*�w�غ>����L�w�U�_�D�����'�o@BI�
ϲ�n+(�h�"��I)C�g�bgt�t,�v�W־�E���4�$o��ul�r�X��b����.�m��v��#�䣘\v\�$�n�J^�r���W�m��
�M,�E��(c%i�MU߽��	��ү��IH�;0nN��eZ�y�tw 
�.�Z7�nrb�3Zz a�L|��)��?���8�/�V3�v��퍾,�'ǋ�=����j�	,��v��n����I`�,��2{��a[!�
�_�X��U�h����?r8��Y�㱕��IQv΂oѼ�e��6�א)f��O�'��p�u��"���L�m����������F�c&x�)[B�C®[�������������?�E@���9�&�	(�/ԏ/�Y�qB��U+��ӑ�r�P� DЂ����ϼ�*�=Q�������G��k��2<f�O��2#��jP�J���eAM.���4��$��E!��lbNE4%�,fBU��M�g\�Ïbn���u��,u�n���R�%�խ��C���J�L��.t��*\ň��m��j���ʊ�B�b�Dx���a�R�|K���f�v�墅�fy�;���x��܇N���\j�Y�C ���׎��<�$��d�7���D�~o�ދ��Ʀ�e|X�y0'��[��]::��R��@�5C�^ކ/�shb1�AM )��L�q���^LʀL�����Gek4m�
8�ITh��J�~���x�~�ω�ó���Z��C�%aM�͖)����ak~��p��ޕ�5G�ow&����/6�Q��G�;�:���g"n~�Λ�/'� u=�m��y;g������\s��������;/Jh�:I�2zY�al>$�ANO�H�6h�<�R�2��k��g� I�,�'�"b�<��=�<*ˎ��'�Cyn���6Ȕ\�i�2k�IAs2����Ą,�\��Ȗm;�Bs��f���G-6��DI#�H>��p���*��:s�J57�g&Vz��,������=h����D�Bj�dQ�����g�z������n���?5�L��F �cNS<9R^����'�ocb�7�2"�j�(�������#_��z�h��{�:�d��wnk�Q�/���j�mH��b��%�Wx�]�&�y�*İJz�ZF$fEl���\�2��#0�|>��QV���=-�#��Z��LjB7Zª������H�\T�[�3���a#�TōexE&>�t��E�P�a���aQ������(ϣ%!�P3	��[�ݤ�%��猟�������񖴣���{f��������}I�ʻz��^���r5̴��ӒM_�?`�&�	^6B%��o�O�j@y�0S(��P�HBA�c�����}�av����7�@U�����>g��k~4�.㻰:Z&"�ƶn���r.r��}�/�@�M���h9������ i/��$�>��x���mv9�I��V�Sd����z��U�F�u��z����Vg�3dQ oƧU"��ƪ<G���N�6��
��%��B��DV�w|>��UU�5� 6���w���"����1�¥�����WEr��1�q�%ظ8M5�V�� �+��Y^P�ڵ�{_�w��Zj����S�0���G���\A����̀>CSqwv�?-X/� ��[����/��'�[-x�K���1n����Y�����6�擻��l��"��Hnp}��ؘ+{<��l]s ���SR�~/b{��f�!�X d/X�m{Z�S������))�!����'�E��2-�m��h �]�úol�����InA�����?޺�_`ܥ�/L9�n�W�/'�!����m����fp`C������l�.��H�{�z��O�ǑU$��?��M�}R�=���KB[���U3�Z�{����>6~1j��u�Pց*{("�Bf����3����7:�_r �*�+�l��Y�-=�� ��A��q5`	v`	m��Z�� 8ޕ|p_�ɷW�~�8���j:��
�ћ~nY'�Ǎ�KWO}b"�����勞PZBt�C�#j�aΔB�`�|$i�C�aC0\�_��N·2�i��鏠��O'���Z�:_8iȥSC�i*@���-�~����;5e��z3��kr#��rV:��+�y}���|���Z��u��f��XY�u�@#9q�_s|�U�V-�x����f��ea ��r��vQGb� �Yp}���MS�m��ؐ��p�;���N8�ߜ��c+�j��,ԁ���ǻc����E���d<:�E�Q~'�b��q��%�2��t �äor#�s��Q|�P��jY�|�R��\�@ӏ]Ǣ! S_,j�]���������|��=3���KA�0DÀ��Ƃ�t�P�˨��ݔ��=� ��1M'�b#~|�`�c��&)Ҳ��Q����i��� �wfo�B/��F�7tv�~|�!�AZ=#_�/����*�a�4� �>��uZ��T�U��[0�ه.O��z|S��zA=���@�SN��O�:�a�Ӗ��Xf>��Ȭ+lՋ����`&j��G�}O���$$8<@?��i��?��3e��` ��99��}�v���GJ|Z�T�� K����?z�J|ȹt�!�����l����lpi��B���QZ���+���2'I�t&;_ �����W���F>GcϚ4:ڄ��9���R�x؊wI��v@�.�4h!�C_q��1�+Jf�i�]�Xhy�-)}��G6e�?�ЊW���5Y��Ք12;Q�$�܊����2��`�,�U�L+�#���6��*."��Rq/m���N'�ܾ�|���v\�ٺ������ʖ�;�b�8�z��ֻ�Ơ�Z
���ʯ�R2<�VƢ���d����1�o�,c�#r9f�_犷Lp���[Z*FC�K`"H�S�Y�g��)�T�b��z���K�eX��+0�6G����G>*3@!y���j}1�әĹk�`/�rV�z���:y� �s�2���)�㢶xv�=u��lⴾ.���Ċ�{&�� �<�l��9�o�R\��X���g��N��'T��� �,m(�m@�ϕ���l@�yvu���x\p�@���S�b9��`)�2E�Y��_^���&^��7s�#07ox־���$kέh����w+�=&Z_���l���R�kh��s��Օ�qh�j�\i�Փ��cN��SL���8��=M�j-�N���֯�У����-�P�4ZP��lk��VI�[��o�=��Õ4I�������qPc���{*h��nۤQ;M��ZD��,T��#|ԇ��%��4LDѲ����>�^3�$����
<۪V�t�� RƇ%b&M�-�	��rGz��H��α͞��K��]�����\��	�İ��E�ٿ���bq�sE��
��䤼-/��e���e�����m��b���B�?q�ו:���~d�A�z��]0�)���J�8둏-�S]Ѿ��ŬJ��:H/�O���!�5����O�g�|s�; �˭	���~���r�%��k�+�D2��
2�/1:h!����9>�|�v�����-ܻ��l8�g}�J
�|��xŌLd��� c}oh�� Ñ}-֑�p�ԍb��Z�?�$B�N!����&�>��"���֜]���=��ڛV&�vq�+�]*��qm��l�r!���d���^T,�ށ�+�L9�w���k/[nsw))��y?è_)G��F�ǆ�*���'�h��Vv'>��0�������0%e�K��?vێ~������"'MNQ0h�4���Y!YJs���|��̬�{�+ûI���r��ϓp<K� hY�z�oق^	m�_���cw�M��v�}�gP��w�����g�g ӽ�s��`�4����z��I-+��P��H�_H�p�;��:iմ1���D�Ʒ����F}��cr�yϢ�>[L�W�����p.���]�?P����Gq[���F���(v��M�H>Y"�047�wW�ŅI�����ˍ�N3G��>\�������ʳjm�"�Ĕ}[-މ�_>hM���`:��V�z��3d}�@�
��`kEp�W��i �nk㔰5CP��1���"Vk��m�G]Y�k�.����\�zR�=u�x�������A�N� ��u댷�R��d��7��l7�$��F%li�+�{���$8�s���Y|���r��g���#��O(�t�r��1l��L�r�O�k����|�^��co��������7�;^�����`�	�O~��!��2����l���ѢP��n-�cm���I�LD"W��mқ�.��	�S�)�Ĝ+��$� R��;�&�G��6�2|1n`�D-|��.!@�˭!��Ό�����m=�MR}kXQM	Dk8����7�������U�ǻYd�_�B�.�]=b��U����S�:7����SMݵ��h簞�lf#��]&�k�[:�߹�z��n�G����F�,���>�7Ч����^M��"2Tw���҆�[a��',>|���7�~"O����5o����6��Lx"�z	��f0�0W���Ÿ�_S���rwk��3]��Ⱥq��硓���8)J	���^���3�ԜZr�N}>���ǚ��{t���8�0��f9�b�W�')�ڷĩE�0LVldB�Dy5v���_#��ٟ]��X:�E8@M&��<�o�Ч��Z�{w��:/��Ғ�/nL�ب�����I^��¨ض���Ih�QO8A�#g�(Q+��a׸_*]ݷL�c��2��8y�=�ټ��T��+OC�V��w���>5\􀧌���<�N�#;���lX���|Q�%�ր��o[X��e,d2>a>j�2��V��qr��?19����?yR�-Hm��ne]���	���>�h,<`�
�`@]&lrS������x��P?m�`r�xꃰ��x�3�AA�Y�-c\�e#n�&��׏������5�&Q��;
�G[�J)7a��(_�[͒ĹH�;���<��	��޴��
'�����\=W�ΧIe���� �(�3�'��p&`��t췢�}#-��$�����H�m�Af̓r��|�,X�*��4{h��(�nn/�/k���տ��T�<�'�����	 �����ɪ��ỜK�z����o�x;��<a�xY�� ��I��I&���M[�+���Y�H܀ĵ����4�������0�V����}0�	m�Rԟ��t�.ϸm�E��x�Eda���S|��-�]���:U����&z8�iA#�z�&�5�G�L���`�wUtZQ���'��٣S4B9D��>'dą�gbB�NW.|5�3.�O�'2~�׾u�����p���[�7�M���H���������"�������V��̘6���r�s�c�YQZ�xb�u���sdp�Y��S������`�����09�ʓ���N�Z������yih��Gg����ca��^��7�s�x9)����nz������@R�� [�9r[=���:����$
 xš���b����y#�&c����p�Tp_y���pc�t���5Te�{3���4{���tmND�z��l}�VB��D��>%EE�4��?@K5f�44�
��g�JR��>�XǖloWL�G�_��I�*94��*Qb�m�%�us7�	�� ֥�hCcqY֤=����8':`!���ki^�j�Y~�eیʘh�鱧�Vs�j�2.�����^�������$˱[N^�Mm��#p���F %AB"i����mU�����'���~����q�T��1l���[ﰪ���1�n��Q�\��SQ�ۤr>�f��B22�]�i	iabq{�Tr`�!@�f�
&=k���L=(������k��ЀN#���K����O�pK�d&u�}cآ$t+|G�6Ik���r*�346(M{��T*�IR�A�ۓ&몬�J��Ih�.�O0Rc4D'�Ql�9C�Q�m{H�����|_M�kiΕ#�lu��A0F7C��Af닒)y[H�� tt�B�n�� ���q�)�]�XRq�P�� ���jg�4����쉫8�ε<��O�����3��� ��as��O�	c8"Z�ݡ�u8�����ܖC�_n�ά/ڨ���x�歔����ދ�����w6l�LM&�v�j5�����pjF���V����!M�ɨ_������3W��&��ū�������mۗBB_¯��Yy1[n�"  ZEC۟;0E$�"��eM�'�)�}��!F|�5�W��ݞG\[��R8����[��i9V!����N��Ň����(5ѳwJ;0i��0#��`����N�A� �ad�E HJ:D��w�"sb��P>�R\�5���3�rK3�����qB��Q����n�	���/;�fB }d&E&Ӯ�f�����ۖ����N�}Mb�퐁u�Q�G�&���]k���x$R�,iW�a�b/��/o;]*8���1d�	0��M��n�C�pjt;e��ƿZ�G):7%�b�`7pu��ˬ�����	�����~�W�)�ʧ�L��嶺M/x$[�]D�����,�>��AF�r
n�;�[��pe��F�%E�/#hz=ş <lJ����1
wq�+";h'��7p!d������/YqD�rN�R`x��X��~��L�~l����`��jo��l� n�����~k@��΍��v��Q�K�F��P�eѱ�|n�%m^c"�z���c-�n��������7u *K3�
ʂ�rM|p�y��k��V2X@���Iy�U�%��-KJ����0nt�uV��"1�u�=�M���S���0f7�`��=��xU%n�����J9�0�[��G�<��@��	W&����&8q�{�X`r	�lQ}80Zw+mC �-.PT���ȏ��O](�&m��E����Z(�`�>��@YqYÒ|m�z��?]����?#�^	��!}1�:��W>�j*��;���g�]����d�:ū\�z�ԐO��2�E�,���!ڟ<��,"�ƺ-M{��"����t�BG��B�&̽�����>o�p����#��?$4a�@�[�SW�=�ʌ�pr�#�o�}<�!g��7�c�Q
��Q����V�:wk�VKD��O|���gdo|�\`�:�x�[K�jv�{�t<ox��{1;/��~9�<Ny��+�H1l���b���D!pY�V�,��[�KK  �4?6p@5u) m���%G��9� euQ�I��j��5U�Ţ�C�����o��d��G�ɍ��y��X~��(�R%�l��QK��(�]̞��8���CH
�h�}�b��YE)�9c�ל�=`��Zk��B,Zu�'F�a7 ��i׋�n�5�������U�b@q^�����F�t�=���`�s"M{_�xd��k8&�������g��B 
�����هq[���H�!���j�ⲛG|u�d�	|'������Gi ~ֆ'�Y���6{P6��B�K+Y��E+��l�0���Xiͅ�>xV8�5�P�^����ώ��O�?�MԊi#3?�g�ݲ0��C��Ym���p��kyL���f�A��$��p�ic� 1�zud�l�⥚8���'P<�X;<�ڢb�~�<��9d ���\�r�l�s��������3+X���\�R��c�z=���b�P;�/s�xwuڻ��J���6���qQiu����Q���3��ԠG�@B���-+�7l�^E�\�&�2fS� f!1Ih%��7Hp��w�sçu�8�[�{8j�<+�0�3�����3Y��\���=}&�Rn?C�6xM�V�R�l��Ii�}��;0�:�ڨ���|���{��S�ƽ�nrl�R���@6rQ�� �^��h�ZōBW`�* '��zf�v������$/�H�L7^�/FM��@m�	zh���C<N�Ŧ�NgG��d��!d}��L49 b�������Ia7o�
� b�{�)�_7:[�k竔��°y|U���q�[�6��٧���,��t�M��.��"�ǒx�oX�^���tv�k��Q�v�w[�i_�_���M��n���{��3Mԗך�i�r4Q��	��;�9��V�����Q.6��������z���[Y�UM�+t��%c���#i���![ezQ�x]�P�:,7�0 ��k]�2`��"V`PO���et7���V'tC|(�S�}����O�?p�̋<�5N:��q�نo5��<��պYj���+L�.��--�(�B����C/b'��Ƽ�q~�o��*�Ԃ�,c�ڍ��,���%:DBk�W�*������IJ�83 Ȉ���O�F�N �M|�F��}TJJ����dp�t�I;A�LQ�X�x���zڡ��x}3#}(�o��l&��G�d��l�C,�*%�6��F8���8pz}m�
��M��Ͷ)͟��J�����%�p�PAyn<t}���0-:ޙ���1ڭ�X�L�>>�`/U�XNrՅ�q�9�׈�U�ܘ�%�>�bg�}���4����jx'
���f\}�u�mɚ��C���M��ح�3Tf[���QP<�^U?Ɉ���enr&Gw���'xZE�,��5o}7�%��W>_�D#T�ƜF�����iH��q�����H|���1'h+�����k{�lnChݫ�Rw���'E;�M�ċh>�"h�Č��*"���I����'B�i={� $Y愢�Є1� �c��c�'���T�i("�Es�H�+��?ġ��s��0�~�?(�C�򽙸����b4~��Ҵ�=$��J�k�o8H4�K�K�<M�[ �TO�.A4���sjX�@�6�s�
͝��xPW}ܮ_�����5�&6��U������vS3�6,y�pYNXy6�����?{!��f+$����^�F�V��$f����6��a)J����Wc:�B>���}
��@rQ�6���)�8�u\�;�\x8HBtȽ�b�]���T�)�ȪÆ��<�@�$	��t�V�r���7T�,xP>�]Á	.���!�7�`N#1�����8?���GB����YL=�Lj1�"��A暄����oywgU��4$s+��ʹڑ#�V�\i(���b.��&�OZs�a�ȼQ���Pk�^Rh0�����s�V12��J�-���*�����E��
������.zE����y?�t���V�eIj=[4'����,n�ym��X�[�w�S�b��Ҁ-�y˄T�5�˛�+�#�+�i�L���W�p~HAN8&Nl�F{�tv�d*�U6�NJL3Bwk �'�6��^��dD8�KI������|�� pF7�Z9tA�4��x0�v�!L�|��l����I8����k��y�lmTm���|J�s%���Ai�����tv�C,Up$�܀#)�ܑ{��zZ8�OeĻ�:͛��>4��u �y#끭c��h��1�9�MF�#����HB����P]�B�sߺ�!�ߛX��@:E�&�Ż��'�����Q���[
Ȣ���HD�W �ʐt�~��E�}�A��r��m�v'ݢ�H�3�p0t�J��jk�xroh��Tc��.ɣ�������%�s�����HD~�����kY�K��d�?"���`��h6�q{m
��6p�s{��sv�G�t0�ӕ%����1�#*w67��B�=bN��.bY̸�L��&e�Yğ7�
i;H��=�[�$t�÷JF����Ƕ�Y��ڿ�ww_�lff�
��{TA��{%�l�Y"ۂœOI�M�o����T��Tޮ�{�)����jgnX|���fV�����i��9󚰎��~Ƭv��8��H��a[k�b�G	�<����v�/���fa��x� Y���IEG�wЯ$\tC��}�u�W�.��6q����8�l������c
�0j���0Ҥ���N��yN����2��O���%SG��#[���{VAqy�5��Ң����mJ���Y��rw9�
�­�����|Aƿ"k�v�Z��|�ƕ�v�����N��0����gt6��Z�]pX��V�qχ?P��Jq���ok�Nv�ՙ��0���Z#�24f�ٲ��o���#�2����ͺ$�y3%�ہ\n�/vz~�V��*������qcP�%4�����^��b���fp4i� Ǘ�/Vٻ�L�K|'�����?�� tl%�h�h�R�{$5Zm�
dP���6<.�O d�$&�֚ٺ3�W����o�*�[��O��;�
ꤘ3��Ә�O������kR��.sC0��Ͷ����p>�	zɬ,���� ��x-|pX��ǫ ^�����J�P�[,�!`	o��t�\L�,��;���U=�9�v���m˄�"?J"��8��Ji?�4L�P��	�o�Dv�I�X�-iTx7 �M��a�$�qﶆ�8�7��:�i鶥(Z%!"G��tU{������u-�J�1��R��z��7���p�ҧ�V�^��T1�����L��R��AFL�Y��M���	�&A���]���PE��C�gpmZ����Q���?j#c=���?E��yR-�8V]pγ�.��F�1�{J�� �?����G�Ўt�B���!g��s���6N���#۶��lxF.�4I?v4BB�&�fM���5뭾]��jQI��Y']���L�;�#O��zX�C5�.����L3YA(;Ԩӡj�s��ܝ�ۈq7��:8'�����v������U��b������!���Js������3v HkS�ܲ�=t\��'q�WGS��%hG&\�����^Ǡ<GƭvJL� ���W�I�ݏ1�6�Rʸ	��(��vii�~P�'9��'*����w���" ������W?S�������Y�x�w�����ep��tBe��-
�φP~ft��+���F,{A��\o���3���\���v7��ZN�C:��)���E�[�׺@��+-�(���♼u����$��W�V26t4�7o����C+���h�H�/b�͢�e`U�tv��l�[Iw�.v�m��vv	0ءc/������Vz"`~	�$1�f-� ����{��K�S>b9�lρ Hd�%�R
@ �o�nA��5	�Pvac�/�����AYBn�����"oN����nhS���(A0�Gp�����,�s��V�S�sB��1����Gۂ��2(�1wՋ]V���sJmN���2"J,Χ��j�@`��v;쀊���X\�P"��v���"լr��64�l�-���f�>�Ɗ�Zކ�¾�_;�1�!qR�6�*���1S�=�H8�4͎:�Ľ��[M�P�0��إq�}&���>rc�K�}�;�ٚ@��w��--���@ �m� !��a���M�u�J�f�+�ڢ�
�`���n����V��w5�Vz�7E��!�0 ������Xڏ�¥&%6��-/;~3�gD�4HdR(�����r���Ol����uӡ�7,׸Cޗ[���{ٯv�><�T��-/��U�'}LG�X\p���S���^R*6����tť�����	l�-w�ɺ��v���a�y�uMi��L��Pg}�J�@�7r6�Q�xQ���0��E�q{��_����$�_�N�hAb���|�}0
r��	�f1��k�(�d+9 ��h~ Zb��P�����|���~Vjƙ�\�\^֯����?J��sd�
U��*[���1�V[�I�I%�
�f�No�o��9���86��H�E�Y�������[6V��h���||�"/F�.������J2&7�������m�?�Q�IO礨C����2u�9�T(�²l-F0����7,h���6�C�~&�ɾq���^;S`���a��:������oQW��Er�!#K2�7��f7X����_bs� ځ�� ;s�6b9&B���KU_{�zY�s~(��ɍ��6NP/�B�
��[=g_G�Lʓ؊mG_�zg�BQ���54o6<�T�9�#���gޡ���Y�絨A^ ��V��ν_���K��X�G�:<����I�xzQ�vu�)va��޷� ��9gU�ƞuBLSL��7]S`��0�MLKKN�eDc�ʌ���	%Zu�I?k<1��~�P��_���|�\)��Ob���$?����->�,'��t�XT�*�ޥ�A7�����+m�[��wo����1�N���?y�o�F�B�!5FT5�MV:�
c�ǲ��A��& �w��rʍ��!�4@"W@/��2l�۬) ��yUg��q�[��6e�>=%Q�J��#�7R"P�/t���^�K;o��$��D�ϘP<,*�k�q��c@���]�٫":�T��٘5:���3PDuԓ`A)3E���ZǻB�P��� ��h�(Ӊ�+9��(b5�P�	Jt�N9����_�8�KOԼX ɣ��	��rϝfr��m����D�)��Κh�ⴅk��L�Y�����V'�����b,C�<Àt\�>&��+���Ȳňu>%��ʚ��p��78�X�?~�93��%���]-�tp($n�AO�� ��n �/�'��L���Ef���u�+X���8��x��D�	���oh�W��R�l��S�ִ����"ɺ�E� 3���:6��T�^�!���2M�s�B����yV^���o��F�-�~M.%�ٶ5B�����;T�z�49"<�Oiͦ�D�U�y9)t`���[�٠!�^]!j�1��μ5u�����П�=�X���J�?�z�����o��š�>�E��5��`ՕT��7Y��O�/(�*�_&C5}��9M�\4�b��ZR��Y��R���o���@�L'I�SV����-}T�n�I|��UJ1;w�ߩ��sAz�S��Ư�\����4�P���i����R)z���v�3Q�e������JԹ�7"�����t]\P���#�CD+�oE���[}&D	Mq�H��Ag�~Q�}�&��}=�d��j�����G��TV��~�̥z����U����h��%�S;�>i�3�_�}/�����a �﬑��ag��1�"vv$��4�`&0M���[��пn�zQA޽;A-�m�� ��[�Xt�*�p7m�s �_�	�`2cY��8�ϡ?FL��N�p��~˃�����tt����O8^��F9���=+��t14݋c��Q[w�Z8���^R �{�)'A��l�W�B��T�̺sy�Yr��H�n|mw*���R�d�h"�@7�i>��Dh�MfU]����W��M�_��2�O�B�;�~�!f�E,
E�S����xN��}��B��$8��-��a9}�}�.h�O����8f��S�*�	���S�WߙP��&�cI���~R�R�[@Y��~�j�,>�Џ�/��-��͑�;pr]��\��]�̡bU���z�X�s/����f�-����nQS����4��h�d�_�[3���T�x�	EĲmܥ_J�G�ҫ����}K8����j��Z��2�/�U�o�N>�7���!5l�",��k�eѸ5JF�80�i���F�ǃ��#�w����E튩�?�ެ;z/�J.��~��`5m{�?��Σ�]7�r"θ\Rg-n���v�=l����7�B�o�i<r����b��n�R>u�dK���G��V�=+LF$�6B1u"G�M�푄KM�����Kq�n^�*��A-���5Z��]��H��K�\�}�]E���d��@cJ<����j���Zd�.R��ۧ���/Y�6���I��J?פK=�� ���+�Gs'�0�-�B�M/�OJΩ7%?�{�Q�uU�;�A��Q���O,��y��F^��TV�KWv���E��A�h'��k���N��T�!-F�n���$,J_�ɞ�����r֓O��i�0Q��h���d��B���`�=x�P�n��;��������H�W�:]gD��P���M˵w~b�v ���ߩ�����-��19ȹ4�������>�5u�)n���	�祪�j�_f�Bp��f`����ܞ���`��c��m�iD珼*'��,��L�'Ob�+z��FJ������8�{7��G�-���-/���	�J�}��/5�	P�J	B����W���E����3��!�V��.�,��p��H��	X��춍�/��4�kx ������ŗ˪M��U軴����#=��^j<������դ��1��d���̭�ܣ��9�tj�\�[pM9���oG�|��� YG�:a% �m�3I����}�����{����r�6�6�[
H�1#]�0��2���Z�KD�b8@B[hC�Zp����Ա��W�ߎ��$Y<G�n燙�@US�Tҵ�$&A�r�;ޓ����� �AZ�.�\`�q�`ŉMwb��a)�%JR�]��,h�8}J2����<���}�Cd�AS,u�ts�#�1�4+ĔhJ�Y-�H�zٙ5S`�v�+���� H�����������F�	��v�����.BfETv3�$�!wz�����m
�!ͼcU��3䮬nŦ<��+9��I��b�Qw�4'�y����xU�9} "�H�n�b�	��K(F7t��t(6��U�fQ7��]�����%i�n�2R�؉��0�>X<��ΧwY�=�|k��r�e�ڑ����4ޠr��^4�A_/��R1qx �X��vs�����V)�K�IU�GD�%�$�AK%�5�
6��ݦ,T>j�g�7J�NyQ߆���xQ�V�A��󌁫<b�PΛE�����u���$��"҇�$XR�SہSv]�\��IC��_f4��x/���湜B"m�9q4��"n�nZ:_�;�PE�EةP�;���^�{�#����GGFX:���?#��s�����o��m���u��އRhe��ė����@+QϤV��vdkt�6�j��4�[����q��m��=�{#�봟ʵ;��c,
@���7���d�DU��}��𕏥fW�L�ʯz��c�˨��M��?>C�&L��c�I�+�d�R,���^����O$��x�[��LkDY��h�5��q��G�=ߥ�;\P䬫�@#�HQp��D�V�\���6[���v(`!�o�D���-��hH�?�����a�d�f��'������*�qb���ۗp��n
��6姣}��B$)�\{�i#ʜ��l��+�ɕ�S�y:�>���ؙ}y��4�m�y..�wr4:�#c�oȱ�x
�37�ϕ�k<����]v,}g6=n����S�+<��c����^w����i�M���X6�}��~���!a85
s���R���^z~��ز}īN������~�+��0���M��J}�$���w�]��+��;�5|1o�O�E$E�!�ҦH�j�;�I���M��J&�Y�ज)r�]���^şҳ߫h8�Df-�F�h������w�fN�����Ã��ނ�Gm?����'������&�5�]&I�!t�P���1ԠU8BQ�K��H��W�$"�#[�<E }Ԯ��bs(��NY�P��l`����Y��{�C��8��^����&v:�����66�78��'��VjFj�imZ*���N��6��G��ԃ���qN6�a�`U��!����S��K��OS�HY�O�B_$�]��55ޚ�v��ʽ����
��c�e��2ȴ���֚_�s��uՓ'���u�"��d@�,���k	0��.�!76j��2��H9<��n^D��B�u�Z�
#i7iWk�x�;��|��ZT}����"w��������h��g1c�D#��5q",/'�����5��5H���BAm�!/R#�fl�����o����d���� i��Xl����ҭP�t(����~(���8n�'tɁ=��F���P[�'j�|����T�ݭdB]��X�Gyu�y��2,�"��zrѱ�\�u��m
�,ϒ=���JZ9�<?�f��Y��+�Ww�v�E'[67���%A>,� K���?���V:m^,Ҥ�B��Ri��գ�q�Cg������N	��2�h�&t���F#��sb��A�8�$��o@Dd����z���У��_j��*|��E�C�H3>������������a���vacT�kGhl�j"p�o��U\���d3�R�sj���fX��t7�N>!�0A���XR�d�� c�+��I�\�Y8�خN=�*�L�����)o-�6�
騌�ͩ�Z����k"�Z�}i ��G�z���1�0��i�ӷ��!�$�95^ř���Zo�t5~AB��յ��.E�xH��^_J�@3�$L4�ft��j���]�M��L������Z�\�\����eFxsS�z G#�������g��R�j%��:����)Zg:6*#F��#|��̯���[����c8J�o����9�;{�Xi|�/�-"w����#�jD�I{@�Ϝ�gW�Co-]��v�M�e��7�A��R�m�<ML%n�9�#�f��5u���'�����o���q�p��������U���N������
 ����A���D�x4��ɏR�����漈��y��?!�A�No�zcwe�z��,�/<��"k�j��Z3����2�P����h&�D�>Xj�{���
����}B;��ɲ�<a���nJz}���_�Wt���/ᴲ� �#�����@�����-Ԙ/LÊ�)�L�����ţ��N�5�9�=)��ƀğ�?��;�n؍1o����ڪ��5���gE��ۿ�Z$�3��F���8�@Y9�K �t�f��ˁ�$��{}��kꔥ��{@4�bb�-t�B�X[p�z���ɓ��F���P�8�݄�Iyˑ(
�]�ɧ'��$3����n�]��TW�j�����%���Z�bk�7�t/]�|���1��N�7@Ij�>�7��|���3ZE�	���Z'�v��r���f^�K7�\h.=��_4���>lڟ��q��lpj��8��e�\f�A���٩���g1�#FO��*V��ԍ�a�K6wU_�ʹ8"J��)��m%)KM�`sdG���3�����������Ӆq߯�/��D6�0��W���)?��N���\����%�N�o�F9W�b�V_u�$�%���	x�������BG�����Iv���
N�齩���C\ST�LBlD�J�_�L�5\#;팈���3X���V�5��{j���_*)^5x�v ���)��:{�E����YV��3R���Q�o�t�MYvZ��V61c�q�Y��~�x�]_VÝK�8��`��D|V���ܵ�+^O�xv�V��\)�aA-�����8`7�i?���n����+/W���p	�^m7��h�=9 ���L�/H]��ۖ=G�["ޔ��h���ĸ�WE=u%���˻��ĉ.ػlcG���+����A{$q ��B�%TY�c[�ڳ0P�fc�Bޣ���`�GoM��7����mH4��s`���a_� �]N�0�T[��5_����i隫�+����Η{_ �Q�yaC�0�o���'q��_g�?Y�v�(� d���N�z�����{�0�ׅKIq��h��R��7&	��74�u�-t��͢�!!w8���I�x�����Z�~�V�f픆�Ts�����%l֎�
����$�ZK�v�O`�9����&�RL�J���4�|�,l��ϠE����Hz�lȋ�z���M��w,���$���8�z��!ٸ�TWQ#X�ǵ�Ѻ��P�GGϺyG�����h�D[H��^�LY�\��Y���,@����F����\ֵ(cybۑ,��O�� 2�𜃧�Xp�ׁ+[_�+����kk�m�$�[�������3
R������1��-�\�����jp�`���%�����,0XR�>�q��`B�������*xѕ���Vܗ�8��b��]͆ �P�IJ
�)�q�M ��+���^�1�F�k�y��}*���F՝�w
���+}C����:�/R�]�J�4�*���O�5D����S,�.�M&���G���.�?����Z���	�̺-�sb{=����w̍�����)w��%�g���4�c;�����"�E���%�肍�������t0.�K�_��+=�E���=�Z���4�!;c[9�"�⇀�Xb�}�x���+�(Ra�	\��,#8i�=¯ ��	pE����-]!��R#�Jl-0�1�uN�,Y\����l�Kr���{s�d�6̉�1���6 ^����e��\���X,hٌߤQB���m��b䃵L������ܗ�����_$k �(��'$O��*��Z1�T�'R	%����Eʀ屔�������v1B�)��@���Mԕ�tP� .+Μ74\��$��2)��E�/TaE��Ŀx���P��F��o��LN:�Z�����u������ r��9���J���d����˩�����rE�~�hl�Zj߼����f��\n,�m���R�_�} �$���{����?��1{�b�ߢV��@��wX�I��Ȣ9,`�����_2��b]]��[[C%�i޵�6��`F���!&3��⎮�A' ���uj�_U�<���7�l$:O�����|��0�+���\ܓ��:���X$W�oQ��ŏ�e������v�ƿ��F3k^��S����ݠ��m�	_K#�� �)���Q]�f�����Yeȭ��C7�1i<�<�TV���Q٣���*�'����Kב؄�*�>��l_�Z�8�p��L=�*���C�+CE��ч)&��LKx@���@�O�48:��7-��K���-�J$�u�`�
�)gqK;FX�]���������e�W�LD*t��xAZ��)�>]z�8�y7����|m�QX���%��! F���%耿O�q�R��pQ�zԊ$�O/a�=��h�9R^Ǫ�ux�
�:0�c�Do��9�$����ѺJ�-AȄE����RD�{�T#���D���SC$iS��5��{��e�����~X��T��[u &�-b;�N�"�l鿊�{an�x�)�w�rs-�)HN��:*��_��Y�;m��[�`}a�Uq�F�n�7D\I)��îo���a�~wD�?�\��|��7�> /x6����R�#�P��U� oK�'�$_����8����Zc�.��W��L�`��O2��>R
(Pk���ӈ_���)��@N���pʊ�~^���r����iX�"��	��	>ݷ-��Nb�o��(H�S��xv^���h9Y;]bf����$t5�_�\nv!-�B��OB�$=�����d�;����UEO�;���x�$�-��&[n��oEe�؜��$�*�fM�֔�}���+�&�cN8DWD��ف�
r����3����z�A�dJq�Y��1�r�O�f�h��qEm��L�æ�a�f�'��g���V9G\���ēns���%�0|P�!ޒ!)(��`��񇗑 �"pcL���M֑DY�-WF��ʘ�gE���{󦹺\�����Ȅ��]��f����ڞ.����iz,[�\~�1+�2��0���mg�_�*L��D�QV?��B�Q?h�҃Q�B�m��c�"�������gEB��f�8�G��N���m����!���Gq�Ͼm���DPS>Hw�^��w0����ʑywCv�J�Q��r±P�u�P�舜*�/@&���K�I��;lZB�A����ۆh��s���?�������܇|���0D�s�$V;����Fly�o����pDC[1�'��Jk)r��]S�Ļ��p�f��g�{,(�ȯ8@)��Af�N���.��1�	�;�tD�Ӳ���߅?-Θ�A�
/�q��1���L��XŬ�� �<�b�s!�N.OEK�M����`Sq���0 ��	��6�%=2B�d=&���6�;Y,ĪlY�U1���GSp7�JWm&��g#�yT�wà�k-1_�ut� ��T�o4��[+k�1ٹ�ȚѦ�����#�[b�Y�8S�K�e��C�A yƼ�~�$ R�\�t�kԚT'.w�~��nY�2u�.��^mA2�P2�P:�z�F6>���1u������l='���R�$�?�,��DL"�޹\qP�!H�x����4 ��]�~��7���g��;�Y>�x�tV,�l	�Z���{	H ����f,�����2�"?Y-lN�Ǽ�h�d򴤦6��0�����z��x�~A`��������D���_�������~BjBq�I~RW
�?nO�=n��H��n���)��11��^��qoo�w]�͜���=A�H�g#��,�w�R��&Y�u�1�8�%g�"z�/0_f�n1�V��2[_I���j��;��X�t`��9X~�U4��A��.����;)��VB*i����͆���:����f�Ά���<����G�υ�D%빤{V��K����I�&��=�`�v�Y���A��������2�8׹՛�F��m)O �t3R��+�+7�m��nr�g3w$��x��"A������(k�%],d7ϥ�n�i8n�i�%��pӼ~7����r��_��@$��3m첺n��4�:�?���Q��}m|�T�U�YI��!L��p�ſ)��%�{k'�w���l��I	���7�ײ��cN�u"̯�& i��a�ͥ�*]х$�Ğ�K����߄��=�%���kY��^��;�k�}�1����D���3�g�^O��9�A�8r-����=�����{/&�2�߫������ep�v��BO��->MY�h	���Q1�EX58p*��1L9c�ݬ�'��Y��ｮ8Ҏ^X:�]���e���S����͠#%W�za'q�ZX�)��M�+eL��+_�2�Kw6�놣��"Դ+
��	[�=̋�Z��1C��{?/|V���q��^��d�j&h0vR�[��DD��Lv�|}�}�$(�&����NF�E!�}�P�VX}Q��=~6�,j���qԍ0փ���"[�k���曂�#؆�_|C��������N�X�a+J�ʴJ���yf�(!���e��/'<Y�5���pitꅟu!4!�[�d�a�i���/���r�ʊ�<x5��Q�2�����a��U�'�+�f��nDza�
fnp��V;���_�X4�$���=T�F����7�~����hޙ�ev�����^���ܐ*ncwҸ���i_�t�W��i+N�tn�-�-�.}�$E�|�r���ܗB>���?0� >GM�0lL�&�S;�'A��O�@Qc���m���͗��cC=�d35�<M���T�c�n�#۸���ivB0�CA�8ar�a��c��+eV�&S��R �^�8!k�z�a��vb3��a��d�8�*n�ؖ���[T�:E7J����&rH�f�ȈV��	8�~rG�&`�`������oDD"��8�J�'����SM�Z�U?�?�LVu��p\��U��e���LVf�lJT��nm�`j���O)��EK�����&c��o)��֚��
�����(�e�4�[Ե0��{�1UNl��t����3�f��P�?��k{�G*n�����5�,' �x�ɟf3�-Vް���*�M�I��t���PȲ��1AzL����(���݌��738Ic�Z�)����pV)��a���|�߃���M[���¿"W�#8-2��񏨊��;����*C�:���~Q�ަAz�U��x�=v�F���Ѐ�����F�S�����x�Z�f�>�\*�e.a�_�BP��	3H��/�E��:#RĊ���;Ϣ��r�������2�.�ڦ�Q�����j.���9�1-�mw���4\��C����������t���VQL�-ƹ�������;�<�CV���:�~0Zg'LNʩ�/�.���9'�.)�1ax#--c~MM����ha��ͱ�<�A�n�Qnxx4a�����������Iw���2�� �ehK��ٓ��z7��0S6���1�릾���S��u ���B>D�J2��C��i����s�
"D�(�;�DS�h7h���'i����uS���&�?,d���Qϖm�>�n�z�+ư�+6ގ<�96�'~fI#i�_��;�AUXhA������ߕˍ��/��7��򛼑�EV*	tf��;p�[R�C`^��ˮɮj���}�r�+92k�����f]�D�k���P?U�g��7R.T�X�s��$�ǜ���c�ձ��Թf�^s�G�W�g��PN~_7�����n\8�	)E��T�%�5`�ͽZ☕j���1PT�E$��'����U�I��F@Q'[�(��F&�'�9v�(��G&��f�Z>�>��va�WIb-B�N�y��C��ɗ�R�E��B���ژАܪ�7Jfua_#V�V���G�&ca˘�F50h#ٖ�r;]�qc7&U*n������sr�����J�3l�)��"�\�pLZ_�����Oצ#�W9��hS���Xgv����;
��@�9��<Πu�#ԖP� ^h9p]ګ7E��.lk�Ž!�r�U��:��#����`ɀ�+>��+��YC�C�FQ,��a-��ؤF��a�Jt����#���f��{`�}ڏac��~����%�t�Q�Q.���u�ͣ���үj��Nz^��*�id�I8ȇQy,䧆V�/j��̰�85^�u7\FIg��}��]����
�*��}L�a�(!x��D�J>H��#t'���}~|�n뛳��&�Q_sg��h��o�k��<��m�+$٩5<	l���#�!��6U���� oZkݝ�3�Q��|Ț�gɐ�i+B����k�gup�(��-W1a�e&l���(T�e���f9����1oT.|}{0W�dINz/�*]��HNN)D��@�m@^N	T|{�t�7Ke��� ��".N�[���H]��������'����^c+�����Z�U��J��2mY0B��:`Ȏ���\���Y�.Dm��h��[�U5�,6���^�{n֧2�*H��Mc�"�X�g5��?E�BCd0)JY鞏]�ՠۚ�� ;I�5U��	�f���T� �Dy��`�
;9��u���`���\��&w���E�=�!�'����&�g8�/N���Rj]�Q���0�P�:%AY�gd��_U�T�5�~٫��J{�zp�k��Q� s!&�����B5h���m�CZ<n3��g�\w�,��幌�A��g��=�Y��8�����h���ćv���n��yr@�S�"2���@�l��C�����qMXxb���p���z�Ȗ�T��r}'�� s�ʣ���QP��H��� ���4�d���E$.�.09�'t��.iʚ��F�9��`J��7���g-��yS���i��Ot��(�MMo-�6���iD�X�PNc���@���ogȿ���K������Fm�h\K0:�
/'����<z	�������]�KE2�)���lmj�T��ros�<M���Y�&���#�x��A�Lo���.&օG�I�`q��ٹ��&�����5P�d�9s@y���we�� �Ƚt�=���G�V�f���v/�Hye��� ��fK��{�檔�����@Lws�G��VcO}r�f��ƕ5�;ɾeO��d��(C(�Dΰ���g�Т#.w�������%^w�鷊ڞ�0L�b�>�k�Hچ�]���e2�9~�)�YrԦio�7-C揢V�1uY�RCm��+Ί�-1���Q������������4���7�T�_}���Q�c=��[�w�	��C�DG@s��˳DT���ߤ���[,|G:FT<��#�}a�ȳ���w�*r��%������b��C%J<O%��dZ��}&Ng�7�?�x�䙗��_�k+�L5/���>;s�K���Ah���]�{��@�A�q��s��-�s�mVF)Y�MJ{�+v6��O���tHv���JQW$8?<³6��X�;G �0��������U���p�P�j��29��'��� �ȑsX ;��X/�������u���T��A?ّ�� �f$k�o���%(O���4�eE�%m��1������/�+W$8�o5w���g��0�״�)C�6�Pu�.�ĵ��(����k�#�r����W��G���"T�X�tL�(8��J��NѤ�j��z�qQ�-�JUpH�Me���|����;��C�?7AQX��Fz��2E��j�N�o��5��W��v�R���?u�7�lrw�>,Rb̀��e�;tm/+J[�?Z<k����䈂ĳ��C���Z{@�I8o�Q� �KjK�J� ��P����&��-�����A�3>8�[�ڇ��b�2�|4i����+͟U�|L��+j�5
�������&������`���b{Pl\���V�E�s�Hs����!A�u̜]`�L.��WC��{��kp-�{҄�q�I����cO���[�q\u�~�a{�����f�J�1�|]���aWLx3�~����G���ѐ����m��ݼܐ8yd�ܴ*Q�k���FC�E& '�k2� Ņ
����2mgI-ʸ��(���W:�Jû���~%$R�S�ܣ��?R�AX��x)�;�r'�����۸�+��
�<�u�ij�T��tĈj�)k�1��Xv�Η�O�c�2L!��*Cw�_�K��sf+���G�ڙ��.��Fƾ^�<+�L��|����V��0��cZ	���{Uw�C�N�dكW�j��c�	��(��o�x�2I�����������\�����7�����L��Y����(~�N��s�OZ��_Z�Pɻ�B�m��ر�zW��`VSJ����<�J�tᾨ����ߚu��Ë�N�2mU�j[�rˋ W�vCq�HO�Zs2��.�6� ��Ut�$}e�`q��	9�8^���
�)��y�q��Z��c֚��Ibf����;��X�cN��G:�0y5��r��`�K�J� $�L���F��n2D�ֹ���{���6y��2��wp�x��~y�0zA��$��ݻz�N	�g���!��b�� ��ٳ#^V��sK�<1�|��}]e��Ts�|r
��,j�����C��~ig�0e��Σ���h��D�/���X���5#4��K��I��='�,��>��*&I��9h.bIt�l�^R�E�pr\3�@2�=J�m�P%�Q}C�m�����[0�{O\�@P�Y.ا�,^Z}ě�3O�8��a���M�-��Я�o��\d"�M����!`��_h`�M���V�	Ty��[�*��9�?5�?��V/�Sw�NEg�dT�� ���7���c���U����H.b5�Oy�1��Of�?+wR�t�q�f'�v�M���� m�L\�!o�S{򁜀�pFW�r�B��)A�s8VRi����eSbBS���L�Z��]*��n���v�]�<;{��mVë�S}�#a��So&�*�����M2���\K����z"��n]MR	�z�Ui���-�w�Sih���S�C��*�uH��!�	, ~(��g��}=��vi�0S)~��( ��4W-Fҧ���G��B��Uz��*��,n}O�8ڼt�3,��{2��1���ǔ|�6�S�V����$��
�Ȑ����ϓ	��
�~e�Za�V�[��<<!2��MP�s)���'��t�cm�n������F�fs��m�+�}�-�z9�Q����y��*�Fk)T�
x���N��ڎ����u{L�z��L���/_�è]l���1�+��x�1x�al9k���ݙ����K0Y�"t}�ZH�ub��w���x���QC��W�߃���I�T�#��T�R�"o��$���#�(��_���آ�n׹�����u�{`�1T�ΚŎ�s3�7�����og��lᒗ�/9���Ј�~%�����DW���F��3$#�i������+.^_%�y%��XhI�'�M��9�K2Q	5�`2�|���i�bK�z�Q����͖�eAp[�|?oG+�"�����';��(�d�
1[�"K���n0�}vn��o!]��|,�G�i�0~s�o�'6�=�iv	�}_[2z��l;�V7Hlx��ȸ�щ���s�������(�>�����񽥆�|�pǣ�R���_
�v7� /�ڛ>v7}'��+��"��Q�&�̕����J��b���t}K��A"ʖ�k���y�@�O���);/H��77�S�?N7ZE����&f�':'��,?������K�Ȩ�1�>� J��Nu��R�8z���.�5 ���O�kS��$`�7��\�Kƹ�.�ӡ=P;U+�8}O�Gr���=�ީ�^iװ�{W�6���GS;��O��ߋ�����&��7(�-��lŜ�I�	M�'������x���O=�O ��EI�WD�����fݠ���ӊ��˨ �Ҟ�f�\�'����Z'xf���e����ؐ5=g� ���Ł�^�V�2�����^p76ub����g��i�ؼ��yĪ�w඲�F������D��:R�R5�8�%<z�/O�Ƒ##R�R�<Mz� �&���ЄQ-��M�~lO0���9z����Ɏ�� PF��ڼ)�-�.Ԧ�$��9�V��B6P�kp��}�ΤM@�	�7���d���c����6C,�2$�RYj��un��In��h6YC����G2yߟ� ������5i�4��d�X��&�
��Dd~�F��P�\��}d�VM��rc�;����U�
�b�AAn$�O6����N�=��7�X.6��E��mP/�N���Ğ������փ9�"�.��tb:�����s�T9�K��'��y�,Z�}gwJj�fZ���$�J��Je�Pㄅ�Āw��A�;��75v��hEn6q�˚ZB�&3mF!���U��, `AY�"��כN��Kf�cb���ž�},B��usؖ�[ꔲ��C�.L8�"��Z��ݵ1}�9���e܉c\ء�@
�v�2C��<9o�#����V�wM[#�_���O�]�,�G�����8��yw	(�J��<�κ8���~�;3�܎���t�����6����I���|��[�["%���i���B���3?f�\�|��L��ӡ�+K���rkx^���	�wH�/�k�S�з�6J�*�V��"_���B=\��N<��f�M��9
N'پ�D��d� ��P F=�W�aB�d�v��&���2� ��z�醼���h�\���,�"�]0��jB�'���WE���kC>�_�-�\��Z)Ш,lü���LʾB ¿O�,��a���|+hb�<� �7Q>�c��a�Ru���)��>�0��H^��&��9³X����.�t���X�B�mv���FC�=+7�ּ18� �%�u�B�}5-��&%q�b��;�~����6�򐜓z��;״��6 .�Σ�^�ҙ�N'��Ǉ��_)(|w 6�+Wap����p�eKM���΅�c1ȣ��v��~��$D�e��Q�K��\tb���\x8.f21(���HI'�%����PG!���M��2养t����{�OǙ	�8�����@3��K��[��@�6���b���a�04w%a�|��?��eKٶ�r�ʾȎZD9O���m�h��d^�� �?����.�̯Bԕ1↝��螘�V݂��h��˾I-C�3~�7D��t)��F?�6�ÎS4�I�����!NfCp�/1��M�@upl������sE���.��������DF�VG�%۟Hr��N�\��~]�����D�C�$��E�s�M\���:ߋ���D����a3O�_2��7�b�D������N4��;�ؕ���-�C�����gz3��E���`4/}=�Zl����H:�iA��e_D�F]omS�p����$9IL��(g눈c��/���lď�Q��ޭ2q�T'���j�(���'@�Ό�uu�$ց[l*n �F
���b�A�%˄� �̥�$�թ��Y�M>=D~�����%'��1�Z��%}��LDӯ\1�Ͻے�X���T��� �Q)~K�`���ԑA�tf���`4��L���%�}-��g߼d�ﺝ68��
9w
:�;Y���Q���\G�{��c�6.��G�f'R<f��e�8��pz��y�[�[��?~�l���{�Iy�M�r����Z���4]�-m����Yza^`"�^d�������H���,��,A]�I2�Yk{BppTn��=��ݕ�)�VV\�_���M	��u��)����LS� �S��Q4"_�(-(�
m�Ƴ� ֵ����,�w�V�nQ�6��G���m
Z�z���dY|����&�(ggf�u�H'��2ݝ,�
cTx�Z��T�S�>C���)�=�=����n��L�'����V�bW W�/f7���&1�z-�tӫ���-�������Q2�D�(�(b��s���H율�����$��)3�N+�3�7�R_�mYk4Bs%��(���^��ݸ��& Ņj�M�>�V/p�&S�S;��^c%�p�+��"�,r�ݱ: 3MŃ{,,�E~�_�;�0�{؃H5#Y�c�KR�H;��yPR��h�+��lT���L3Y�ka����1x��$���+������a�L�d�A�=���O}�*��m��s�Xr�G��ԄW���`X��}d�j[i�dUQv��@gғ:W{T���6v�
?�$��]W��6�N�L�vY9/s�}�e�$Pi+��ȗ/��]J}h>�P\#�b��f�li���ug�)�*������X�c
�/Q�+����;V���w��A��+?�0繐,ۭ{�-�5��ƺ&����׺5'�܅}z*�kL*�Umn��8��'�"���Z�=�C��u�ۦ3O���3�������%��Lg���v���"�m{_ˮ�hQ.O�e��|/�*�6�<O��(�9�D�A{]�#�<C�R�«%��i��1�fZ��TU�C/B7	W�����@��*��y��Ƣ(�_�����JD#�g :3R_��3у�~=L�О(��	���g�1�@�
�-�"��/w)��Z�d��ZT�5X��D`N�88���iO��/��8�k���Kd.S���[/Z`<�6X9���J���l��{Ud�1&L5�V��%�Bw��mȗ��Q��?��`bC�'����7}$�Z��
��))	^X��BXJ��;X�*$*��S@G��m��('t�ŋ,���d�TE4>�:�R������I��2@ƈ��k��%����a���`�-��bܙ�U9�!���oof�@����y�r��?�Yq�7���S�'�\�����o�e)�p.z$�9߀f��bS�Q�FY;Z
�d'�����L���+B��l�p�6�^ɂ����v`�9��inU�R"���ΉG�$׫iB�e��k�x��<ye��r�2� +�Cl�U��ԫG($�&YIs��=�3�^"@C,�}���C�>}�����&��W�� &P�WÌpʍ�.��&��Y]��-e�c�Jp�xD��ȁYf+l�`�������X����h�a	9������6�Yhˤ>����O.���	�Zj�D^���r�++����p"q���?��VU�˰�"�ꘃ"�É�P�/�l���p�9J�x����JDj�F�����"��p+#]��<�$1��II"����M87�NW#t���)"ҿ����˷��9$Z&F;[��5x�>[t�����,��������
Lo1Abe*��Ձ�G��}�i��\��@i��F�����5VG�6��l��E�TY-��L��n��%�ܙ� 9�kA*��^d���0�1�N���%��H�NSX=U�/L���[����t�.~�x�G��-F����PU��ԏ��@a�R��Ar�*E���r��)<(��H<C�_k��V������ľ�ՖJ�מu'��U�H�t3��l$��0)JP��ؼ��1�4 oǮ�����q`��_�"~X_}i���n������ٍ{��|w�d���߭4nY�z��q��Q78�1��l����4jA�g7x��H�h/�r�qc@�`���[�G�$�~�& �{�t�?�R�n�PZ_u/U�K�sh�1�ހ�bI�S3<�N:m�pi�>�+j��*�7w�CH_E�p&��E�?M&X�%pu"ķ�c>�/R����]��bH2x�f*�p>���'�pD��'ָ���s����{��C�o�&�S=�hcg��E����b�(��ܴ��J���"�	��[z�~�pk��kY<�]�Z�S��WS���q����Th�B�0���/�R��rL�T�s��H��KӶ�-����I�Ž2t����Z6����Ԗ$5��d��Qe�[hIڵ�ԯA�c_�-�)�j����%�ju��%��(���+��qb.������	�r�Ӻm3�CS��;��&6����Π'_�3��*��,�l�Y�����Q�L"#��A`���Ud���uVg���7��O��%ĨX�����b����K�T7�t������ȧ �b���:��˒RZ���i>+��;����u��(@J1>����YH��*�fK�ָ�zY�T�o6ugU�v:R-��<�����P�P0������y�r��������������(�,1wpe�����V=�c���H��.r�%D������Ӯ?��Ǣܫ��]EGW��г�9� �Ā�yֽgKq����*�?�"�J������RC��
��#;���J+5�^��H�	�V�Jȯ��>����FqЯ-뭃��Re��#B`����胣�ŕ(�G<
���J���U�g⫂}�il�l�Z��$g���F�Ĝz��&�	�~l��X;��&'s�<���.G�'e�{c�M�z\g�����wɤA��̣�84��Z��M�U�nr��0�|��ZX;�"<O�a�C�0�B�" ��ji�.松�ǵ��5���1�}�L�	��ָ�Q��myM�m�T	є�W��6��`Pu�g>��(b��g���Yߜ>È�d�Uν��Xg�{�	�g\�x�K�i,�$=�/� 5�6���[�zv�#�n��8��<�+H$�H�LYo�o�����U�k��6R��?���Hl3�TV�+өZ�G+)=!�P�����'5�a1��܉K�Z��^�i.�g�ó�`b���GM�ss�9�l�i�9��C�wU'�?<�<�/��Ӑ�7s����_3�C�9"
鴨1������?��/l0�����E�r8~xM��-<nzk��ʜ��;�`
]�BuHuzci[�x+Y�꺆YLK�+7I.�|��A>�����,\[ypMt\1O4_@V-������˨n�١^�V��ǝ��$hS14+ftV^��%�7g�F̥�ӂ��=��N토�6	0��p�{�6����]�;��b`�V����f!���A?hh;E�粘:�|aa�D-*���e���0��0�Ҁs$*���0�F�
�v=�w��8H�`3��ԗM���u�Y3����%窛���c]��Tq2��d����yP�����9�H�\�l%��z_$�!��+���� ^�"{�1ǿJ�l��4+�{�W�:dF�k;4R����C�d�p͂QR���U.����:��ȉQo!H��K+�$R?.C�w�O�B�ķQB9������u�O�_~�T-�v�ǔ��kP���ڐ�Q�-*ħ�Cy]d�G|M'bX������3���_U�K���U:k'�G8�}��d�z1Q�֗��Q���od��q#h���6/v���:��c���:��?7L�WuC.�����{�1��՗{��[T��U�ͿH߰����kL���9�iV�`�y���g�?��V�xzw�Ǒ=���^�]m-�����1��[ᕲ�Y����G����8��0�/�}Ÿ�k���4�?a�����G���
%���Τ[���֜qS���I2t���~B���p�@���SQ�\x4S8�k��w����%6=�n�A7���Dr��׼eQU�Q,Ǯ��&]��j�i�ɼN7���&�@+Q.�����{�M㔛j|ů�T��}��9�?�`�{�P�%�� ����dg
ŅB`��	f;pX_�߾R�ܓ�v�2� ��q��ě� ���o,�}�E[]`D��&]"�@�e�!����{U��I���:������X!�f�B&��gg��8>>k��N^S�g4Sή�MM=b�3d�C�ڋ6��q�~3����2X��@�ހc&��s��O��q{�?yCi�2[����qPX�6ԓ�I����Cʯ�v[�i�D� �郄�pj�:����S���v�p���
!�����Fg���k��ɰ�������AM2���
V8h��Ϝ��i$+rl�EZ*%ALhz��p��/?�j-���=}ާ�"���#��)9�fxE:x9�{��e��U��=hO��T�3$5������!���!Mi���><����F���%�.pɖ�ڑ��6\eZ'2[�ی;%�}��j�D�iY�%��U�X4�����ǙU����+���[ފ2��������۱��DfgS�h*p:�c�/��>�2*�)�u��{�eA#���