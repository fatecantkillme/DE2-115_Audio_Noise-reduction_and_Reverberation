��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>b��z�P��d�d�g����WG��򈣿ҫ�a���GZs�o��K˖"ƺ�ﺜ�e��$���NdS�L>����k+<7���bY�� �q0���\�aR'H��m�+�r�p��n�NT���,����h%���h+��Z���$�51f���'X�J�)��Uq�fM�rH��	�[&ME��&����hF�Z3ܕ���~�,���l:6Йye"Ɩ�m�I��PѠ�<!Pg-lV�����
��ݖeV���M eC$����!�Ւ�(���y���U���S~�r���xL��T�֌��~�2T�$�*���sp�Q�{9�4��]����\;34�R�\rް�'B/0.�5�=ʇ����.�*x��[ۚ��l�W%��|㱳X��M�ŝ�b�r��Gi�|�y����>��ԃ(|C
�	���g����DQ�X��ԉ��nEgե<qr��"^��4�
��l���ǲm�	������ �#��|z��O�k�&'AV�� aU�J�"���&ە7��%Q��+��cW�s��:1�\�U���4"�y�)�~�����l���O��J$VX�ԇQ�0A�UD\t�*mDط���x�A��Fj?=�`>Nʳ�����f��F覱u�����Ōn��s��w�F!�3�.o�;�ݫ'�Q )��W]�0��<��_t�-����D�S�
0��B���}��9h������g�/(��ȑ�|�8%��ֺ��#o��Lm2V�e�+���U%�ƛ��#/�j��-Vk��%O
X!^�D�y���!�,��]�����i�p]s9Dº�T��$����Ì�(�V��V�Q�K�I@��6
,��1ӭ�1�T����~����	2T�U{ڒ;ajy��M�h[���9ސ�n,��H%_nƬ���x,�Ĳ9B���9<�6'���K�>�@
��^����c��B�Z�fp�zV��T�����>.��m<i�E�+�wZ����a�ړ�%�Ȉ�Uh�j�鶠XU�s�Pɓ���vj�D�z��G�o�v�+����QMY�uN.vH��[PKܲ���9���i�-F#�ThA�s��C~�x���9/�L�E��Ҥ��ۂz�t�g7�7���	ا�/���֕�jl\��[!��(�/��m���^ą������"Ȥ��{�+�.���,(��'�vs�� v��9����d�)�����G��u�I(oD��,o��ZPVcMC��}@�O]h���}fi�@#U�߭A)�d1��\���N�qAK�I��i���H��	�� E�U�qE?т��iwA�˗�<�948z?B�F���nJ�G�/��D�ɋ��6`�p|S&�98�x�����z�KI��4���.b��:/L8=�L��ԥ`G��K.�wr�M�l�(�㓃xa�&<��l�L6��R1��0��A�[��*��������T�s{�x�������12 �*�!�Ў(V@;8J5"K��:`���8z��^��^[�ek���@��J�8'z��yd�)EԆ'�I�{���SȞ����8$BQu��7��~)�;�� �94i�vO\�M������ToÜ���8D,.F��C[і2Go���A�rE���]�0�m�bB���7�J]g�?�_��j��{A��L�O�+�'(���]H�Pތ D(V�L�Q�ęz7���'c�gS���吏Ey.��_�ZY><�Ѭ� 5E��+��	-���tϒ$�٧S,�����6���(P8iJuDE_7�yc�5`qR�B��a:��\���� Oԟjj�I�Nt���L��BBm�P�\�!��8�GR�i��p|.�*��c�ľL!nٴ�e�V�$�#Ե2�F����|	�R�$	T�2Z2�,�S	��&�n�_bg��fݴ�G��)��=�'+Y�C�e��X����z�z봈%��G���)v�40.�s�4���hb$�S���2&-F}��xAd}�5�����P��7�N+Ȍ@M&�m;�f@���<�����@�9�z���|$(k0�Mɚ,S��6�4e��{�#e57�Hg=r�(=	z�=�i�]6��2U�N��$���U<2�P� ��WH�\-U���2�?3�;E�-ƶw�Ø��;	�1�
�����ͧ�Tt�2�gL/��H.�:��G��r�N�u��99�M=��ꨈ�w\��-_݂WغX����v\���0a���j��i3$���Px��
*��x+\�Jȇ�'2��Yuv#Y&Pi:$��0	|&��46��Ⴅ�}���ygX�.���\��7y]��VD�Q�8|V��X%F~��������Թ t���87xe��+i��j�Uq���n��u�VA��Hzt�����}t�ك����t�C�ܿ�U�.��]Tow�wQ��vm�a�8+ 
I���3`nba�+
�1�֨��z8�'Y,�u?����@wa/hi�d����fX�ıs�<�0d����ރ��d����3Y�m�K�R�����{���DA�7�T4޷��}{�������ɱ���[��S��|@핏?��px}w_Y
%�	��y.K�kK��*X�J�����^>�w&'y���U�	�3A���L�����Nћ�����m�Y��'~�-h\0-yY^�S��R��>(dz���Uq�5��;T+Y�ו���Q���x��a�e��cD;u�F��GW��I�ճ����+Vs�����i��6�b����yY�O{e��J1[�Bߒ@m�����ؖ�� Y��Y�pG�3�S�xT��k)z$DJ�1%�&�Ĩ���Fݠ�u������ZFȿeN3����<t���˔TF����D�����h�%�(�B�p��Â�ς�l�'���\@	�M�	4�ȱ���@O��s�Q) ���v�%�nG]�L<�/���������A�$��٘��_�"��������ڽ���ּI��q)���8F�!>�l�߇�T��#�޺����1+��jƎ��s���j�*�}#>7���U��a|�(:2����12��6,e�3f��,�ň�R�Y�7�4��p���>���r]���)d�QW3�++SXG�,��d[�!]�6�!e'.� ���MȰ)�iW���#7O��q�M��cǓfn	�^���Of�?�ٕWI��d�jVӓx5��@2""��7rI����U�j+��MGrC����Ws��r5����ҁ�=ֿrSˤ6�wB�(~~�E7�.���Z慯A�j�'�s�����jq�q/��Oq{�������eȞh1C�Yk���M��ц`����Q�?�ն�Q�7���0b�R��i��y*�3F�J��T�หFw}�K48��-z�8*b�~q���$GaH��#q?	����,X������N>�%�qs[�v)bs��T�vP����&�wC�>�&^.i�A�A"^�!U���V�/����%�!�_ۋ1�J�7|�i5ĨP��P���+������ݣ� ����~S--��:SG^}����}8�m����P��tA�d���Tk?��H��XǇ�nL*^�D�X0��q��)�-��l5�)rH�[��#�k�pAH��6��B����t��ا����5�p�)�f�W褏Uo�^�m��}{�j*%��*��;4��$QB�K�g��&X�D�vu ���T���E�G 靡6w��Ԙ�/���{e�c�J���nT\LmK���G�a��/�۫�d<{�ɝ��u�� �4��2D"}��l'k��o�kI� G:����<�ۂ���ث3h���rTH��=�7���󩼃�N�b�4t~Ϝ?(��7�o�`w�z�J�pL�����y~$Vs����1�S2��w��'郬��^�}k�R�l����=(ýw�c�5�������ؐ�jK
��uP~�����Tۘ@���W��.��<zC��E�g�h-s��I��&yD�ҠB��V�7VD����Gy��/T���_��r2n�8�T�mտ�������� Kb��B�
nXh}4��gV�զ>bo3�'0�o�Jn�-�>�x 1.��*�������H��>u5�#�n�E[�-y����9��	I/Yu	���M�){$u�e�l��؅*�eR���Њ T
�5?�X���l�@�]՗��s@|fi'�,��B�0��#6#,-b���7׶p-��8~�,p//��n�!H��tn��7�#��1x֪	�q�1?��VM+�
�zXb�:��x��WM������D�+F��8Zf/�P����Ѝ���V2���$^Q$oE��X�u$����$�H;+����S����1ލ6as�A':���(t�y-i< ��g�a�*Y2$���d�ۄ&RO{_�����>N1�ZoV|�xH��s��4��N��0s�"�Odٝ0̀�����`�w�+�]�UiF��*�c�$�K
��b>%�� 'h�rut�R�{�U�k	���HUlBEnuk��ל�O�F���p��̆7���	(�Y�.I�o����C����ؚ��� ٠��G���%R�5���������Z�vgO���m�876�
�Kt@����21��n�m�C��hxt�&¾��@��S䔣��%m��e} ^��e�f*�DWߐ�'���l�&�q��A��É�׋���[	]~k�y�[*���<��t+�lm�)60n1�e����5�"�Ɨڿ%Ḯ�K���I�"d�J���Q�o������pX��@hcDVR�9W{vNb���p�]0�E�� g�Y�/�9FqWBʕ�PGI���7J#҈D��}Q��Cw݄�:fg���k_DH A-�Z�)�U|<�d�l4��I�Md��~f�/ξ�[C�ר!6�1φ-�Y���[*��~ޭO!*�s��A�IS$û�T��UN�B����p,O�\|��ɯc��I���}����O�-(��+0k ���A̘0�ݒ�7��.}��ڃ�rtyIK}�2��<Wiرa�KL� �;iq�����=]��@Q���f�<��/�	PE}<�R��D�����}B�+�U*f�f�9[E���eO��9i+�hz�5��X�����@1�����dD}���ŵ��qW �4�k�do�<��x�X$b^����U�h����F�IΫ4_������
�d�9��#�o����:��${|��mt��z�@�I��[�I��0�)?M	M[߶�''�u~�+FM���A�i���C�� = �L
���m4`g  V�HB��)�3}9u���u@����|�ħ����ڝ<�oN��
ؠX�	
�ɲn��'^H��zY�.FE�5�=Y��ׅ"�K�B�v�3��Kj�]�݌Ԟ'�)�<6��s��\h���!�߾��#��0��V�3��o�3����vbKPR��n9�и�'ܱ|:�����Z2��ZRW�-��#��ت��$>���+������$t�$w���(�AT��`7�u��M��	�MOQ}�(���$~^ ��	d�:t��V�§0�q/�_ܖˏ*Z�.��v;]do�Ď��^	�^;>�&���D�-8ɍu�aN����~�?[jX�.+�R\M啤(��3e�c��	ם+��Od����6�?~�fK�#n��9�jy}t,�V��Uj��n�2��/�RP_X�<�l9�M�Ȯ1��$Xl��a�]��Ia���w�n���h�	/�:R��8�//��Z����$���Hw�x2쥇9�bi��-^p��[:;����o#��89;�s�E�)���Ȋ��Q,��پG��֑�3q���9Ic�G��0�3�D�1�T�ل1XOt���2��o�צ�`�<Z�ϛ����ɖv�ĉsW� d+ɨ	����+Ь�����DX�[kz�e/.Z#p��Ɯ�ul��f?U�[��bSx��ro��3C=�̗V�ϰzztˠ��O!Բ��S=�k�ڇQd/ECqM������X�c?��T�
vn�#m�^U�d������<ar����WɋPH���.èA𷹸�s\:�ݲ�4�Ei!"�b�]ҾX��~�8�ѽs���i�\i/��_�?g���&�$i�������@㧣8�.H�����TT�U���Z���<g-�-�K�y��	��=�;��(��&3}1���_��� �2�v�Ã��U�B�凯�w�޵�"��(o�����@�2��їz7R����,P�X���O�����?����Z���M>��<�Z�Ӹ�c����?\)�rYOF�ÿ�y�y��KJ�T�1�nz_�g�^��h���Q�^mCU_�΅�Pas;GmJ��ed�Y�]���