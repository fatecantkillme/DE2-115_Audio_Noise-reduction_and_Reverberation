��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|8���e5�I��d8<��.�l~GjqG�F������ӷi�FՑ�!aX8l��s=I�* �3J��y/��D�)�}�űv���D*�_a?��!L2�nN�L�4(�p�-��M�h�B�~f/�S����@�������cpd�+q���:`�D1�~�$�4[?�� mp��w疶�T�R؎�ޕ���"D�b�X�Ha��ʕF����l��7YY�*����� �:�/9%����A!�(?��{#�d����Z��>&r<~O�ks]$�r7"U��u�Ķ��������[%7��Ӿ��),.e���;�aoS��g0�C���l,�z��eN��-���e6��5kt���G�3�I��7ͽ#ͫz%nt'C�J��0'������6a�M��H�o5�g�|%����P��b�yQ��H� �+4�ʠ1^�v#5���ɻ����4j[o����V�%��[�m�R�V^���@_-� �]Յ
xe"Ha�{n����m now rB߯��7y���-�I��
2>Q88��VRo�Ɏ����}����K>F��
�
�1<�Y��IaV����WUPA����&
��,�;�1JV�Z�L�a��u�$�#P
@7��jg������(.���H?"��˩jLCexs+�����Ir�Etb�� f���l�˻vӟ�����\ԫ���Ȏ���q[��*��Ī�wG�x�I!P@�!6��
���C�W��aXci��u3���Z��0u|��#������x	I�Y�A�9{PU1Ȅ#ݙ+ޒ�����uWe�_�'n�Im³�B�F;6� �U�F&�=���d�h�#�%���L��UTZZ`�=r#��ıbLn�X���q�]��r�]��J�1ʳ@�]��7���*�[N�ق
w�U�Tc�Pʟ�L3Sm�[�*{��k�M�5�x�0�l�����̾�l\��q/''Z��6g]0�^r)}�>d��q܇Ϋ��lj��TD}�/�X:�Q;�ixOj�E�������4�����g��6������5�Y�TA�aN�}e'�%���M�0���PJJV�7ŀ�ة�:<����X�N�5���8��I�_� sޮ�L��A��u���Rl.&��4Iŷ��Ы��E��u�.�9��'^F-�3p8��];/��VGZ]�GO��R9�j16�����5<.����TrKC	�v����̑�b�����(�%E�-�Wx����>����P��V~!Ɋ�2(KHʗ���"6!�
U�0���/'���p�V�4EA�/�򓤪r�F�:ˆ�_�m΂���̱�J��Я��F~�]AK$�.�Nݭ(D�{t�(	@� �1��u�(E|�;�������q ����L�K��N ̊�{�ۋq��Zn	���-�]S�X���kS�C)XF�#�u�8yl��������;h�	r��a�v]�<�e���ACjm%�G�ߠ��|d���)�})��z��p���_���Mh��-�^�Z3߆X�:E�<"�xP �V�.B=�0��Y�N�FԸ=]ܚFz��li[ℿ�D�k��5���9y���ˁ���
MJq�t���/)��_�����P>8Ι����������b�U(�P3eO��1��|a���(k�-��J��0��	����v%��w���=��������%��[jA�o���D�N�77��{(��b�g��_�m�]�%�=�,�IVT!x�I�0�<�R�Ĝ��	,� ���	�)�	u��.�d�CKl#�W�31T3+� >�=�Kj���d�'�H�Z~�FB|�M������޽���q�l)֛��G96/��V{�)�/ڦ9=ޙΉ2�z��4=Ӥ#ݠ[��9��3҈�j�ЄУ�O�6�V��z<�(%��)W#�\��à�:$7:��P����� �wT��+��g��Mw��mo����2��#�P��=$� 1l_zb~\�<�-1��o=X$i_O�Z�>%F6��Aw�N�G�ې��f��B������p��g�� =n�P	��3yf^Nٕ�"�8��]zYܻ�����{ ��5쬄lm����	Hhd K�"��E�ZwC��
�#xo����/e��?ė`�x��#)�D�a��=C�!&� ڄ�D���Sm ��VJ-Mз�
r^�	��r@����SCٯ���լ�N�ˑj�X��ｃ�<2m	pp�c�&�5cc9��e�*�v�
ѿĠ$�Pk�E�x?�E�x�vJT���y��"7o�g�Mh)�HK	��/!�o?���#�3BN~w@T,-�:�3������-Ց�Ξ�e�C�!�߳���{���麪^}g��M`gA�n�̻�; �/��(E��U��*��;3�/���)��Ag]D{���Џ"T��	4��<9��hiSZ+Y;�gJ�̲�歱�	���W莎�.r�1�Y|W�7D"��=�*�D��5��vx����I�|a�bI�n����J���$ �R�2W�=���<�.�BH�Rwv$Wۤ` FFb��|���ՔI��Q���"�C���D"�Չ������I�"NN��.�$H�3�Y���M/�v�S�>���j�Z�3k��3R�D�4���H���'%TfC����`%'epꏏ�V	o�"�؞w-�����-��)����D�� %�ţ7,O����^G�m�\`��y��P�x����M�r��`R��JLy0�-t'H��ڥб{j�r.���/����7�&��d���qb��f��Y�IY����x <zu�~C^�Sе2I'�ne��A�F)�*�.7�0>��MB��/fJ�79�bv���)����Ћ$�I��x�N���e��U�
�^1p�{yP�����E���G}��{�7q�EQg8��o�X�$9��l�O<f�mA��V����[XD�WF��P�+|�:&HP�2��*5��T��ΣT�5��Ɋ�3v���qe�R�����i��`S��)�<�WC2��^�kwc|�� X[~̊�܀�"^,��M����1�YX��FxdI�q���R��`N�@�? ~j���	JSU(c^���%?�,��-��C��>����nN�K'\i���I��Q��p�ӯ�|���N��,�����\�w��l�&�@�\�f.smu�!ǌ�>�%d���k̢Xg�08�S�w�܀�RT��#���Xy|�3J�H���RQ��N�\H��_&ɵ�/��d���P7�O�?�B-~�^����8���)������?��a��K�ۆ�����~>r�Q O�h.������Ř�	�PY`����J��������f��-.�Ha��������Ph\�hW�>!��)�gլ���Q��U� ����u��Wf3�^%�÷�g�w;���$x����/����!d��Qn$\�%���NF�7��T�r�>�/��B��2���|�T;֊���������#[mc�ΪN):��g^�HGb�Ɛ��)��5�F����m�)Na��o��se��@�C�4���
�M%�c���E�̩��H�Y|,�
��p��rٹrc����<��T���$"�ؔJ�\)kkM�L0$��>����y���4n�d�`{�n�C4ͭ�<�y:7�N)�h��	��2W��Cx�[��Z�0��9|~��Û��kk��DR���*�ƥ@r�|�߭�t	m%���zh�4��-Д��+3K�K��:m˳��q�%B�`�5��|���������'P�g��"�Z��U�h�O�5X�(���G�-�E,�?DȶZH�-<Wuj�p��AH����(�P�X�����E)�����
�+�?��x�V6dk�
VbP ِfd��ڪ��)�&�SIR7B�;�w������[6F�()8&h��������5.B�މ�`�]{�X���J����T��Z- 6�Q	�=a����	���zc�<�tܝ����|�c{l�*%ZBH�-^E	R؏��s?���+o��� p�jɚ=�`�vJC�_����D�����o�c|����W?ƻUN��,�R�����S���%��t�*������g�͏|��S��t|$~q,�E�}A���(��8�\��
��q��'K���&< O$��:�"2/x;?1�x@s��4�Zp���'`����k�G��V��5ȊC�D!5���o� ��7R~��+���e�U�$,����{�*FR��>�7���O�k�0MN��j�\��]���������X}�I��y��h�b�[$�P;s	��q��e��~0�jK�]8m���/J����竒 �?4�]���72�ʏ<J�EظQd�|H�� �����t�
-"w�ѡ�I���XL� ���k���!����P�1*~̋-�7���v��,]^�﹌�m����ZWFw�����}�]OFA����Z�T.��[�x*���2�/�n'0�e��vȨ�Я©��)�7h�g� �L�6x4�
����x_�=2�~s�v��9r����c�q��L���.��*l^3(����D�}�j������6�����3�GN�����ӱ͖<�,�^���s�~��t�V�W�=P�`h����`M�a�xq9��m�8^�^]�:~2 �6�b<�N*ڀRb+���S�S'Lţ��I��:��Ȭ<�o��F7�z�1`d��4Y�����+$H~��M�����V�4G��;
� ���h��`k&�Y�h&,�4�q��dY�՚���|yYZ���Mc������o�z��D��a㾝���.S���MZ(��&b24��"���	�0i��t�y�(�VY�f�u`9�]?P�����<^�ZZ�2zipH�[؈c�&_�ˊ�;A�� ap�5����G	b��M�<��Ӷ�Ϳ��+��K���w���8,7��eׄ�
G�V��$�_��z[	�)",sU˭W�˴�BS��
��,�����k)�.[	�� @��ጀk��"���m��L[�di�a�	�ԝ��2h6���=��Ɵ��G���!�Ԗ����-̕U�#�/_b�V���4
1Wi��逪�e,v'v�J��g�����Zs_c#��]�R�i����>��ڞ���-��%����2�RԚ��}�ߖ\���>c6*�T�,��w��Æ4��񁣄���2Ӵ�2MPZ�PW����_���|\�:2�݇'3T�
��n���M���:���[��Z�M����$>�_d[�=M�$Y��6��l콙� B��6�J�F��߾r:i�5+�:$p���;�T�"�c��N�k�@�<.�v�0�t��WI�6�C�bzd��b\��.�J��'^1�6��8���7zˁq�0�t���.M}][��yJ�T��8b���^�j�l/e��(��o�31�h"=�}0��:)m�
�[X�L��Dx�d��PBU�M5ȯ��?i�ٺv��!>�`}.,	��#�}O�:P
����NL��F-��`�=�k�i�����O���]!K�ÿFFj��Y�g<W�mc��I=�d�y�b�F�:F�ΏA�����s���8:����7��]���#=��9P���>?��(x�>m ��~�d���Py�9�&я��^K�|w8�E�`�`�w�@+��#����ow���#r�ɏoQG�Sg-�"�}[��Ŀ+����a��L�E�]S��������Ϥ�Y�{I(r�?̚���t�0lv~\ٹnך������FC���̑��l%���q�F%y���v���"����F�s�sfb��o����%�j��s�����e�YF���$a��11��H����8�8��h���R6]�H7�F;����ˑB�瑱OQ����漛����2)"�k�b���E�����,��9X_�S�'|pT�� �d��UtP�󶆥vy�ئ&����ԯ�2�UIU)a�U$+zR�QT���h��7/>�U}uW�fF�������J0w8�My��r��Sj^t� ��v=.!�+���"�c�3~č��X��������rTO��	�Q/T:J�ǘ�sZ
1Ȯh@�P�p:��|��y#b��Ck<\�*L��gD�z�xbf/�F][�)eN*�b7+�Y�x�ѥ�����E[��#���C
UF豭�
߶������&�*����R���Ć�P�����#��1�y9qkثZu��4���MS�� XٯJ�9!ӝ�������h��O-�~؇OǙ�}AK����_iku�4�Y xo}��m_Ɲ�I�A% m ������֬v�%b�0
:<9y5� ��`�qmH7��1؜����M��?����P��W��?nDO<�X����
"��'_L:.`yLfS�^��t���^9�������l��{%��cO�Q+{!��[��=�f�9�SrQ71����e��o��&��Z����.�TڸT���Ntt2&(W�˗�%)�Pv��AL�Dׇ��p�1Mm�T�+{#��o�
W?�C
���d�*�[SĤE|��a���\���a�l=�T�E�^��}�dq�`[L�N��t��iC����/AR�!�%�kSk,��=#�Ԋ��(lNN/Ĩ��h�\�U'��(K .ڦ�3��r��_�"�"��\#��h�_������]�f���'�|�Q��uV���Nˬ��1U�P��%��ͩ�ʽ:����VT�>��]�䗟j��k�Q���(�\� ���ݰ:u�l �e�TG	#� 1S���l�Cӯ���
Z�uJ��+��s
n
�;�vc]S\�Y[}���3�V�^}S�����iIa��J���D^�^�8Y�5�<;��
]YQK!�[1 ��K�%�l�1��{Z�Pzܡ���g�SyY� �nA�G�T��.P���&F��a�6�w.'�lw�}!ъ�ѷ~d�����׌��&� V�����~D�5�֓���B�O.�(jOn����+4\���Y��ۜ��4����g��E���W�W�(f�OT0�� �>B�� ��ri8i�jg"
P!����Q2�Mg��w�p��	N(�Ţ&w�tTF]|�uQ_���'V��}��_j���K
�Y�>�Gɓ�Ի�H��kFd��͢�U�ă#������K�16ϕ��xQ|dۼbE
�����H�%?�/E;^��v}ؤ�k��>x�Q��Z�ap:<��9��;� ������߻�)�TN�����,�r���;{Z+H�ҩm����4��oA��<t��O�����;4_�@}~ћ���t�0Tϖ4�� ,%�ۈ��%�����Eu�6�h꘵ �^J i�D���!�~�(eI��&�l:���'*��k4�4i�E[�d���&5���yۍr�(��L#�R�yV���|�EP
��z�,+�<��M5y*z��Z�����4��sD@�.,��e�� 2�T54\��`F\~��9�1R��K�{�<�9Qݲ��;��3mb���f�I�+������ʷT�S[a �j��!鏟��uV���-W�*�����6��
�Ef�k�bs��ɭ�0���6!�"	��p/y���$��-�bQ�(g�*e�쾺�J.aۃ|sC����(� EY�+���x'�i�>-xF��`͵u�D=����.�-��	��/��l���G,`��H�*H4��4������^�<﫮d�I��1��F(e��^cw�?�Fa���oV��Oe�wON��h��M��	�=XIs	��CT�%=�#�d������C�T�"�7����G�����ӬI���q���P-1g��������j�x�P B�$�v�J=�}�{�� �aH�����(F�cfB�?4V��|���c�%]�K�2�5bhZ��oP���B����wS�o��h�[m��l��D�Zy�����~4;�:���g)$��VT���M��^Y�a1�`i�������ܢa�M�^����E� ��������M�&d�p�b�1#U���@����JV��j�l�W _���.�!��G�8S2� ���M)'�j-�h����BqtdZ�yV���0�9k�g��n����S����_�V��2�k��vC�@���'Eu~CY~g۔�j[�+�I�^i+���%2ko3]� ���l|Qa<]��m��7�@����*0�[ЌT��u$a�_8�A[ ��RY=�-�������K	�/���`7�3�Bcs�^�k/�5z�M~��*r���U���R��Ҋ���ω��Iq��� ��D�j!��%�֗�gEBB5	=��yB'�7+��1\\�VO/��_���q��F���q�����wv��@8��CF�V"�"�oI T�r�δ�i3��\�Z��_�i��Z'���'fM-S�e���΁����GA��	���f�R���{��Z���-;�;���v&9�'��UQ����[�o
�_R�xG��U�ǜ+Ô��[M=�+zSY�}ꫫ,7���MWgکy�������R��1_��1y��Rޘ���ZJ����_THa��j	�=�������K��I�`h��2� ����?*)A�Д�����nʰr�g�����H85��_8%W�ݤ�̓" ���W1�G��,�*��L��.���C����0�
둪����'��7M�|Δ�\lpB{#TgF�M��.ޚ�B���h��a����W�{`�V�:��-h�B��O����������x/�.o�Z�Y�_F۲��e/��k�8���4| Gפ�}��Bb�A5�oT-Y{N�A|63��54W�w�70�*��@��	/@�����l�Ż�Ĝ����M�Y�H�"�;��L�_�b��JC��6���$e��Fײ
^�4�8�윚J?�L�������}������Z{�&!H�B%�X|���FI?`ت��ʩy��^�De�7AOB([zC�<i���c�L��0������k�����?WOM�Z��ye	��u�,��Zo��v�������̮&��˥t�t�u����f�>�3��Ћ��Ͻ��%¤Na�=�T1QG�7�E䎃�*��<�4�,?t��ʪ����WΔ;�g���<6)ls��@��X����#���N�|Bx%��ð���k݆ͩ�>L�a7�2I�����q���$��d#(��C<(63���4������g�fd�ʹM��Yk��4MS�>�L;E��������gl<��|����t��>����nD2�h��?���儫�{���������vb�b��f�x�Q}/)0����0y M"����y2�<^J����=��H���Mq����}�+oy����5%(}q��Yطvoc�g�ӽ��ܪ�gi��eu�ƃ��hi�B��ѲJ`/��~�	�i3�ނ��y������"��̣(�k� �`(g���+4��� ���r'��u̴>s�(�[K&��8Ƅ)�Q1"8�U]@d�����
�_��s���e����z ��"L|���:>{����a��^u���_��#,�5���k��t�;G��܍�=)�B���6���@N��]ڶ�iO}\�I�풫�l	p���z����v���!��p�/.� �1>�YItc&��<��6�L��;+ӝ�4��)u��� 苮,B&PyyҾ�FKm6:7�*�drk�;������QQR:�WME�L���c|���4��v��0)!�H��>Mm����ɣE� v�Cc����;�J��@Tu�8)iC�2��Ќ�z�5�!}�;�N�ӆ�@�9��M�	�U�/�����e1Mx���pKG �1%�d��
��tY��[��eݻj�y_ȫ��@)�`�4��Uh!6�ʺ� `�w(-S�>�n��y3NpjHbnn|/�h�1/�ܻ����H��7Q�c�{�1H (�Q=.�+����E3��H~����\�F�"U�{��SH�Z�����S˂_Ͱ�E&w����sxw��YG��w>��꣒?�z��?uOi%���*��#1:]9��K��\l(h�ɹf��P������og�\	�=eji���W��vL�7 � �}ԑ	Z�q~B�k�~�1��Rg�M{A<9��2�E�Y�yY�U�fp���'۔Տ��2�p���&�k�t ���v�3��}�+
'��_;�HKI-��ZN� ]��U>��������cMR!L{�f�cH�QKhă�퐋���	U�hü�VхQeg@g�$��_KQ4��./���r|�Z�i캂H΂C_bD����p��~_��\mCqiO�T�oQ@LeM�[)�$�.��/� Y�3�(�� ���V7A%�6@�4XEx�k�FTO0n�暺.#�Ww�� �Xm;*(����!���sI[N�Khf?Y`�*��G���ϝEɸ(�k���2��Em^&p�fi&\Gf�9�Z+�E�0�Ӟu���pͺ.�v��p��܊ϸvS5*\�'�b�|��ɨ����B�זyp�M�Z�1�;d�(��}�	2OK\H��?�i���{
z�a�����z�қ��	�{���e�0�f�/�W`B�ݍ(��:��x`�Z���4�k��ծ8��.�����6���C������@�k��-��R+�E���iڡ:Vx�0�^|���ѣ�Z�^! �W��.�	o8j�;U4M�όZ9Ll�\F�l�f� �W��x�="��ξ��S"N�֘����șW�@L�v3ܨ�|��u[Y�kQ �g���&�.�Ћ�.���0-.���\S�F���vu���k��ܞ���Hĺ�� �����WcS��'�5E�hX�^�C�Ǜ=����CIu��>;� K5��y�*��J
�)��y����Ц��P�`"x�1�.���`�Ҡ�Lޘ}��
a��c��V>H_�R|�n��10 #�߭d��&�����be��v�C

�ÍQ)�|zk���s��uP�W��l�れ���.@_���?���pe����4��<�aX�phuF=��$f뽰��-�5�ߖ۵H6DV���`��?�F.�YcdT �B��S�n���5�T��p�(8~ೄm�h��Dǌ�\mq�eFK'�u�1��&��k�K�4d���IQ��I�X����2U �>#� ���
�g�"V�kvr\6�W����8,5�J47(�#NyI�>0�g��4~k�B����g̪UX�w�S�J�D��8��V���o"d݁�EzDY=�?�H����)Us(��4E���@���I0�IP��9t��#�Д�Rg��sO���h������$���{�=��Q�ITɐ�HVaF�+�'���E��&�ZXRҸ���3V��{"Ƹs����
a	2�wi�Z���^�V��m����}�E*�D?x0���F�gRH�A�sy�.��ǀ����y1Q[֗���n:��V���iK}@�C��K������ГVa��Q2O�%�8���"�[�%7�z���>Hȓ:��aC����q_qy�����B������&L�t A<�Uf�ߜT�L���`����l��p�[�wvb�f<SÈ��?󽺴�5kq�>��G���b$fa��æ�#�j�z9U�Ӧ$o�L�����W/�&V��'�@�>�C3rw~b_K�h�C�}.l�65�H���4wCj9!ݿ���9�Y#�#n�	��dH�pZ�ݗ�[$Eհ΢/�>H�q�ώ�O|d>u(��:�Y��X�Q���Q�˞j�D;v���򡁆2˘���q"_Cu*K_��V��f�~ļ���,�;z-��b��ͯ1;Qjs�mgWm�xt��_�_�F=�+�^�����ĩ��ۄxIbHk���y8��N6������"#d�Um	�w�ݚ��}Ί�I���0$8G�q���'��+)t���k(t�	I��'R�#kIŵ+�6�I!�K�p��A-A @C6�7����=%�ڏd�������~AQ�s����WaNۏ��W���`s׽�ZF��@lQ97O����փ}���l�*mh� ?�P�B��v���p�]�tp�eg����"�+��r�n���R���}ӹw&2�e��숢�h�&xRT���뎝��(#�Ta�� ��lh��W�U��:
6�ՠ�7c���晒�5�*z4��w�@�n��jjB#H�L�?�o�I�]�k�e��ոMs�ěT�NI�����K�{S>����j��O/*貎� ��RA!��!׸�?��0tGxN�2�l��vJcK��i�_䍥0oת��
�,U�V4}�*� ԗf�P�XT3)&//לb{7�6����"FJ�e̽�����%����{�~ݫV���$:F�鬵���Ұ*�/�{]�Q5K�;"J��܆}Ű����dW��>b=3�E��u�菱�J�����6ӝ��xWz>�����Lį\ȅz��h'�;t��������¸Y�R�)^�"h�R�O��_��c���lt���߿���b������4�Ql��"xڕ�I��j���4/�-����V�����J�Kv�=ؼ�+���#�ovE\�8`�d�o��.	��G�ug֞$ui$x`[�����D1�W�؍��5u�R�����l�]�GU���C�G9O1�	9Y��+�z6,ᱭ�m^�pKZ���� ���0��^�{t�2* ��Q\"H	��t"��~��!�v
2:{:��K�v�k����;�v	�?d����d�H��4,Qt�ݳΈ�%��𒻝X���V�g��tp��o��o�gP�ОVsݺ51�&��r�Us_U�a�������$6)
Y"�D#}4����Z����D>ٕ"��� $ufݒ�`7�Z�/���U�[�g�7�Y�&-�@��KZX��^�re:S�!��T���ۮ{�F�e3���
#b��2V���Y;~c����fH%V�ܕ�T�J)���+��O	�����h�hH+'����Uv�����`g�}�-��Ń���'��`>
Uـ@�}}"P�?$rsF�o4����6zDpF��(F33�#�=����P�b�\�@P(?�'ӹ��֢�vV�k�z׺��kM9q �����Md�	��>����$ڛ @����0	!eұB�oR4A��:�ǚ�Ⱦbz���AHbu+�����7<��!)�����Su{��R�0f��B�uzK2�ʾ�I=x���A��A����VZ=������d��*}ӞN&x�p&Zx�U�C~3].q/(v�.�jv���Q���b(Գ��'���W�Gn:�<���aiž���LI{$'��Y}��$�_�i�i�Ҿ�rb��K֍���h5�׹.����A������	��.�<���Kֆ������~�?��Ȅ�YCWi�&-�P�ܙ�;u��o�IHf���`�k�tD�	akU���>Й��p���.d���Rb=����b_�l�fM4#�	ĽhzI���_I������� ���D�S�4U}.[���?����D��Ӯ�)w=�t1���CJ�^{e�,~��_��ͦ� ��p �d�n=-�2�]sW1�S��j=;�cw,�������&�������^7=�2��n�ːwإ��u��b� ��E�92���~nK0a���S��RZv7�$ORU8�}E�j�ڡ J��K�����>��iA*l��7�24�� m�گ����Qj�P��#f:�T�+eDٶ�÷���u'`����#vԌ�t"68�������w��Kh@��ؗ�{J����$]=4o�	P�n��q���m�������ݶU]�hǂS��%��A��c�0/�"�~Ȋ�ѭ#*��0q`�R��,�fߥ�:���e�h�����䜇���5�̾��o�5�\��_�E��}z\��{@���\��k͹p��G�����	�C�Ć^1��!xF�Y���	.��ޜՠ���S�O��>h�܍�9��u�̐{��\j�n�+	k��I�Ƚ c�~<��Um��P�ފ�������A�%��O�Kv�@o�^��M�����G�ƴ-i�T������������V�4즋=�v�+Ꮝ�t\�+?/N6m�`�g�,�'��g�އ?��Y+:���ԭT� �����
e[���׆�m����=�p*W�7��k��Ǌ,���Rn���2�t]���*ȗ���d&[�P�U��.p�s��}��p�8F\6�$��7w!@��%��۵0�C�����[,*U7U�~1ņ�����0{��<��S�4e�����ܔ�~ү��NC/_����cku�ѥy�nnW����e���@2�Ĵ�N:(�G���J�~�#m����:(���j�����SWI��֑kqm؃�5^Q(!,t֡{1v*,wV6Gq2x�!�xY>`�����&<=��`f�r�'��L ϒ���S��G]�:��Ѣg�~��Q 7~.X�y��ί~]*:������asY6��-�~��:��C5+����t͢c5T4����=�:�k:mI�e~8�LAQJ�2.�yz���|��4�Lw&ETT2��Jӑ��)�� �]%IX���������g/
�VݯhI��2�#�v�:]	��ˢք0�-O��$F�>�l����\��&��&��><����[�Xk�C��TJId%��t��|���%�ϟ�Y%X}^��0R�.�6�GI{�̐����پZ�T�~P��(yf٣
'�LI��]��y�B�~��iT���Ies�1ļ��[�]V#8���	[���㸿���E��ĕ~�o��<�l
a_,�}��m>�
��';tN;�)��O'>��	#7�|Z�5�ΦS�h���,L�ؽ�t8�ʕ�MF�/V}(ԆW}����j����d]�\�x��$��eL�	���7 t w ���,�2/��(����xS� �GEd�λ��%��A�1~�Gj�z[�i�/-� `7�Q�(�s���y2��Cr��%��7�3���3{d\%�h��)5�^k�.�O%�7W�Jߍyy(��&a���������!�¡�\��KX/�]rx>5�\5hD�2�z'˭?��й8����0�n�k>�6��l��״��Q�hL����jez���f+�
 8��7����(�ɸ���e��
��9g|���2��/śhTae��f�z�	w��#�mM���nȋZAKMnM{�rp��b�����a�'8��!s�3^-X9]���i�Bj:U�V��x���>�~��z=r�Q܁�y��(�O�\纻�e��%�6dJ3��<f��T��ĸ����d�	�E8���P}���ZJ�N�bx��{���7��l�^�����[4�l�9	XDp"�l�.��r:c�/M�N�]G>�ww�*�8��$E�FFԥ�de���p��4�d;�4�z�IV+$�������=XI�[�:��¹��tW��Rj����柠4
����lZ�W�>{Dk=Tp|2Q�����'�e���T�G�o�0�7	Ds��@H��,�Ϩb�ST���>�r��=-�=݂��~;��:Ńh*�?�@7���4lؐA�FE�=�dX��La�%� J��fy2 ��?�|��l�x��xL�b�PPP�|@�Cх���S�}����D<�)��6}�/�>��KT��"9G�Z���0��$��N��^�^<�g�4��S��}s�5A��+�q	����W��\s�gE�g�8N�׼��l<�&cHZ�\���s,tD���P%�%�s�ŴΜ�8���*]���q�U�NS���"ۻYPj�
��
�].E�4����c�Z�>&���Y�4㨦�|��k�{S�n��m��pZ���|�RW���N�t�����vO���V|Sә��\�L��K�j����UԒ'��k�D|�G��w=�Y\Gڗ>˳Ol�7��YH�⅚��T��G�ܪM�I��i�da���qż=�����9�4���-��!� =J�����˟�OıJ2��<�<���4&�g[}i����1bϑ��>IkXr�D�b�����L����h��G��|�02 �� W��kK!RN���*��)q��F�����Ѱ��>k�{l.�O��f��i�>.|H8I�j�e�a�70���JT�˔U��(��?�;�Uˑ�m6ߎ�yjd�S�je���h�WE��m�8���&�o9�I�~x/D&��u9�����4wA�A�q��g�r����ݖf��9&(9��%{M��t(˨)�M����ٜR�44i�(�3��5��(_�ʚ�4�E�6�1��E���ޠV �����ɤM��ĺ�Wf�ȍKJ&�	�Sy�Mu�?�H�C������B�y�)J��,j����71j��HhG&	{�.�U�������*��Zw��@��������u�l��2�⃩g%��ks|�\a�2,7ش��~xa�����}Pk<l����^��"�1��kBy�^,���R�h�y����%�wE�1-:�	oyL3 ʸ>iu���C��X�{+Gĸ�1+��YZ�n{F��0z�A�4�9,)�3uЌ���J���U�����UmR]��آp���lw���\�n���45��7��k��R&KDM��'�j�gJ�����r� X�bz��Zq� )c�ά�����߁��r�Q�y�ո�>q�J�
�����Y����d��Q�rj=L��_����7G]+��f��F�b�v�^V"g��i�U8�Hf8f�tA�]]�v{h\�im���v���#��m�o�4�(���i�����q�.�n��N )�y:�a3
\Ȅo�tv����3/HN�߿�h��b��_�j�	�HH��"�`�.�&��A����pE�0HSX�]r[��%��vFv�W�Ვec1�b��5(G��,�4��a̴u�B)�d�v��H�,B7���d�#}L~O�B�։j�r�5��ۋ3-�i�?�M������:K�#�Z��g��$SH��;����sn��m�52E	e.��,7��R@�i�	��=���ěz�c,g�����
̀�bTu���ջ�� ?�����1ؔ���C���A�|<u�o��u��\��r�|�e~�����*�eCY��T��z�Υ�/�=,F�`�v��@���+սH��>�pP��#��Z%8�CYr�����ȅgt���<?�>G��),� 3ƮCT'��,���J
37�殙w�Z��B�G�e��mn�d`:g�LS�����^Ƅ���k��nT���*��C�e��B-baT喇Y��S�gv<VL�+�%��͕��R�<+���X\לR�P<-J��9V�Sy�V���~���7�!�	�8��n��ұP�������&4��x����<������[Tٵ�W�e��4��Bm��қ��.R��0�Ǖ��޿6LCѴ"^��{��7�{;�u��x��Ûy�j�Oh�KT,�������P��ڵg��b����J���V���O���"w8r�%e�$�4�'����
�d��H�w�k���&��i^-5�U�ځ��;j�L�4�^����J�v�����d�`����L��;�=�-z�Pn	�Z|�>��;vo���=���s��+Ɗ|j1b�'�1�ɑ��	yO#���t�����z��t)~\���U+����PCQ;��b_K�z)m��Չ�u�u���+���BFd,7�4�1/{�n�j7�Da�&}��f�M3:�E9u��yL���a@#�h e���gq�9R�6�hxk��ӥ�xY���Џr�@�y���Y����=4gX���������Ew
A�U3�*��׺V�i��u�	o	�p��ѩ	 g$m���B8��)qw�E������$�|���ӋR]�v�ƝY~yIO�4%p-E�Ǚ�-[
5��y��L?���t�2� �kD�|���A�Ӛ-�;a����hQf1�\XT;���s(� �t���ֆiuY=�"ư?� �5wc���`�[?��r�	e>�x������U���o�Y��&젙#:�6�+������9�������$��@��� P�Uñ<�L��y� i���4|�����k6�|����t�}��["Z��D��6=2jy����
���/�_"�$,�VI�B�v6%i�0��J(����Cu$�S '�.���x^�O7M�Y�ג(Ģq[��e��g���'Q��|��n]�n��W\�����M�����cGU���Qr���[T�>tu�"R�LI�q� N���Ɗ�A��)���6�9�n�!��x���|4U������� �ǁAE����eY��w��x_޴�լ�(�4v�Y}�Nc�
���Y��cMA-�D���WT��y$���?���`����w�������T�\zɽ��A����?6��ϧ*WGmy9� iB��AJr����8���&�N�P �����Q�>�i0��ΥB�^w��q�<i2�������pLFȣ(��U����JV�e�L"d��[6�\�C.RT2���H��v�ؒI�G=9�Y{�*?��.6�W�n�D^�u��TJ�Kj3�5�ns�V���8�9>%��]�^�Z��@��q�q{���/x@�.;,)v��5C�!r�cl1��j����;����¼n�ʭ�\a�>˷IB#o���|����W�PU5�*�≜?A�Ws��I�Â{���s*Sg:��)f���/�,X��O�mΕ���ã���]p���Ӎ�[?W�97H^c5Iʥ�)2W�2fo� �O��q���f䶹HK�; I��25��:��>w�j���q7�8�_�i�w�Qn�oC�Z>,�?�o��@��m������=�V�}R]xwR�LL'aG�Yg8�WA����2}�yn����ƀ�����K]�٩�;�T�N�nJ4|Ü�0��"h�J��y�G�*c3�9��ʔe����RxH�.}�ը�t�ћ~��(�J��l��P���h>�Ĭ$m@i���E�;P}�eMl:�y��_�)7��ڝ��o�/r?�&��a��`v�c������z����Yd9�?W
!�> y��
9w�1��� i��A.�I�p�7���6)&qٽA/o.��
���`q7QW��󀽿c�3*���	1���8���p}�2��??�Z H�ģF�,c��^	1�Z���ygy����@�f�����+���%?Hn-�90�L����
��)@Et��%�^�Na0�~�@I�i�\�b�OV8���z3�U��Q�x�=�����G-��K|��8P�Y��u�������D���eNd>O ���\��bƸ��
2�#@�p�KA��]�M�ԭ���(�cH� '�������S's��<\�z�!|��B��#�_�_�d�e�m|���?�6h�{�p�R�h���P�2=iqQ$V��A%L̓��dV�-���Jg վ,��~[�8�2�6��C��5gn�z�|tJz'sHO��
Cȟ���I��j*y�i�I���t�V!SH��Z��W�C���?�/�z�֍����(�40�*dC��Q㻻�km��D�^N��+�W�BF��_����jz���yL8Q�4;�`�'2��'w������!ܨф��O��>�+�R*P]~�8�.���a��L����/�ƊϬ��0�@z�ǅ�Oc�T��Pė�/ҾɎ>-�	+�V�am�v�]
��|if�{���3�V��x�-�:�%&�a���j���bUQA�wZx���j����e�#���n��;��p�u��~��Z�\��t�4=�B���_bަʰȻ4"��D�Gة��"GH2{�'���8lIZ�u�L����%C�^��o�d�"���Ti��#�&��JO���*��	�4�m�-��������IR������������@�( Ĺ�|0���NW�J�%�1A<��8�՚�����Vz\k���m���jW��\W� #���KI΀x��?�!���5���%��h��k	8�	�2������y���2����ko�~
 �jqz�;98��&\f��Ct�����D �ҘB��-�Z��@V��R�ji��;�#IO�y#tVϳ�����va���w˷�8F�,�lsl�~1*e╼t@z }ބ��ڄ�B�U�ơ�7��K$�X��2� �[��	�q���r�G_¦�͙P�lՠl������Z) �e7[����Y:� ֗Xh���끨�`�o" ��%��,R�Ȗ+��kJ�Ӧj��H؊�y�}ƍ�HKI.j���=9�*\�^���w�<o�G`a4DG���m�j��4"\[�o�\�c��Ïؾ���T������K�cH�^
��H��y��ѭ}�.��B��C��=5U�Y�A�g������<�X�1�C�0z��_�(8ƀU��i�U�͎�u�P�}D�?l/Lø�T:�f̔��1/��/�ڧaEݼ�:䝧a7\��)=F4Q���w!ߪv�rn!�@2�K��Ώ[�}6:u�9N�����NoG#)����H��8����� �#mî{N���𷕨�\��Zب��h�k��?S���ȸ�!膽&�T��Y	��x,|��H��O�\���j�Z���̯���A��#o�����hhI��1l:V|q��8�[�s�Qq�Eu�vGY�u�aFk�t���@`o�O������̽&,k�����~B9֭8��U�ǌ�"o��EZ�rW.L� ��[%��3|��:N/��^z�+ q�"��e2	���p��A��gw���>69K�M�0�\R�!��p���9R�$�l�G�,`9٬2�Z'ح+=`ѣ��<�E|���^6pX����P�OÍ����/�/:^�Bvr��K��JO�j(�'\E��dX�an�����H�~�!�5*Δ*�g�q�!ϋy�i�m�Ո���62S;�A��Fcb�&bU!�Jڄ�j�_��Y�!}CcM����!w����9�K�j�sj�B�� K�'x�<�Y]��<�)� 5����[|�K���_�ŽLU]П�1�;#Vb��#o�4��Y����v��s�ڶ�*��K]R?Ȁ�(����%v���0a�K)V���9倥�E�>^J@L�@�cKmf�s�"��b�+JD�n�p_K�<C%#8y���t�H��+,j�Ŕ��P��[�Pur�L��LS�!UY{d�NI������k7����VЏ6�ZA3cPBP��#n����ȴScLw4]�1H���4�ӌx��~�K��_q/�Q��ɺ��*�`�xϞ��/��b�o��i�PP��MI��Þ��q�g/�l���v2!��b�	a�GG�v�L�5�.*����Ó�5�G�d�Ȧ.�p���z�DUu�s<uR�� vÑ��ɍ-�'�vLq�?X���=����r���;�`?�d�qsR�e��/S2!�D|9:����ZU��QM=)��MI���b'��3K1?琟�?�Z�'�J;��F&�<���I2���nvY� ye�SD�9ڃ�2��~Pwۜm��*�Z��<�3������WQ_�����m!C�x%ٔK ����� j��:n�G�'����0�|��f�f�� ��W�L���:��/0�?��Oc�s&b��_k��:ʕ��_�E����GǟPO8.�3�qK܏*��X�!��[����y[�}����`7k�]�T��/3�>���k��%(�_�`�(h��7���R���`6���")l"y�|!��&�GYa;K=b�H�Ϣ��ELC��������;Ʃwh��&8�U��2b`u=���!�+������k�KI:^�)���O@=>�r��%�.�:��΅�+}��`�1�伮C��V��?�bl�t�4r��V� +��k|�o$I�".���5U��L`w�r-6�8���:���������8��|��A0��~p�j,˚�ۚ������~��n���W����R҉v��(��2�����nӤ/�z�q;�0��C�j�b�gB��^�Z��Y�Z(o��8�D�N���e�O���?w�t4�gZ3"��+���ۼ�ey[��.��#�}F�m��#`	η���ٖ.���^D��M��x��ǐ�?�+q��dD��x_��ʋW�uD!0F���P"��
�A
Ӭ��HSml EV�E�s�����c�� /xa�E?P �gTAn#Yz�S߽R@������k�L/�填sp0���\���d��'q�:+,��|�`�Z�^<��~3��XsVo���5/���p`�i�L��˱�ݘ���2�P��:��w�=Xp�]�ͪ��L�D��: $���w�UJ$�K�aP�/Cl���r.Y�.*O�Z^��}���Fc>�w�S�¨,�t�"~���m�����\����3���L�2X� �A����}���O�L@�b!�㶺��������ME��H�<𗭿�φ� x�Y��ǋ�F����M��J�:{��'UW,j�]�g�br����7rL(��TY����-�f%H\��/rA�k9�+��I���e� ��*N�1\%ZةG�{A2U���P��.ʵIԁ������n�y��l.a󛰑� ��}?6�2�Gc/]8�ε�8�9jz��my�ʾ��ɽ�X�1����[ť2G�����͞;@A �0A�d�^%��d�=����b�9{��ef����8z���S,g��F���<e������1�3?���@�p���ݹ>8��<z�o����X��\��I~c��z� +���[�?����(kJ�Aںi�8F��*`���!k3#$h�<n�����)'�JᒻH�Y�����M:(��!��ym�^�,	��X��ƑT�dĀ��u+���VF�'�'bn!�.tm���V˝5'P���0�`B�J=�R�i|���}�:W��	Y�eE��	&җ��J#�_�B��y^L]�1�f�B�]0t̎�`3\Y[��	5��G����~Z��d�T
M~8�Ο +���Y�lⱬa+���?%38G�;�m���	���r�ywA�e(��Y�ʲ��*�D�&ԡ��%/]?���4��m��NFk5gя�����p�/�&]�(�%�e9a�*�1"�`���mp�aᅓ��Q��L�;����	u(
�̹�w6$�XlX�7� ���w���T��,��S�8m�k�����Nm1�8��*�֧��C�'h���sG#�R���O4��vX�S�z�Z�)�Wg嘂��ϳ[�|�@�q��4��.�������t�-x��U�/��fJ@Trjm{&v�lM����:�3.<3�[��~����	�i �J©�q_�:%]��|��������A��\;�bj�?�eB���L���eh�$��.%��U2v�{��􉄶�e*�ˆܻ�no���y�WT�@�w�JЧ�F	����S( ��os��p=�
����f>g���6F��CT�2���(�*cY2�"�=dckp�ٜ��\��s��op��q���p�p����q�N�/p��YU/S�.S��~��7SuKiA�p��eh�q��t;fAyV���X��?�P�(��1尗N�	���l��,�o�������9^=g���\%���pU���C\�-�%c��jy;G�m����Zc��Q+\}P�G�eT�T�|͝2{#A�;z�Җ�L@1v������q�k9X=b�xQ=P�oϩ�2n����A�5N���;�]��dpP%�7]E!������ޡjj�ʲ3Ȕ7�L	�+�Z��H$���L4��)���7R32���	��B�b4@X���q��څW{X��7b�/��1|/B���*'l�*�q���>�bl��a�&���io�*��Y�yq:����3�����hR���.ޙ���`&v��͛ʏ����v�8�Cr��?� ��r$��DM��9��5�?�w9f.�~~ϱeT���U�D�p��ҷƯ�&T,�@{�'�w=� 
�橫ߚ��ԝd��2ɋ�?�o!�X밑�O�O�)1i�Xδ�9���uHR�)-&��?�,�!z^I�b�Xحrg�g�Ѳ���1(	f�߯i�ʽ�|�,2'���rv���V��1�
�?f�v�܌�1|T�)��������vr�p�t����(Иk�s���aH�N��F� ����;9>y��'���Ez���P����9&���������ߡ��G�jxm��+T��\S5�\���G<�����+�{�O}%�����M�/�u��ۨp���#�yڍ�5S%���uO�j�u�rI�STM��y�k�  ����{[f�h';���d��~8�Ճ���Y�ZM�(�W�^���vT��ۑ2I#��Rd� ��f�9"��zȄ�1�/GF62Z���*r����vb�����=͙�V�o��(��@��S�Kq�%F<4!4A[��D��v��������+ Ӛq�+	��c���1 yX�p�`���
"���!���N����zȖE��0gn��7���];�6��I���
~�|��A�&�6�G
m���[z�U}�E�vzZ����0r���^,�~凵�	�pJ��Q)�n~i�6�-��bQ0c�D<�I��th8u�UȐ�ߑ�����>{BR��`_���ƭ��8�cʟ�ă���z+��!���Yǩ	=�>_ҩ8t�!�z�З���P>��n��G^oEU?�}�ږ5�5\ �p$�8*������"��N`��`{,��b���>B�VZ���V�x�3�0v6���� UI�<7�I�H6D��T�#S�����߰\�Ł%
{A-MGkn�3�M�I�C)���C\�ڢ��41W~S��D��s�5D�?��\|���!xW�Bz�[�vjh�ac��(�'Xn���Dz���]xJ��<��5:Y�TK0�H}��Kҏ���ui�G���nW��������J7�oZ�*�8F�C�o����6W�����Һ��X�1-\ħU�]@JpʑxaM���⛻~�B*K��i�@�RDo�A��h���n��$i�oǽ'��[R������,�$�����I�Zy�͞�:�TE�hW: 4%��Ⱦ�p������Ƴ��^H�&���<0�
D�����}H#iT��8��o���@6'����6�g���g�Nh�����	m�X�v�۞o��`9�t�3�Jd��k´^�V�)Q؏x��@i7m�D߬��x��AɅ��-jW.΀����{�T���sp��3�mw�@։g� H�]�FI�w���)%��t>�����H�2tѢ�{�.j,�[͢j
R�$!�IY�=(q���ܕn��bKk���1]3��AM����j�]�)m�6�*Im��':2��(k�����kE籮.,u�dD������R ��N�RM�ЛZ�R��.vBٓ`&��[�>��Kp���4ƴ�2�^7��Z��><���je�(�A����#��nۺ�?m�
�.�����-��#K�7:bb��8h3�Kv�e	)@�E�9�v����Z_�� �_7O�9�Cv4�=s�J�u�vܦ��#ۦ��d.{_�4�,9�Gal�TZ6��VHjn���E!��UI$��>]�y��j�j)~��bjw��݅��{�|F�b�G�R�:�P.
�������7�T+6{g
d�V$��,F"3>�fP�$���~+)�/�D��=�C��i|��ԥn!8�0v^����\����7Ψ���Oz�bQ�]
o{?�k%�����5ysM� ���׎���Q���/dAN�:�' y\j���^Y��7�z��zE��$�y(�4yh~#[��c�-ޗz�*1��)�R%0��u�Ԗi�t�74Y��8D��a�T�b�_�8.r�	W�/n�@g���+�^-�"VePV��_����9�%��G��J����}�9Ėc@SB�S��y�I]�D��O�S�q�r�&����D�o�{�T��(�6~l2���)���B֩�)� ����h�+���X8
_=�%1�Ok_B�`�[tJ�D�� O���	�g��]}xZ_�!���D'�I��0�'��RI����W��$�-Cu�@_QS=�q"���K�]y�l��.B(�7�W�Fˢ�U1�H�@E� @(���@�맑t��2��\[�t�R��Y/�}���z?�@-/U-k14u~�n�;w�@�>���Ԭ��j��$ҌEd�%<��A{\:����=?��ײ���"Z��^�
4���W��uV���&�2���ͦ[�ұ3�{5��u�s��2+��J���gv�'t���	�M��>��(��#!�Ϝ0)�=��	�: |�q��6C��ؔ��D�k t��Ɓ�<Ug�p����u�� i0ЏS02c.�ꃶ�˯Ld�A� !��L��/HE0�F'ҔĊ�A�[��Mb�3�<ܯ˓�g�i_��J�;C[�/�d��4'�gt�!�$.�_cz�[R�xí��߹�!����*6*�\����6n�4c�p���<����l�4qUM���~ؽZ*w<u�7���1��!6�Z����Scd�gE�}�8�����q���u"�`�F��^���-_U%����Gi�u��^���Sd�O�j�/t�E^�����r �*d�;_��Sd�������_���9i%��?W��(�W��T�[�	�\q�mspV�