��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<ꊃ���6�@���P�8�ݲ�A�U})��A}�x��}э�_�𨚚���Es�sP���XL���>�$������.Vf��pj�׸G�W�&U�No�� �̻���2YOf��cmP�N\ס�(�������.Kb�#��;v-< l���H��đZ���(S���c<�٭�e�[��5	m	�A�}�>�M-7IR�Mz��O�۹� F9e�GC����#3�j�4�*����¾��	��q��px$��G���E~�:���8^ޝt���(��{A��̡z,}Y' xn��C�-���	�����V+�#���ȕ��zP[bb���v��a[��jU�5h�*z��Cu��P/�Ƞg@]�{�ƎҘQX�[`".�Mm�;��Z���ܦN�3@�����f�@f�_���˫���
eN��\fS���gm�j,�Z�j��������Q+F�g ���q$WJ�m�7��V�;�۪�n_�G��c p ~�n�(w�h2�2��c���lxL�}�HO�O(��ff�_���0��b=Xr�X�_��O"Kv�1d�ӧ����g�Bw�����ӇxW��&��ą
�=2i������g����̱�J�bF��av#ʅXT�_�����gO�;53���7*�|���nѩt�[W���l8�>�g�QZ��>Q{�S�U�n�.��a�D�6oȚm{I�v����8�(� ޗ|M��4ҕ�ݞ3V� |a�)ծ��Qzi�iq]L���{�ca�ǹ`	�E��РW_��6���
��b4�]��̭N�-��V+��(�q�3&̡�VYH p6�ȱ0D���%r�X�0'+�}��L��,�Cdvr2ј1�m�Ы�'A��zQ���x�D�`A[1���6�j"_����9���ś�������$��ָ[�L@g!��Ʀ|ฅ���0��@0�d&5�:z�d�	�,[x,�>�y�qqO�x&����:Oh�>������j��:S_uq�rx0_�I��C��r/N-o��t~�f[kx_���jA��hG����y�\�U�y���l"�&�nD�=��u������	�}G�I�&)�������GI��P��w��p�x)�����*��B��t�
 �jP�+κQ��2�z��H���0�T&��I5%�2o��H�g�o��3IY����~!*5�Ռ����;�;�'��~���jLyG�Mk�p�Y�����%�Hչ���O��sM4�\:�_�x&��^�Zjlr��T�,ĳ��~��b�{�"!�Oaǆ~u�b+iE��[���Hs�*2�&͠�%3f�}�L�[��xŘ�3^��DW[�a@&�~�9݅���I��~�((� �%/{�ίq]�L���������Z���FM�y+�=Ӎ���BWm�=4a�>�o0����M���z��4��
���u�"Z&
U� +�R�V�f�%H��V^
�ֵ"�?P�Z�����xW�W�A���ȏ|js�(���Kb�f�v��(sFWCb�hC5v�^(AJ�����5�|l������A�3���cqa��9%\Z��T�o�F���
>��F���D;e�h�^��7����.*� �޵���3�sb)���
�uZ��D�J;�Dӕ���P���-���(D���>eS	�&���C}�.�)�O,�1$@B����; ��l���Q�:���	Ws�3��Xc%̦���z'I�Q�6L��~��(p��̣޻&zl�1��RKW���*>=��.��_l�K�&KF�#����"���O���A�D"�H?�&�(~���)�˽�[@���ܳ�W8�_G�{p���]C�e��X�Ln�>�4䟓rͩ�^���5tkL
'���i3ɳ;�-n�����Fo�wa,���_�k����L��؋�O�:M�����\�T��S��]��r3fe�C�~���Υ�Ts���n�v�ҁ��ʾ�l��*�^tM�.0-�%!x�L��.�ƿV�z�v_�����t5Ut����� ۰��{�De�.��P3�B��c�b�P�(HB"���s#��0 ������Oa��z���*0��KcM��ڣ[�9�X]z�G���B�b
@����"v�EĪ��9X���� Q�wF[���1`��J3�������0k���uu
IMX���dds���4L�d^99]�i�
?�C�9FLPU�j&���0?��^��`[7�n!p���g�]�~C�����]�ZF�B�2������<,8<��l������"�4s�j��*$��9}(P|<�o4J�����R���E��gTU_)x%�<�����قQzwŔ���΢М��-X��k�(�	z�0��d�z�>O)|ៅ@�t Wf��qi �m���Ѥ��(q����w�I����A� t���͸z�A� g/�!D͟
[�7���֭���]����	������>S�����<� -��
3��Խɍ���^6�'�X�9;�x��jE��^��X��^vJ3�Òc��?#~��6Q]�kPӃ�'	u�U��-��g��{ڧ3Nc��Ԫ�kL�ؘ�n�>�R�mw�.6�/���=O��oK����-��c)�p��	GG�	v�Ie�o����+V�\�U�bY?�� p ��M���Jk/�4��T_4
`�h4�2�3��Mܠ{X���ia8D��\�)�_����{o���y���]�;�Di�GY6Ł�����k��E�����QT �^����UXD��fB׻f�T��^���Fh�O�X*���"cb����D�|D�yñ��-�R���x�~�I��,v5~J����G��6�n�^�NŜ��WyB�[�KoHZ�;��7\s���yNZ�'��I�����u�����ÿӌ��nj�\	S:<Fy���X��/e���"���Y_�F)m�|��s�&+�mDۄ�o�����ä�b{x�#�⡖T$����������U�\_?9��>��i��
2`n�K���zBN��g� FQ7̕��Q�6\*�jWWZT!���F��ݵ�;��ƨ�Q
�4��=܃Q�`eW��s�3���$#|�ET�8�m����nu/�xx�?�Sw���l��Fq��A9N��5�yL!�=�khe��(k9�46��3"�b�[Q�m
�TV�x��O���������_�TC
M�i��f��"}o�X˼4�3�,a�QU�~�!���9! �^|?��
�Y�%�rt�	FE�n�m�F�r��'L8��M-�F��Y1�IUUEG��a���./���fWv�r#؀�;
��A��5�נ��������u{1��ғ�k��tH���BI�G	��2�TU��D�k8#k��`�+�8��7]�*�L�<��0��>�i�j��J7��9���ff|d/7b��x�n��k�e)"a7�����" Q|3�V��
*7J� �۳����r0<W��F�<��Eu8K�v���1�I��r��5���_AyS��cu�x��.~�E�z*�yhZ�I�E��2�-\T�i��"}8R*E�Q��/����hS����q�C��̶{��=��_��K���qwI�2\�x� <���G>�{r�.���:�5?���WT����(tz�y�g�o�m����/��r=�]���L�᰺�ʚ����+d�˫V��=�DD�kO�[
Ok���A{�.�a�mN``UG4A�[U�`��-�n�&I.�����;G*�fS�+����p.�B%�}4�FM��QHu�Կ g�7N��Z\�{rC�W6��P�Vr��.�߳l`�U���r"�ۅ�W����Ĝ�[r 9T`����%ÖE�_�o��>%�����GNPmR!omi�b�8 ����q�_h�
�j�R��rB�J��w��f,�z�	w�v�qq�)��������q�>�Mϫ�����xU/�Ĝ��D=���
�t/��XG�	�=��;�7���՝4�����/9X�O<3�훬��έً�����T	�cѽ��� �����|Yf��J�������:���
���_��\���/��'Zx�)G�_�FT�\�����Bj\$wl��%��^"Dt���xgW���4N�=�*�{R�ɳ1s}��=��6�2�D,T������m�㮾�;�I��0��z^�)��ץCf=6o�$�����i/3���Z	԰����c�-����;is�dYt���O�/��2cd��:���v��%���^��3h��B;I~��YK�jd��
�4|B-�S&�f�KS����U�:'<�� c`r��WLH2�Y#�H��	��)H� h�$G�RZ�>�i(���lgRr��kN��U�����@�	%(ށ��K��x�6*�Թ��44O`Yh����I�v�{K��"0�)yPWrB��f� ���Z�YF\�8��]��Zby����5�q,d ��|"�u���/� �S�S+5�u���"gE���7ب�<}^�ŵ��ڈ��5�뚎���?�\՞\�G��6li��򹸀��u<�W����G��ެk�9�&1~=�^�U\ZB��W��`��������<�����v��q�q̝��Y����,r�{�7��Hn��j��L��.�_j� ��m��aC�Hm|�8�RF�QG�&[��a�W�s���+��3|q/�f"x��K%��"o��ֆg䷳������櫙�܋���g�&���Z��q��EU��"���s�E�������6G�lX���l�����N�[m��E�4"�;�´Bލ�Nh�Yl$�im1�W��$$�.Ｈ�ڈP�7FT�Jn�z#��p��ζ	t�<౜9G��
p�Br [U�\Q�`?�>2)�!����#e:�2��1y`g9���^��;#��f0���^/�����U���lR�Y7�ђGn��R��ZS���5a�c隀�<V�
ˤ�FF;�%�����b��j}	��ޜ��BvY�4�w�@���㶙�̈́��̓�7pc�1�h|_`�ŀ��Xl�^ub�pq~�~�u���zZ:t����bb)�}q㤭��)�)�a�p+��{��)	��j�O�c$ձs[n:|����T��O�����ʷ���ۣsEL�!��$j��c-��Ҟ�m�ZS:z��ydG�ʶ����o�*:�b��v~�F�δ����14��N�?�g��;M0���ǿGDe��c���.r\h��3�I^.Q'�~a	W�
���/���^�}T�K�V�0='��A��̉:5�}�L`�iC��̑e�k�����Ѝ
H\��D�4�w�k�x�����At�Y���"��Ĝ�9S��^���kT�ػ�(T%�¶�<"}J��dsw̥�Ÿ���P;As�ҸS��R�B�D��IZ yVNcZ(���
�2��	/<��l%{\��y҈�Z%R�o�����9t,K�%$zn�#m��T��k_�l������P�k��T�j�.�w�6!>U�����R�� Јb�x���\��h��[���azxi%5��eKWE��@}��$"��rO��Y��+{*�����oR:L���"��j�z\Ƿ0#E�x��ߝ��� Z�:;Ё{��!�}�V8Ub�:�{} �3�I��ũ��b��r�ìv���]���Y�?Ԟ��x�ΩO�"��=tǰ*�,)P�)B���O��v=����$�?�\ Y�Tˋ4+6�4�+��8�7%x��P��e�gC��>6S(��DA�%5Z]X�TFV�j?m���D&Hzq�mk��i]��RM4���m��?�8�����nv$W������ws�eN�c�`��Y������#D��!�XL�yx��u���7f2ӝk=���n�TǳF�T��sb	 �	��T�S ��%�!��].��n�w1+!�f`��YMFVt�(i=���_�G�(Q��v2������<A�^o����L(@'�t����,�g]�؀��QT(&�L�鴋8-�BX��Eb��e�R��]�G�!�Nc+�h�v����Y8<�Fa%sW5c�����l�d�(�Nx��	�Q���S��&�����O�gIn!�l>���c�"��6��h�C:��9�3�NI����`��ܯ�!���,K��[���(�_����g�����92f�J�>׏JcH�����$�<PL�dY�</4>0���k��� �ۗ� � ���Ծ	�r}���❐�.mK
"�/_��������u��|���)Tk�;������O.�f�ŧȵ!exT �ٴ��c�ճ��ǽ��$>�e��}Q*K��������;��ӏ�Ώ�����q�!�d}g_3�MF��((�§�����YY/C�i�q�C���Z2�*���F�]H���3AwKۓE����2ܢI9x9��o���6����#��{���@?-/���hA��c�[�kXQ�);������3��O�y�!�z�u���=�:�\S��smU?Cinp\�5�g�
:��Y��CkB���h�eݞ֒޸�g��b��;rX{{%�b1�����bD��@f0�J���i�L�_����M��<�h�v+��+�bN���paS��(VБJ�6���q���e�N��1��mf�nI�
�W�V+Q܇������F�Ӳu��6΂�*M@2�����e�?��	'�0����;�u� ���V�mraktM�3���/�r����s%�ZH�����_��X��.�Q0^K��X� s�}�N 1��aԀ�P���;�QB7�7}�֑�%0�����ZT��Є���Ѭ�V��P��2�9�ĵJ<M���`�7
��@:��B>.���	�� )�Wn �;M ��۹F���Lޣ@�*=��JmI��H9�s���9�6���"`f�Q���A���nl6-�)} �l��2]�D��Ww��)�n�3N�D�^1Se�9!\�/��zz*��״����	.��X㘰G$��"��y7^���%� 
f�A�s�z?��B˽|����շ%Q����W�H���MC�!���[��x&k}�/��g�z�g�I��q�a�~Iƅ�Q����X#�*�<��1�����^�^��DD�)��'v{�Q�ӓ������.��2ɡy��-�U� �`�����>�R�Ae4=�)OΓ辔34A��|t��U�,D�ka�M3'���^�Q���T ��������8��f�6-��B�'�ΛT�7Cp�+�"��ga��l�-2@Da�<A�0Qz3�h	� ��#�i
5x�q�[ծ,L���G��u#����VZbh�cHR�\��^�OkUԣZ&ۡ���Ux�t�^v^�x��+�bt�.~y��I�m$�ӕF;9^l�$�ZY0 g>R�'#�����v�w{ҥ�E�v�G�IU�i��WK]P�&M�?���|��u�ݞv �k�%D�dA�����:տL��Mn)���F	�Y�V;j"��D�z���D�;믿�q����=
r5G�XE��;{��Lн9Gvm��G��P��r/;����AN�����V;�h��Sf5��+��`J��qb���L��D7��ޗ� �E�B�HO�)Q�n+�x��h9nE5Kk6�5�Z�ђi��A�T�8Z�e���Z��z2kߐ�5�e2QE�Z_+��j�Z�(+c�߈��qS!���lo�'���E�'ލ��DԼ��c�
}�Z�:����^]�ZʯIls9q���-����|��}�fd����Q�zp+Ǖ/i��heIe1�I�-�}��'�``�}\��!��ȩ���/d�ŞC�֡dP�~'���]ٶt�����rS��C�t�\*��C��F�ˮD7�?�%2d�O��u^��7'�bE����V��[c��U����!|�%�(כ5tN�����H��W3�cS�&�J��Wg~�zY_����� G
E����bu���H-!AwܫV�ژƟl�U��ﾷcDhT"��	k�`A�^�b�y���Ă`�!kO�cEjr[Iq ��Wvж��c��_%�s(m�s�X�-����j���8�'.����������A��L��i�'��+�*r���3�,NF�;��f�)��L��&��m�C�n�����fjp�5h�ޗD/�'��ʥ�N8Ay���������)@����:^ojVK��uѐ��*p�!<$~���ѭUZƮ�'lTWi�h���		�d!��2��9T{������?�w>�9��z_J@?�3#�����>D2ݶN��;��r�u�q%_����ʬ�)M����:��*Q����P�5������O(:�/�bo+�����?�q��U��b.G�4�$�&�G�F� �ր>p� ȑx��M�|Fğx�w��o(��%$���7�h璶7]�����H>B���:Z\ݥe7$��<�*�i���'���&�F-�J��RR�o�0�eK]��? ���Ф�P���C�o�g���k�5�gl:HF$<��\CO[p<3��=��� �]��`��Ⱦ~��Z�Z�h}'�%R����K��	,*���ّ�>U 6�Z��i$5�9�|�(+���g!	����?���Ӣ,{%vo�/u����2*���B�N�%���^�}�\�>����� ���Ih�I�O��̈́_I�c�_�vj��Ų��:��V��<;˰���l*�~�旆4�Y�����ʥ3�lt��]>n��T����'�S�1ἳ��<*vF��%1��D��Qc��{/E❅���B��ꒃ����6!g.��AX�U���	z�:tsq8�o�H1�Q�����yg���A�_�\k����- eU�;\]����Y�`�*#:/\��n����{���t�f0%�}��a)���Ufc���P�A��41���g���0�����~��B�����`0�_��*�U ��/7���s��$l�8;v����}�QL�ѐ��ooaNz=�6�6��N�&@���N��eɪ	