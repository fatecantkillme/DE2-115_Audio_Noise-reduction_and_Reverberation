��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�uwC�5�b ��ϴ�	+�
Ct� "�J~���z����<
�����'k�z��ߵ,d�.��Z�Ӝ��2�x$ҟdL��h��ʔf��#
����;�;m�ȋ��[F��E� &'{=u�3jg�b�)��LA�u/5{<	����oiܒC���&�'aV7������~^��ލI�e͍��;W���������R��DI7t��9��1�(�XS��+3�l�ɤ��{T[���L�l�vH��7�*���}I;nF���T��7v���4�9X��Dﾚf���z(��)�ln3�4�kJ�ú�{�\Ed�m@�;Q1�{gT=h���T��E��~%�T���.���vSF\@$�k\#p�l<�sㅅ��_5�C��G>w)u���
�>�݂�Å�}�9۟�>�U<�[F�~[�b+�[)��c(O؟���%66���2VN)g��++C ��@��'-^���z���=ّ�Oz���率���$�I������:2�h�B�s��Q���Y�-����=�BXd�eϤXtSsa�qa9�(������j������������A���)8�4�ͣ�|���%��!yuU~U�{�:�?���4�2:��[��+a���	�u5|k5��~�"��sU ۈJ��	����]��0\��C��6,������4k���D���3.weUX��Z%�e�J�uKf���j�w8EI�Ns�k�����j���ˑ{(*��� �|��gb6ǰ|�Z!�%q�%�o�׷���rzd�y�DV	Z�E��	(Jh3q��F���&��?p��L9	�q�C� ��K�39�>U.��벍�䱥[�(FC���ɓC^�%�g
�C��4�˻N_ӂ�W����T��t�}ex~�Ql_�9n��G�o�Ǭ�V�H��~�4Y/GW�|�ڄ��N]�A���}�Y�Ӕ3[�g�#g���At��&�����P#,/D��J]�r�^���CQˎC���7��U��!�8���nR׼Mg�44U&�q��;�tn��[�d:P�~-��
�����;y)ti��H�"��`�4��|l�~�.��#a�UC7U�Z��@x���1��~���J2�Q;*�����Cw�mZ5�����T�7�/T��J�5�����[�����B:f��輻`���u��9��T����C���Ө�;a��8��j*�}Y5�rj���ܹ�F2`��l����m�=S�2��\�����@��W���1A|�V����7^я�U��H�]��c���G;���*�:Xj_<G2ܒ���D-؉f�>�~|nD4�rQ�hsC�y?6�n������$������dx,�9�B�m��J����j�V9����0�J%���U�CƐ ^(	
a�peT@9�����?�
�������	���i�� -t>��ZZ8xG�"����/9� ?���auZ4�*Zƌb^xo�n/�g�p�k5�!�R�n�w4�����YC!������x��J�#��P�<VXJ�:� ����پ��x]���@62�qIr�|*g}�ٜ�<��S�v���������[ы=U�
ngGŎ�TV�q5l昵�����W	���č#�jUa�-������z�e��kl�^$)���4`m?�Z���<���v�Kbޡ��-[B%�>�k��	�s�;���LF�j!�󯟧L��}qR�n�$6��P ��������!»׋�.��'��)�yg��=�� ����m ���)����4�~���6
BZ�5�!�C�8xy�ᖣ�0'Cs�m4M?�$�F���7����u���-�����S~B;=\@���V��BPi��7��b_F>�o;e����r�)��Z��h+��ᶄE�����k7ZRy��OtfCg��LӁJ��_����y"
T�Z����w�tt�v](�p�EI�:Kg�i�;=v�<t�vX���9M�������B��ï�q`��d�euk���>����g�>��A-�Y`þ$�;G�AQ�����K��B�PJ�ɡkDݔ�5zZ��SRb'Z���_lԱj+2�3�$����Y�S��2�[��pp|��*�Z���G2�lO;De1���c7�%�9�SOڕG-����XXi�
D��3� ������c4A�9��}4��?O]��@�sUF ��lͺJ4U�H};����� ��w8���RP)F=�+&�,kG���Q5m6-�kY�{mE�g�O���wL� ����j�E��U' �����B$���w٨��U-1��}{w�ul���7Urh�8�v�m����h?ꔹFG��f�<T{�4h�<�
2dO.֪R��:ׯ:���zs�<G*��VP�Q���C���n
LR���ύO=DfJ��Ye(����B��P�7��`���s������b��>+6��2�͗���幬����K�����1`�T-���]|^��Dj�ӻ�D��9ݓ��M_+�����{&E��.h
�r���ꓭ��;=�����x��1�mx zC�!5��/e^,�%�����u������Ƥq�7|j\u�#��s-簙d͜� �7���BYݮ�[��[ˣ[uUH��ϧ�~�}0�Ƥ����:�k�H&��$�#�8�t�4�����p��^����o�<�ŀhM����F%WC�c0�4�BHFW�+� �ʒ�����ː���*�0�������t��x�>N+@�I���P���\��(C
4�h4�
]K�Qg���8��cU��4�?��4@��ݦY�~a}�1�c������M�����5��_֋�Q��74�@�dfhS��F����@A�t8f���YOZ|%RR9��t_�=s���j��	!-A��h�
6!��Gf~���l�A�}\J���D �a�!��]�ù��2$�Y)I�h(�&�������%���|�+��o8���u��P�`����%���`>��RG�^�D�ZpK�N�_�!W���y�����>�(��θ&V��7>�ntJ�Vx�ϥ]"���I��%Vj��}�n�u��lg�7�,-�`�fL�s?�P�\$�#'Gm���N7R`�ZZ�d, ���#î���|��h���h�j���VX������d��)ʤ����d�eO	� ��c�fJ�* �^9�g��)n��rx�ړ^��:9�g���F	���`��M�q�M�-Z�3�$H� ����ȶ9yk\�\�&el�@O�;�<� �NWa����^:��2�R��ǎ�g���Q�8��Iqy��]ߧ��ܚ��=�i�Q�d����I!�lqI$J$uUO��I`=��ϴ2��V�z�W�N��*�ހ:ͻ��5� �3�&�?T���6��QS�#Q>�����Y)�u�o�X�O����A��V# ��(����*�@{��Q���SmP+�0�Mt�:Q5�/���TV�y�)������i<��/���eA�a�߽sN(8H���/��F�i�u&e���(�����5i��&�ȳ�c�殦���emg8��Ń�A18�2��um=̚�#�Y3��W�����e��mƼq��{��V�H�8=�ND���n[1��尢Rm�%�5锋���ī�R�oݩЛc�P�� �<���*��j�@�O�6&��+�qF�2w�7;�`،D凌a^N�A���~Н���n�,1����XX���4JV
�&�Kb�:hO�ŮM\ٚ���UL���8��kͺ�3���< S�ʜ�to��f����r�'�������'7j�#&�*���d��^�k�b����y٦kn�*<���mzLVo���Y���_r�w~ś�{�=
R�ܤ�~�vB�5�~`�f^�zL%r���pv��,���d�v���7�k���y�=��}�������Q!Ad���m>e&�1���<u�$ܵ�����lݛT���03�ʄ�}Ԁ�O�T^V[�{*�o�mؘ��g ��n�}�UM�&���o��$x�]�b'�3�	���lv�q��L@��g#j��!o���s�?����(��O0�,�R��P;�Mځ�KT�DtοC�L"2��u��	��q��5�4�#b��TS�\�ќ�훃n���	"������f7��Ҵj���=��״�m��e�C�'Fu�H����Mc�����U
p��<Ť���w0`l�P��kVo�?w?�a��۷O/,�d�\%:�و��ՏjL�l�Bc�J:N�Z{8��l ����yփGԕ�7[���5^~Lz5�*�iƿ��tа�E{����a�4q��j�p���R�8���$ҠO�#��U�{�������U!4���!����,����,���zD�|̷<�d
A���h�&lS$  P�9\ S _I+�8���	���'P����u�������#�uw�j���2٣���A`!biJ��g����\l����dPU�BU�f1w��U�����Obg9l&��B*��%���$�`Y�n�ߥl<Gf�Co	��GtZ-�'ލ�~��ZMˮ���oz<CB*������*����Bem�����$L�ۤ��TY�}f��~��qs��W�&�z3 ,��9��u�MGN�`�=���5ϵM�M�9��T^BG����J0�Z-�;��Y�V��i����X�mB�V�Gk�����+����ĩ���(խL�ă!���)�)��d�wח�8 h�ƅ��r4��y*����K�w8qKx?)�L�]l�'�QM}0���%ő�����2��_*�1�,�s�6��y��*u�LP��=O]� ���)�E�@4E��U��� 1+�gu��v
U���������x�5J�]�*��HcA�$P������rz"�s<ۤ/H�lȺǔ�qu�Vw�u�&���<]MEh�,5k	��n�����ɇI�M�mH;)F����dV�k0��ߒ��ָ�!��w�����	�{��8��KG��ح��y�Z��q��@�#ݭ04x���^B��y�[4%���
 {���O-�`��G�
�����D�����8� �tŞ����Z���p���Z}���uL�v��v�5��=v�?�U�j�c④�$6�Vǝ�nG���ҥ���"z��L�=��j]�+
,=�R/7�	�����l���V]�S��z��i��^���,C��و"����C�xng�{|b��w"_�Iv7���N��#n�/�0`(�liX�.܊=M#�[9�Xm��;rC�uB�J���
}������T��W��2��\?z�Qq(����^�9dt���dk�E��$���#���)NS�ɓ>�k�}�Q���TfGv���RX��$m"M���ʈ\dA_�Ymgf,��|W���*��A���.;�vk��3����f�șF��Q+�3V#3�&vX,��I/fkт<q�}^��D:]5����D%�-O�F�;��4�)Q�V�h�p��V�d��킌�MͶ�:B�G�b��,��Rs?%�!<��:�3h��٤Xi��5d�%Gس 9�յ���؇���AEP���\�>F"�J��E�(�e@�ssX)xA/f����3���I̟u�����D�B�<�2�I1�,�M�U�+��ܢ;^��ʲ�}p'Ħ(�S�=_DG�I��Z��Uv�z��JN��+��N���������_:÷�S��q&s���}�1m�QH�b7�:�-Y��w��Y�xb��v�S�߁ ���&��E��u�ܼV'$��������������$0�s߿�w���Ȍ���_�?�|����O��[Obn �'�U|}�q.гW���|*Q{;�N�T�'#��MY�j��]t@��
�T0�����@>��7"�vG4:��'�_v���'g'����^��Qd�(���}�z�m%A�D���R�B���'zGf�k��C���%jѶ�wGf��Rf���"��o7o���ڴqk����b�!/l�K�\�'��d��hae�M�����V�j�\�ke�b����=I�E�
�JŶ�5�QE���Z��;M5������o>����ѭib֍Gw�����FE-����@��+������_�N/����u��q��@���~�}>��������قS�x~'�j����cz��[�!�/��˘'(��J��
��i*9e~q� �vf4�L��F(h�;�I�I�X^�闌�v��?�7�b��CΚ�/stX�,C1G��2�m�*���O�,����<�����;�c?r,������4M��L&ug  jT�Ԃe�0Ja���.d�\��Q��1��z)7�.)Z��b|��/ܰ���d�G��:UCv��	K_� �r)z�W岇��ӣ�6$���m��h4Bc�uz�|I�!t�nw#���o�9#iUs����*M���,���oFuIq�l��m�+�Tq��c�T��P]x�&b�a4g����������Uf���I.��÷�����A�H ��_h|��D�~�T>��w��Kj�j_�M;�y6���H䥟���~.�+��e	ĸ�'|�z6��`����t	y�AL�N�e��way��0q3�:(^-�vO'�y���*��b�;��
`�`h/�*��,8n�̷�;8��,�ӈ8�s�:$��?]�R;�	��?H��M��P�⁂��y�����9��~a��"���\��bBY���^<�cJ��ѐz�;ev���Pc>�"�-	fi4���!��� 2^ X���]H��w�E��*4A� 7z���q鳶��=�r�h�<ll�q~�Z�|���gdF\�I;�rƤ�8߁G�h��o�4GЙ�6ֆi�8�W@����y�����x�$P���ޕs��^���K����%i���W��vߋ$���G�w��%4\�8�t�~$x�� )�ٲ��)5��Pw��`��̕Mw|��/,:��ΦK���W����[@[ruX�zy����i����Sf�=�N:s�w=:�
�J��ݡ��tG0�g��
��v�3N�P�.����n�"����p����U��+�aMn5\��|P�i	�����|2���v�H���sc��6�q��<muA�*9��/.��A_Iz��#��V=�T�($f=�M����Mh����jhC��I����	0�xщ�_&��JXF$�*q�	ì�?�wl&������:���PN4�/�`�si�o�U/10�� J���Q]���d�mM�]]~ܦ���q��)�~�T�76�fF���_
��ќ�0��$VD��~�/w�huBo�����S\��_��N�yLI`!4=B��C�#]e���"�ɟ���o+���,�%>�㏅���V�HGI��(�b�uG�;s�Q�������N1w6�x�@P�@��h��a1�T��/������ٯ�� ���v���� 	��,�/v$���
lG��G���G�u�[s1�cG���#����(�M�@]/�d�Q{
Y?&�B�hS��O��?[�Q˛2�8yv�g�Z�E��B���{��
Ӄ��z�� sî���"��DȽki4�+�v%g��z�ҳY%+/�i���e�rb��EP8�N�����n��o�颮��>��y-7��� ��bJ�_;��/ w��5�W)��g9ɽ��#E\�.AL�_9lS�E�dQ=�K�HT��P��'�Kn]S��L��ƣWe�u� ���9�6�rt >��������J�'���m�l�H�[rч۫0�$� -�`����04bH疂DA�H����ήn�ݳ�掹�IM���.BfZ.��f,HӞ�>xi*��é�S��a���7&w %A�o����M�$�(W���Y'-&EG��챚�X���0%%a�W���W�;G��Ȥr: �w���������i�9�&��9�"l�w1���G��_���莖`h���}E5w ��_�e������o�Vd2H���l��fr'��P�������A͡��LH�9�I����4ɉ�%�|Ύv]���յ�}���^� u�a����T��������,�o��/B�x��Z�tkb{Ա 3�aVՠU�Ȫ��J$�\I����@yC`rEAE��8���d��4���@�qg�� ĞzE�On�׭�ׅ�C2�\M5����Sa��'S�p�=�����1?<��D�w.��\�Z]��п�E��*Ա,�5����g�w}-B�� ����q2����5�Tlo�9��aB
�z��v���&	g<��|��a�L2���jԨ�8oz��7��*�e���.��s;\�&�[�3��%X#���o ���4�<�d>R��`>�s+)����d,_6M��S��IB�P�0�Y뽀�)1�AE�|�a{�P��W�P��_x�>l!�hl�_�[8�@�0��ʡ"���>ao�G1��7��	]-�d=w�Bv�h<�b&h[y��a��Ap8�|مjR:��\�x��
-y;�a��"�����A>m룅��`'Y~��d�Qsi��T�P�߮�<��JC��ciL[����_����_զ�;�ŝ!�)��Ӊ�2]u�	���z��*�$Sxb�G��o�Y���[%���{#�A���t^���Zb�"miꨇt[Zc���#�E!�����FT�ױ((H���Pt@T��h@����N)��&˥�Dn�{w����\%F���׺�Y�I��}�C��_|�%��w�A�R<t��]����K��@ʃճ��䨖���Ŋ�����G��%��/#�>)�.�h�9��(�@G�@����`wP��cs��q.yK��ݯC�S$���͢Ab��,ՊI���zi�r����#E��\ES�#���b}�y�F��9�Sal�v�-���C����_�#��id@]%n�^& ��Sk+֝�=��.�,~&����4�� ׿���x�Aq�C�ŉ0Q�=��
 5,�a��"w�il`�r�Z��^��n�%k�o)��z|+E ���ԯ�T�<a����IY3 ���X?
�������M�de>o}��[ji&Y75�RK2Z5����25���Y��t5B�LK�c�a�Z�K]�R�^`���	kpug;���w����=ݡpeuħ�ذ����V~�z���ǳ
�v^D��;F�:�B�*"$�L�|��6��E|�bw���2ju4�Lʨ�5;LS ��cA�f^�A��\���B�T5�m���x��
|j�ypP�.x�4!~AGR�V��YM%/����QxG)���>��݈{@2:�up��T(Ē1�n�4�)Y��}Ua=�K�eb'�!٣�r�j���L����̽gW���h����Fjñ�w +ޠ��؆��g��GU_�_��#��&Z�#��^%	y� ^p����f>�q�T(�ѣ:5�B$�0�Ë^H��w�{�Lu��WVE2�ul>��_�m
�ǫ�kh!���)٠��P�����Q�߄�=yL�z��ͦ^!�`ek;��!I:Dv ��>��Ь>_$��P�_��n7_����{�;���ǵ}��#�]���e]��%���v4OQ�j�;�C�%c@ߏ�@I���#y��tf��vޖe�m��B�Kຢ f�z"�I*�N^t@�%��aڷ_X�ac�! ����f�����ӧx�� �4��[қb�i����� e����qH�vѠ��F�5y�`�����$Lh=�S�`gFc�R��E}Z<���̸����C[4����T�R���h�'G�v	5������oR�"ȧՈ� ��Oy�N��=*_��aW-�L��.T��p1���		y�e���eqE�T*Y��O��ז����0f2�����(�fQp�P",�AB7�2}Q��U�+��"��M*jp\2A�ů�bG4���A���l Ey"r���$m���Y!�Hp�O�B) $?���Nm�5�J��FZ_��g�C7�������r�N#��[TK@���\֜�I��\��a��-���I����̸}d��#�-K��a�V�P��&D^1`���6M�:FV���Z����g�M��S����[b��%�U����U(��>3.N��
a!JX��]��n�P-����(����#Kj���"ܹ<�����b������L��}����ˌQ��(�m��C�`��Q�/Zr��>�I�Q��c̀����W&����7���~��^_����Xʴ1��;(�Jq���U2��p�|��qK���V[gڤp�5��%��{=��ㆤP<��+�u�EEj��yQ�#��Z���~/��UM�ꃊ8i���p�`Re�k�mT�k��g�@.D�?_��_�y��3�g����U(K���~�1��g���i�ph��jIl��>�w��|<)�93]��c�s��1�,eڼzňFY�qr.�l؟Tܻ�W�5�����
ԏO�U���㓵Sb��7�To�W�8���e�����M���7m��+�'#w�U��'�ZoIP!%���ύ�#>tN�+V#��xyr���R��=��1���~�E�"���͊��Ig��	��½󩻝��y�4 H�{�����n�=�� 	�^8��I{)UR8�TB&_�a`�4�����E. �>�{�:�T��U����9���7�{�>���w��2�=��i~�2d���"���@��}�!+ɀ��D�/n ^$4U���O��|?�:v	�-��V��h���v?=|A\	[����@�!���X�D@T���R�j��������8b���້:�	�ڄ�
`&_F��=f��S�_�N�6ߝs����c��,Sx���<	�բ��o���q�߳�bܧ���LZ
b���7�!����f8�:^���P�� l��G������ �s��8Ǉ��-��V�֏N�L�-��3�b2�a+��U���&i��3���Pg%M��H�� ����a��j��J}�sl�UUB�1�<1Ζ���fg��xD��c'6S�F�I����K�	�A�}��j�����u��:~%��,nt�8��9;�[�w��tH�?ƅ�J��X_��DF��%��>���*&�f�I��i`:��(=@��9�E)�1»�:¯vj�.��N�p��m�ʻ*�XԀ�e
#�
�D3���l]Z�$�5�bj'�!��+2��[�L�)��[Mk�s�GO��DHAyw��B��NO�6�ܒ=N�4������)��0ʫ�j�,I5�PW��F�3hǰ�~���g^���Ҳ���΅ ��5��8�1+�.K2�`����sH���Mr�EK���HM���׹��G�Q���~}��e�\]�:���!�3�� ��k�\+�8a�[<��ŀ���癊�_��qbIw�l��;�{��ڦ&L��c���z�f�i��a1��y�`�+o�����������5�B�{���&�h*ђ�>oI��	Q���=���5�8M��X ��`,�|r���!��*&�yB2�4=;���@�\h��ҕ*y�i��b�R��v�h������L�����({!���r��
���;4i�Ӝ%6Â+c�g@�
f$�	�]
Q�_� iҥ}C��3��s WY(�lx�u7��МK�u��d����Nr�hk7^�2���f������vS��"ufƊz5��б��-�(�7jS��G���d�d�fPQ�Mq���� X����u�{L������o��Wy�mߞ��4���W�l���^僣�J�ui�Rg'҆��׷�w1t�E��L��~<�6�8�9#sNX�/�%�:J!��_V%D�L'��Y�_�Iհ4��!`1�U_6���po�$h��4�(���p0N�Sl=}���:�S�Y�ŵ�K<)Q�S�~�4-&y��8t4���T��2��r�/���Л���Vװ��3K����l���U��[��'����?�����~��R_����h�n���eM�I��R!������	��f�"��-��x3-��ٖV����x�A\�eK��\���� 4*��D�,�E�}QX4��֠���� ���6���zǮ���;1���;L`�6�ٝ`[v�7�o&�d�=M���8k:�3S���[D�Ζ!w��lL�8�78[3�Q`�~FGKЯSb�Qj~k�	#P���l�mn�5}`)��{[O��}���>5x~�ڶ�6s^�I�4W��ј/�ɩ������IP�Qy��%�Cf �U�~�!��MUUMx.��` '2�M�<^��IB�F`�3�z׸3�}���^��珏��`�'��=XAq�J�� ���0?8T�. �js�W <�!�1�f�\�HF~���4!K��^4����r&���Ih]�mkQE��f�t���0��n�sw��(���^��_���C:a�.���������٣�|��_$衾�l9|��EY�9m:�o�n�	��A'��3g��RmX[�O�2ޑQ�*a��&��l�5ɑ��m�׍�����ﱣ\~oO���0�ֺH�Y��-�$mr�Q~X�3������r�L�݋��.�hDq{�»�h	�U1=6sKp߈6X���m�Ϯ����j2]x���-��k;HcE9P�@���by,�f����@�,�a������]�=�땁�yوC!������i��%Zէ@�P���0B��#E]fbƱh�tv�7�&=o���0D�e�c��d�Nu6�ExMh�lT9H��Kۼ4��q�1�V�
�8��֭�>	�'߾���v͵�Y�{�_�d��5��E��f� �������tH_ai2G�>(�K\O��g��aZ�/s𽘲57�$��Ú�*��G��{b]NXy�EϬ^�m:�J,�'���>lL���2�Nх�cQ0[�vM�����(nڸ���YY([d��~�4$�s�L(��L1-��T�ָ�%pZĬZ���̙� ����0�q�'�h�Ā�yｆ��n��C��Q}�d672 �i+&�;u���]?���&��6�S?
��H r�$f
�̾{��~p���p�hSq�<&L,�
jP�C��l�k��4M�M�</�F��A���^����c���7n���=�o�}�$��a�����.!_0��G� ���d���O S�I��iD��Qef�q�2��9�U@�Y.��"Bd���U�t�Կ�4V��(��E�P��������9�#�E���C��P+�Ξf2�جQ��Lc��"��X ���/:H���[���}���#�����@0�N�9���?���3Vh�`�ƘB}j�N����W`�����:�FpM\��0-1?h���G[j��b4�@��;v���T�����Mt�t7�P�0 ��6'X).�3C���n�tHr޲h��F�Di� ��̯3$o��~8hgzv�!:T@� ���Ƿ;"ր^&�����p��<X�����81Hg�[��ONa�=Ѐ�N�*�zr���i�#��X1'ˠHG���99��>������Ws���kڐ�.�@w��'Y���}:�VI�E�����C�M�S�2Z�l��p� ����	�`�y�k��|���(S�v�U�b�����q�2H�����p\�[�s���bO�;�
M�+ h;��p:}Û�����B/�����AI�G��b����Hr��?[���&h�%
uT��h��TA��Ϩ���� �P�"�l�V��G���Ń%�FR�3,",N���׬�������{��]!��T��>�w!/ּ�M/��2�g���ؙ�7��z��*KM!%����ȓ�x>v$���}�>�*��V�1��$�$y��M$o��7f~�J&=hf�=��%w;Ȩ��2S�=��]���V�)�D�SIuc�XC{"�bNU�9��C?9if[d�H���K�R��Ɗ��Y� w/Ꝟ	�.Q�j�s��_q￳�����ׯ�J�a�u��/_G��#�<f��پ���??�qlC*�h_���;�^�������n�� �v�9���n��۸��Q�Q :�V�em���^�ν[\'>l�u��_n�K|�ϑB��joi9y��b���h>3��8�[Ò�<�(����V�4,i������w����G��t䉶�����H�JB���g�~���c'��6�Q��k�|ʹ�ii�D*�p����bb|J�����Wv�)'x\[�_��&at	|�ǒ9��s�����W�[�S�]��{����(���L��t�2M�����-�*(N�]M�A���I���B�T�Z�D�V:�3y��6�I����AĒ��P���%Y��\G�R��p/]/M|��.wHF�ui��-*�X�y�ĽQx��:B���&�)�&���a߷��M�'�"�x�!n�H�Ē��>�iO�QSq��{�6 eZ�G_�@�G����k@Bn����v���V�&I�Q-����-���ջ�6b�⪉ʹ�|��J0���/�Ґ�Ҍ�VPr֒����o�A�q��)]�1��b���w� 9�BE1a�_�����AfA�~�B�Z^Ǆƞ������0 {H9�jan@�<ah�#����5��C:q��Q��j�\�1�~��B�3x�B�Hte���6$����X�X��"_fM�<},��n�6���*���"�*{�� ��-������?�$���D����3�wyA6=����{m��� H���,ck�HU$�EƏ������%���#lf��&	�~�^6j����#����H*�	����q��N�N㪤h|Ӽ�]D�����0�����ƺfehN��4K?�>��'�]YR�Ďq_	K��<~�e�8�iR�rm!�)���� *��m 0��<d����>��;S�Ce�U�+6�z����m+�P�n5ke����[�G����d�:���A�:{��e��#�Ӊ.$+���;J���Kݼry{�D[S�j���U|8���B;B�s\c�x1�j|Q�#�G4�R�j<-�C.=�;�a.P Uǁ�Z��T�:��z]�k�p�)"�����A�A��a�#%k�r�ĺ��:>�-IH({¤����s����#��:� >f�f�mr	ɦ"�>��xߴZ�w�}i�I�K
�O�)�2�a�56��L:��Ip�b���xg�f)���#T-N�X�ص�� �D�|���b�%Q�:�Ǡ�OC,a��MxZ,��癶����o���܊;k���[�������q��>]����[�:��~ƅr�Be�tu.���0���W��ׯ�ⅮylS��]�44�_��[z׬]S|߽��3 4k����v3*΄~�kB���SCO�k@Q���,�]@���E�oV���t������_��s}f�q��ZP4n���	C�L�y����|-�P��8�l��A!F�]�����5L^��<��/mm���:�A�׿��3�F�ܲN�������y������Tjc��S��t����tt؂���i�x#�v��~���M�c/�a���9�`ɓׂ2�c��mۓ�5z�g���-�[��U	5��ѼaP��xAh��)8��kqɇp���N�|-��!(���5�������H�9+��n:��U^1?d��LQ8@,����;��)ߙ���Bv���ꅺ�(s���	HT�C���m$�5�3�M@��W٣i�-�{�~ҡÿ��ȷA��x��[�O��<�6��ux�P��y������Ih��<�y�ʑ�Df��e�BC��J�������T�M EP"
VD�ʶ� ���
�5r��o +��B �ƴ?A��	4n(�%�H	�{�C)$љ2�((4�!Z6D��6�b6��t��<�j-��C���B�(?	DU�]0��L�u����1{A(���f- dL����q�Q3��u��{��\��LaE�zӽ��A�
o������_l��%�-�� ����NF@���w��*n����&ȉ�s}uB'r���H*�	:1!;}�#c��m�[%����#7�j^��#J��T��a{�{�Glָ��D�RK��=���0����AE�b�r�۳��<�d��J�Ẫ�&������N^VD}&�s�]����#� �	����E�N?(��g��a%u�R�nT8H8)d��hY��!4+s��=�|��I!U�[�uQU��؎ "lD93\3��+�RU6Ⱥ�B[%����喂�=iCH��_^����Y���%��#��8�H +��7z�����2E�u	za���؄�Ghط�B�-�a��8�̲����r�yF�pXj�=�����M�سL|�r��F��2�l	p���XcR:���oR{�n�~(�N������FS_t��랼TL��
�i�#�z�!���*[�	}"9�5��v-��ld_+�jb���Z��d�e��q��S��y�3�꣣��"$ȥï!��<f������LQn{.����"q�h���\���N�b��e�]�iX��e��
"�ѫ�����Z��+�a7	��b�r�Xfq2�ط���+ggͨ -?#�}����?ҿ!�y1<p�Cƞ=i\��&z!�����`��MW�ꆾd�q�#e�'!��2ݏ4��x{�k&\h�1�;��E�A�ʓh��{���#뽴,Q�pQ.�xZ��G�����������`��� ��X>F<��� 	���Ab5������l�r���KKR�7[-l��t�`��+��t�T�N90����w��[<���i�v��	�n̉�O� ��Lbo*��Q�f(?5+�؃ipc�i�?W\FY��0�
�C�)����!N����>���*�o`�C(��G~8��I�O􃍾���]m�7����r�1k�UzM��G)�!�NQq��q!.�e��>���b�(�h潤nE4NM����9&��l�ciK�L-�mꊱn�7S�d��"�m�����qOڟN�7Le�� O�0t��¬���EL;�������R�E�t���c�	�r���%ɵ}_,�G�y�"��!��7��.D�Lf��hh��Q�,�˴O�+����-�����;3f��q=�9��떵��%- !��ѯ�`��o(�_�˾�2��F�2:hi8��-������C;�M+õd��;�]l�yvA� -l��S�܅�+fI��a��Q݆}&�����I�ɑ��U������V�u0l6�
�ruO:eo��5�J�����
��Ѳ`*���0Z�G`�=Z���L]����~j����p�|ј���-��y�?�>�?4C��B'�0ur�n:yʢ���� gEs���ѽa�j���%���dR$�!��@|k�b��b�t������E�պ�����O���X]Ƿn��N8h���59��K Zz�h�B��҈�3³��p�1|���9/���?���Ve�E�B�v_?�8�͉=��(��s�����u3t7x�=,�sqv��@ ����jW+׳#%����Tc��ws듀�2>7�
�6r������t}�G�6��y�j7��\�:@#	��*`A�"DwN[��[jC9r�b���������N� ���� b~�	��n��]����odaz�<�r�m,��.��{7�������Лe����5�4'1��R��D���Ri����{6 ��}�r�Lҡ3U6��x��7�}mUƨ��
���V;~�U��Ȳ����S
�v�D|J��h�-={bo�����2�V�ʰ�[�с��q@���o)�`�ɽ�W�i=�Ȑeȩ#T�ǆ��%���C���}\R�βp&"�����$��H*1E�V�U�\�6�tF��䮈s�լŁ�D@h�T�{����kʎVa*���럳ȇS0N
���2pAce��G��F@m���eQ��"�`�ї,�dQG^�����C��/����}��<��W1.Q�!Y%
x��o׵�n��wy/�9�o��]s4I��oV��\�v�縎F��XE5#^�����ᚃ��3�������H��,��<ٖ-�Վvڻ��x�������[G�sLh�o�g�P��U� �kIF�X�|�I�$p�:��<���"��X��u�d1ZrgK��u���nk5�ކ��z_E�7��T���/������+D]J�X��7�^K}�&�p������0�u$��NEa�v�Ӂ 9)\�#�,Af�Dg�U�̉^��x��,:5S�� M�۴`��𮝕I�=�s��O�0�i_p���^�H+
�U�(���J�UΛ�J�}>��nKr�D���j��Nѐ
�~:(�|�Qx��>'��t����!:r&�jd@?t�-o���07_���~��zE4Z�tp�[�^{%+!�Wz�w���`Z~Mb|(s�����^Ղ���|`'����kQ c8l�h^�a�ZD��T<���"Ɵ�q�2iE/�tcKc?�\8Xל���tt�����)*7����ߔ���K�(�s���z4/0����}.��)q<�~���C&E?ą�P��s�	t���^x@�,��%&g̖MEIS �d�OF!�o}��G�&�w�)2P^��/2od'�z��5k���ҵ���u4gG%\o�a_�ܕ!:����JC�A؋
q������u��[�:�)�]�(HY`�o�	"��HtօRf]��:ц࿳8�@��И1RBW_�����<��-l�/�=��pa�<"	;�P>��*ϸ�+�d�>��<��Ӡy��@r(�@�N�Q};<8B<�UYV���;تU��d(�Nx׌�ѧ�7Xr;*ʊb��P�3#Av�=
�K;�Q�d+������	kP�o�3��=O�s�4���gu�A�K�̒����:�J)b`��_����p���T�&-g�]�j^�d8�+�(�}V@[�׻���+�l��8��Ka����^����V���&P��Ȉ@��tB}�f�DN^{��n�+��ƉT�څIi���K��������˄I^0�E�eF����oqp��%�o��u1�#H�y9����{ޖy���\�� u}O?�����Hl�:][*bl�^?C*&;x4v�k����#Y�����ԭA~���e>'I0̫O�?����ϲ��5\���Z �y�K�}��Gl�80[m�4�ڰ�1
�{E���uY�
ߢ�(�jV+6���?�U�z'7y~��=[_GW����V~k�cm���E~=t����<�w���c*����Kf} =q7��@|B���!�q���� D�p�O=�-��Y U��������OO���|Z�}~\܌r�	�)����}����)z�:6f�z�y�����N���9�f��5H��^"�>�x�jL�(X$<U�7_ �_� ��Y��1�^y�Vw�\�i��֛P6�s@Tv�Y���`����:�>P⸋@A���p��j���4�p�[y2���H���ښJ~��I}� s!��D\J�8��ȶv :�V�5�[_��I�2�['Hv������.�禂�q��E�\C�?Y+��u���X=��?�K�ݚY��a��V����>E�j`�9On�	iRx�kLK�g���7��Z;�0��N�;�޳Y�t_��J#� ﶃ��{c����v&8�kfܕ��.o]�q��������,�N��庙���C讎�ʭ%32΋ÃZ��N���'�]+/ځcҹ�i��2�����b�������2W�����b�HY�:�F�!Ϩ-n]��D�r�س�[�����A�.�\}m��H���6P���s���9�f��E ͸4�ά<8w�Y9�{6�%�rNQ
JKQk�\^�w�x���������{�Q@����<��8/x�9a���%�"B
D���8y��L8O�0Ka㼴�M�=?G.���m�ۍ����S�^��K	�$E�}X�.�k�h]�>�RS��5��*�p2^H㪉���j�m7�t 6]O/��>���T���ʥ|#�]l%7�5!Ћ�\�g���/��Rν�������m��ڳ��~��-�F�v���ł�� Π%>�D�����y���� � {�Ԭ\�4{.���,΂׭�ol����(�8����܈/�x�8��wHv���C�H����ckW`zQ�Х�������r@z�y߼|y�romD�Vq�^�ӳRx���ǛЌ(���<��B ������l�*s!�U�ʹW;��-��+٦����F���;QU�X���=�U�U^!R��>�C9dT��v8,�вK%+&���f�����M���&��<�2/�~Ʀ�#�k�ڸ �J�_xxN�E�-�o\�O��}�gIu��7�=��X*��=1G\Xnz#y�f�n1��.�9#��g`�}B�@�KU�snZD�����)��?�����E�����ApGM:�O%����G���䫚��)�y�T��@�
ҥ�2f'���G�t�	�L�k��d5�:;���|�_��s�A��
���� W5����0��	��S��&*aro�@o�=��"D���~Ց�MoؘA�M�6eH^Ӝ:g����Ш��z0�V�p[��D�������D�r�zd�A�j7z:vZ��x8-ņ���M�>��ig�<�9�H�bYGGB�g�]ǡ�i��SC��NwI"E��xq��)]y�5lx�c�M!;�Qr�.mz����c�n��߸�W�<H����ч;V
F�L+��u0C���~+P�ڂe�0/KKbx�$����%�q����!����q��3.�{��b�h���}�ڿ�Y�<1�t�\ad&�z�F��)��^{�A #5;PJ�d������Rg/���`�?��F��uS��5j��� 6�C�7[�^�4ʙѤa��,0�V�@�����?�hI
�\_��Jl�kT��j3Yak�nO�w@HB��Ի�Z8�K�U+�,V�$yU,��!s��8�#ׯ��&�)��4"����Xܬ��l�T�ɔ璢I~�a��f�c��k�'z�v�����*v��<C���y���D���:� #�H2��T8�%�����S�`�z�j�ϑ	���`w��Ч�'o!<4��z2��@�7n�s}�9�N��W��>�8�Ƞ]"� 
� �]E����Y��Vc�VȠ������?�e~)M�\>�n���%a��LV���*�V��	fۃ�Lm�Yޏ�&����lD��~�0�A��+E�*#�Vg?y��� e��֡��m!�Q���@g-=�^f�n��iV%&Nb�������.\/	ۍ���U�M�%]�ջ}�4ȫ�p,�st�nG�֞^KwiϹ�'Rn��c��+�/;JZfh�k+���H���wj���#}G��)�M5���~@+�:o�wNV�Ѷ�����?��=�G.G,�G�6����*1��6S�9��_/��&?W�.󱚳�8d���!~-JS}�� � �M�+����g�b���&�u|���:�&��H9eMשT�"sGIaG��T�}�����괔�m�y�j0QlpV}F�����{�t�V���O�<��.��̲�:�҃x��ڊ�N6��>H{	��k�����Z������i� ��/��l3녂AtlH_?�jM�'���j&��(��R�����as����+�ow�[m/�L<���8���(��ԾR�����od+%P*^f( ^b� fVЪ-s� H捴����-��9d��l*��U�����iM�5܉����R�:�r�W[.��@�~�C���RW�K��n.�?����)��[�<�J_�{���s��X�{�U����Q��b%��3���Ψ2S�
Ku��sS7�X��M���|���#}�ڳ�b�I&o�����ܝG�_�h�㦺�jo���ur��,J�?8#����K�	�N���vE�m!l �C9�(��'@g����e�1��;02���2��V�RAl9�s��4ү�D��k��cq���N1�"���~QIK�ݫ\���\F��TRcE�6�MD���2a�j�Q��@�s9��A�H�
,J!���k�mS/;(0U�庰�"����;��-3D/��6@ ����r�`�
��좃`��c(�Z�|}����
i��<�:�k^�^�&���;���?}�sdFW)
�5�����5���]o%����~ y����cQi��0�rG�������#��]����BŜ �(}A�B�g�#1�S;}�p�[��ܴ#����6+c\?�8�!F;b�M#�&Ēρ.fZd	���z��/��p5<��z���V���}8�&��SXն�q�Z�9�%i����:ҧ��ֻa��u�7�L�ņ���6G�����Cs˵TI�4w&d���O'Ƌ��IH��r�Y�M5PF�ȱH5zd���ЊL�c& �N�D벴�j���M�������L���� T����Y����"Ug[��Vr��K�KK�]���K`aK�"��kۥ
�_�	�k�{��HW�Ǽp��Qo�,�ȴ�T�����Y��*e�m�����f��b�;��[��mh��* �]r~.%Rd[m�ZGJ(����ߐ������%_�L"��H)
o�pkS��&^��LI'� �+n�pnx�}�<!D�K�z��{�īx^I�+T!��}f�o���u�|0�oY�Ļ�0�'�&��v���Uera�i�,�e��u����U8Tq�	��{���nB�FGJ���(GG�pv��ll�+��X�^d4�^���?5<�=HW&�f�^W�ڍεccU���ހ(	�&�g���4�]�s�j�){� ���N�t�K��ylo�1�x,�[�-��!�20������Z�&��>��pN�#�ʠ%� sm
�a����73�%��l^��Ǿ{5�:��?���
;�˥}�qDC���c
�6�_��n$� �Yo�#�F�n��ݫ��k�'�<���s���{28�u�>М��-�AGP��Y~�\��w�-q��!�n Ք9M<Ŋ���ͫM���˷q��O�K��يa�n�͒����R�K+����0�j�#���y~�~թ{�(��K۠�ڬ��"ܘ������ԭ��;~��n�c_v��м:Q��Ă!k#��j	*��1��$���סj�Zon*�;6㐂�n�d��2��ը'��r��Y�Ђ����:�-�w�y�\��`�K�:���'<���O��/�FH��1pu�S(��N����nĥť4���iCN� ��N�ۼ�FL������{�B.�}SF�y'�+b$��S�%�[��!��rd>�M�f�{.lN���P֐ٻ�+WʼN�^����'�/k/����V��A��z����ǀ�d�6���A�8���+T���K�IŠN63���'�eg�|�/�S\��b�i�$�` ��Y���qo&}@�fմ���r��������1G�T3룯��*��ﴤS.�]#�2i���(�D���I�&���O�%�͗�����mvܒ��j��z�h�E�N�bs�����V�bAߝEe'|��E���|� ������2����L@���)H�K,	g��h�ck;��w
��ɵ@��6�Zfu�T�S?#b*
pʇ���o�V�ߍT;^º��M;j��ʋҶ�����ē��c�cֺ�&��P������Ȱ6I*=a>̓�ц�hұ�+����2���֡ċ^Ӛ֮ z��ey?�(m:���1Nv�#�Y`|���N�؁����&�����P"=\1�2�
�`���/�������H��=�V��8U+*��:>�ɪ�s+�\#p�ZE� p�mN� -RJQ=�75u��
�����J��b����l��2iϩ؂[��;��|����MTN%}:4-��Ӳ+�*��-�F�@�'ƯG�E�E�⹤Yy�%+ bhh+݈,B�2l��32���KQG�`�E�G��p�c �fw�w4p������&l�Z~���y�WV;z�3��Ev�F^��)��)�M�Gk�2�+���Nx))2rX�hsB���8H���K璂�AYL<G{���}_g��機Tޞ���N��t��U}�,@f�S?�U��!F|��X��^���R\������00 ���>G���ZXs��.��f����gc�e^�iq���+�?�����%�?��h�N�3�2P�N�j���;�N��`I��\pN����0�!v��~6��<>�wH���D�d��[ض�8O�g�-���XER#��Pc�"Ա!�ԐV�X��ޛ&�m�ޘ�m�$���u�Fz1,���n�"��?`P�k̖�8ˀ=����\���}.lkˊ����;�w���#�w�b#�e��ظǢfC�Mo
�
��(ɬa�h.�x�k[����v!��A���0>�̡�́c���ߣ�t���`J�I�1�%g�]�M����Әb�ʜ$DG��?
�N1S���-�*��B�	��"[�U>ՋT�Tq6b<<4w�
�5�3�Y��S1AMdp�5���*W�Lu���[����w٭!L�X�����( ��aŧ+߮�(�� �5�����^����_7r�Ą�6z��5Z��Lq��vzZ��NR�%��;�s`{�w�w�x�xA�����B^:�"?�0�M6k�0�OP��6?	���<�D#��������Y[q�� ՚���C��/z�(��G��H5$���<`(����A�g=-
��k�}��������>�e`��pY��� \�ti펧�Tê*)8�#�Y�%��7��2��,R<���s�3�t���k���M�n^A�mK!%��jg�:����}�m��/�6�s+�>h��X���'?��C��E�#A��"O����,�v��7�I�=��* �#�d��Jt�?�%�p�l�a�I6�_T���Y殯�� ���_��(�sGZ_L@`�]�� �xV�H���4�v�r����_�jc��Ո1ǖ��!�DӁg�M��ʾ�-�y9��F�_R(O��z]�`nC�t��u�k?s(͍�sH��i��E@D�	�{��̧;�:�-��	��U��b	o.<4�Rк���&L U������ل�4@��������N8�ݰ"ZR#:�D��|2��{P���06�-I�ӌ>Ux.1͞�M=�NP���'q	�/�硏釅b��c�c�k�#�elr֯3�X�D����ƸE�w�R4^Ga\��E�ic�������1JT\O�a�2T_�U��sƃF��f�b)��2ep�fE������f*�3��h���Dɾ|l�ܯM�B:��s�8$S��
p�M��F��:f�AR��iȋ<�!,^�O��Z�	%�zv>[�t��p��9�/<�,׏?���KQ�a��"O �>��?�L������(�����4X`f�'���t.rq�)w�Z���c>��	�i�0�P��{�$��{�IŦf����@�ˈ�T��1�#Nd���bQTNRʹϿ͒�|��@��;U��fIA� ���ƜY^��?�t���` ;����/ɮ� ���&}��^�۹��F�]�����ԏ�\V�d�RGl6�
�<)��\���D��u�4ɽ0�#:D��&�b:���k�ɸ�9�7c�\�_C
��>��8��!���ۓ��ӆ�� ��cz�M�v�X�����_�V��RN���eBTB��Jbv�����s�'!w�ɣ�����_K|{'���Q<#�O:��?�,�-ui���!��C���l��D�F����K$8�`x&��1 ��n�VR�q�+�%��2ؗ�������qӨ'۬l����t�<�"��
B9_���:#%��b~�f�X��vj^<|��? ��&���z��� w'��.'{��O%q�x �3�q*o��ۡ	np�N	��zm� ���R�q=䐕����L����.�[}�$ܤ��t���^i��bq�0��g�wYHӐc���iߗ{t��)zzm�]`��o ���.͔�CM��ڹ�Ҋ�����}��k�xiu�c� �.h#L:�wa�1��[����*�ʹjT$h���\�����y�!z.F��JH��}�KQ�>c$�{�eAh�#T)]��\������V>F� � hM�<��΂����X*K@�Wxо(G��N;�6Kd&	|��6#O� ��
mX��]h�����ŋ,iOB��݄٪��F�%�����k�s�1��?���E�W��^�y�쁨iEV���y�a=�\\��u���f
,K��>CPyNK�) �vʹ�[NS��6�8 �ͻbpJ��4�-=|7���1�X"��a��gߦ8h��X��a(rO!U�CE����c��҅}�����_���I�g���+�V�� JT��z���[9r<[$�3�{�	1��u�h�zA6��\��G�	�{���,
����(�:�C��nݹ�(VT�^Q��|�����̒�C/�����5�������OL��?����� ��>	>,:c�Fz-�c�[�fW?�5}J}#�c�f����V*u�^��1�V�=�3Ϳ�?�t�k,5d�L��S�P �5�+v
�I%&��{k�x���3�񯭺�`P��.��R �+$l�8���S���J��g�(�;���c���������`���%���9�ZAI^�?CS����yfM46�{ݶ� N�
�����,Yg$�Qm-�W���s�k�h����n�F�}�a�@��S`�����6\.�v��Tb�Bл�d��2�m� ��γ�J(���O���`�(h�x��6W��Ȇ��i�����@�:	V��3� Xjf.�=,�0@���T0����h�~�%��8�Jk�',qQ{n��n����:��_1�z����M����Y�p;��ʄ(
Ƚ�C<޻%oq�cmAk�8�u]L�@K�>��2~�����0��L4W���uϰ�6�d<�
5�D#[�Z�W>�F�����m9����.���I%�z[��d1�(�;@g]г�q R��	�$����Q�I�I���P���&m��j{{W/�_Sop0��!��.� �%8�߆�͌ƻK�|�NF���߀����c��`֌U�ɣ��C�+#3h�q�,E�C�y����D�J���G�2ZW��Z&���r�b���O��]�%�2+Zd�)o
��0 �����>߭���Į�%6�:�����Y��CТ_�/����gǺY��F�GP`7}Ψ���F�QF4�B��5_����C'v����"�f���CS^��%��pi���ڰ40�o_@�W��U�أG���o�t��W�z��Kʨ�Q�b��Ј����'����#�ai���g�:���mvQD�>p�?�8t�%�X@�>��C�vt���D�dO8Pˤ�:��Sjp��ZË�
���r�)��]>��Z"�F�x���諧s+d3�-s�M&�;��{���XKZ����E0�H�]C���^f�Ma��:gu :u�*V�CBa���uӔ���n�U)=K�'����J��y��
���H/,���Iv;�z���.��v6����vG�������dK3��K��SIZC6�oq������#7�36!,�Lc�uXgn*kT�ɂ�IIܜsz�uڇ�U��*�d�멙�~}c�I�8�T��gQ�3��
�s=q�o�+�*T�T�3p3�ك���� ��Y��L'di�%r c;�	Mޅ�t�W_�M'�<m.��ޮ�Z4�:@7&;�b�W��g�{��MT�ć��
وF�`$���1�4}<��T�2��G���&&,jQп/�>�M.�V����m��d�;[{��j����t�*���[!���bF�i�Փ[�%�{�-�?���Wv�6H=[yY4�P�[=��:=+��V.��P1&��C�>��n�vZ���8���x�L2A�x�]-�\j�oi�������9�=�e��\�����@�]���͎��{�]m$���Da[ǭ!�n\;�^��5m��[[@-M���fǾ�j;�Ҝ�eX�b��3s) ���\��-K�riF��"f�����g�ߤpI06�' ����SUZYC4����S&9�ly�8�>0��������z`���2Ln�zs�|���p�`���5H
X����o[����Mf �	`Xy�@ݽR�L%�]��ޒ����;DT��R�Z�����K��ڐK���L66GN��.g[Me�K�����0s��~��l}�p��;j\��[s
�Hr�?��Q��c�UR����X�=���t6l���~x���s0 MjT�K�]ו>�3�A�Q!p/�N
��3_��6	���x[��nᮉMfT{B5�ƄEܰ��k�;?dU��l,�k.aj2%�����X��jBiUE��:��;�z��������(�N���g+�{���U!��]�ʞ��Y�ֺv�}�g���;��Ǯ0�l,<q`��;��f�j��u� �N���ͧ �+zA�N�N��	��}���X�Jҗ�����o��L3��d0S�*���8�GP�;�O2�T8�\�͵afD�������G�p�H��,��˫��������� !vl�&.˭q,�d-]��CGGƚ~c��v�3�T�u��Zk�༞��b^C��u=1�
� cb�b�V��~(K�q�sS�j#������zN}�"̈�6�.�3���R�T�H�Zg�H�;�hUI�RLƠ�J��opI���by�#yv�7��C�$}�!{a�+dy=�V'��n_��_��v&��Ղ�p�:�Q�1f��q�^�Jc��-X��-����eϏ��8���b�lήb�6'�!�b�k�͛*��+���f[C����3T�Hd<m	>/�*&r�x
L	d;����TMR����P��Ӻ���	9	�zD�ɚ��o����%U�?V�!2)�o �q�����-h<�����y�K֧�$��/VUa��Ll�&����ainX����k��7�y�T��x�v:m�#��V��Ȟo�۬F� w����t�s�:�1�{t����m(򤿒����-9{��oEN�0���&�e��D+'��j�������X�)�rD[��rB�s!|b"��/`�`�v��	#1���q7=�S��a~�,F�6��푢JO=(�S�#��[Z@���B@q#�ǝ��a���]�Q��N��i������G��~N;����;8k�~�=%�����d�܌����!�b��?$�9�y����x���F�,�;bύ.�ƨ<3_r�z�nב���v����Ş��Bѡ!����wX�c��(V�b�m]73{��ϻ%� C�M�Tc~���k����P�l>��ۛ�ӄ?�"�]��e�"w�"�ډ�j��'/�V�y(�\P�BB����l�-h�?j�̇	�Iw�Ƒ����
��&_����r��D�C��߸v1R����e�uu4�DA13x�����g��������?Z��vg}�:(�.uʣY�b�?P�;xÞt�HA�-�*J1��S��H��I����N��ʆ���"�����A�qr��OZ-��K��Ҽ�yݑcF����8����8�)ǹmAk�x��_#QB/���,�O������+wf���MGd�'����=n�0�1$�˩�Z�=䢷�y9@�EP1.�J���E�M�d�R^od��M<�����M<#u�|& �=�8�V6�ʂy�i���#XY���;���~ǻ��s�����AT)DrΛ�N.փa��j3���^�"6=�w��Xo�7�������HDP������ȫ����4�0b�Fc���N��~k�ʇ�D� y� ���er�Wk�s����&������ԍ���u�ҥ����!Lq]rJ�%��x@���3l��xgZ�a������v���m����Y�a� 4�h���Yg��N�܇���A�;h����	��QY��_�H�I�xp��J�����(������'qg�E|w0��v���X\�>}@�(�>xE�V��'(��]:�Lpb����@�u��;H�ē�ɈY6N��U�9��=?v���n4`R�$��i95M�7�2R����P?+���>@^
SI�H7�����᷂�6袸��V� '���s�x,��.	�||�ˑa&˂���|>��@�g��RԠ,lC|��_�P��z�<�N%-��g�n���5��
� ���U,����˸�Ô�oHg�j��zk4�Ԥ��@�[ZI��O��l���|/�KF�����%�g�ԘvC�K7�ف�IDx��;���n:���`�l��أ�t��0{z��XCq)�q7�������fh�/�S3�����ਧ�t���T�]�V��h�	N�m�g���e�r�(x��H���(���pQ���.�W��]�8��^,,cҾ�Q�%iU�U
hӹ>��7zb�2����i�,%'{�j�+�{��[�m�j�#o�u+�q9�	o�t���VAć��n��v�?u�7��_�V�/-a)	J&s&j��B������*i�$�-!o�~I�#\O�5�����E��d�"��kt%l���T{`�8�Kߘ�U~_dN��ۮ����iPr�����{w���#vK�=�ޥ�j5�i���sKS��ZOx�&�M����%����;�������XFp��e*��o|�,ƨ�~����,��ݓ�Ș�W�R��D�FV�׳�b$ޘVx�m]{zm�[1a���~� �W�뒤\�O� V��m>-�,�,��T���J�iW�gX}T'w���3��ӆ	���&���U��ߓ-�:R���F*6�|.�O��l��/�-��Vyj��ee����Lha���)�(cL&��R,�$�����Z�Ac��r�A��ڸJf���GPKY��<k�s�w+�^���9�%�dJ&�vh��	M@R`�Z;��O��"�0򷲭R��^$$N�����c�������kY��d�oY��{��|1�V� բ�1��4'��Ul"�?��.��%d+=�pW��]�R�/�_$��n^vѯe�Wg��+��)�[�`�8��w`�1B?N���.i���xg���}��v��$[�Y����to����*����n�v_\l�'�:%��L�:kK��F�b�Wz�QH�Co�F�q��+��"ǈ�;�!č��[�#��4�!�E��Rw�z��t�D^�S5��WM���A���!��o^��Y���1�lC�?�^͇���0ɫZBc�1�/G;�T�~�����'|ʸ�,���IO_ �8[߮D��cmT�=��L�����_�}���������O�Qv�̌�\8�}2�=�ڛ�	0��^:*a���J�Ǵ�@�}���9�*C���6�!p~Ļo�ECV�C����#j�+�9��{��`7z�ST��h
?�^�Z2��pϬ�F�=:��X��������_��N�C�o�eo��f�뇓�	�c�_HI�˻�cc���S�����9x��(�7k�B��i�lj5@Z��E�v�G�{J�P�	���X$�����*D�j��R�ϳv��W�i�r��®�I��ﴨH�|���2�T�uF㡎�y[�� R����F��nSt`�o�5e���~��-�ֱF@���
7�ܐw��
�翄����[xk:�Mحs��<I�j���0��:�n+d����˳�����Z�UX&�u^�N���Q��n�T�͜X�P�����m%��Q��s�����B+g����%X��t@���{�&:�tz!S^��=�B��34��7^�oYRc�;���Sox����8��J��^��5���ƛqr��N�T5�8�8O=��U�v�Q�P<C?�G���>�:-"��,>[�*$X/u��Q0{�Fv0.~x��1xp	O��u�kQ��
{�y��:��Dk	WY��Z��;d���|��N��i�<��� ���9��f�y��iA�^^�ȫ��V�`_r]���YeO}ȫv�7Y����&?�Π/��$�5+�ɰ�Z1W�T�$ɒ^ ':T���s�F	���鉲�fri�����^k�k묹N���gN�#�M��˫�����A�|$s��w����R.������O~��~���C��36�&���ɧ��_�����]e�?^�8�XݠiZt����uM�����#��J
>�&#&��V�lf�(F8T��r)�"�b�	���wsH���������KG��}w[��r�Xv"!�;Æ���'���]�������Nv�E��t��RX�s���E�x��h6��W��Ę�S�P�!��Z����� \[���o>!\�~G�k�����:�m�S�D��s��r*p��l�A��|f��[Lp� ,�m]ڏЕ�:<+=�F�*ޢAѝ?\��4m7T4��yT�8�f��߇n1���c��.��[z�KOF(Z�/w��O��0�t�
p|$pKLE_��\B����kߩ;��b�!s��[ևw�m&�rY���D�d|�jv���F$�b�r�ON�qO��TS��i/��VIg!���*�B�+9�����ǔ* ���A�|��V��_�dd�s���<���һ�XG�	��y�7�i��'4�����㲓'äM*�+�K��D�c qR^<h?#V�[��	�I�}_�Y҄�����n4���0���8��u�Ґ��LA�6}�^��br�ȳ�؃5��=<}��1�l��'�m\T�.m�zI>�L�������1K=z�8��K��ɲJ֞n�
9hbR$\��l�%�����Wg�0�:���b+@iT�ڭ�n��[�Y/�u���g��!H�f+�����y�X�W�:%�C ݤCM޷r�0�A�� ��0�_�O߉T�QU�����Y����ׇws�FY�|��+9�r�Lev������7����`� 9)eay��ޑ�`�*�ҎE�V�����"(��G�&a�xs�pH(X ���!�N� yXn[�����9���~R��$mI�h��x)�3�y��9���A5���1���:b�=>%�/c#�34����,h1琑�����`/.@�C�����0F��ߵ'�e4n���k��1u2TK%Z��:~�,���w-(%u�i�(3:)�ws�$_kp����LX�J�:Y�Ǩ�$�4Q��v&Jf(r�wGn%k{� ���
8[0�����˺C�LK����DWJ���.��
�68��#�ǧ��U&��)��-�{xFBja�h-T�/V`���kU��~aCc$>b�/�mH:w�ʬ�c�IC��*e�H���V�5�	�<+s���@�9�T�n%��ۂ�n��E�[I��v�]���x%�g%�1�/�*�g�����Y�3�����V�`�S��3à��+�M�ɪ$���I!le����22�h��:Ể�u#K���6F��:RlW�B����`����A��E�x���ۈ;v�%�� l���)pD�a�vV�^V'�xg����
�����W��I8�--p�{�N��������2��Y#;	+oИ�E�`�o �-Z�5����#w}��ks:ܞeaC��J_��<������d$ilxP�ܝu�5t�{�A&4L��jd�=�"���4�wM����q����V�t��h��z�c��q<vE+��*�ZsEɉpl�.R�rC�'T]�[��K��{P�,�Z�k
,�<�_؞�:/����eл����Zj�{��Ӌ��:\]C��#%�c\v5p�,�ٍ�@|sZ#X��6QC�m$��� F���&��f���é�t�����뎸���T��0M*�*��P��?��F l���mI��YK� �� V�׳��Z�����?���b#]
��U:-I�u�B��4E� ��t�F�D@m����'т��n��fb�\���͑6�p>r��Hev��q��M1P��/�&����mshI�}��N�m��%���� *��"C6���*��h�P��!���a��-�����,��鳟�ʨh�/�WP/?!/h[�N�xFXK��Y;�56�Hv"�F��ޕ�L���?�^ ��`rGbވ̨��b%���/,<oYf�m�V+V$w�ߛ��E�[3x��`�w׸��AS�Mimp��C:� �l���+;��9�~Ts�_���	���Ѷ���ң�H ����(������SǪ �Def���*�ܿ)�����z_���� =��{ɺ��A���de��B�s���q/���Kr0�IfX�h�HCs/�m�n������4%i��܎���Qv��?h(Sz�xQ�DTnU6��*�ʡ�7p�量��S�l��5x�p͔�e��([8T����>�q�M��ZY��q��y�A�R��V+хڶ�D��FD����u�l��;�'����$]��aO���٥;�L��_+�C]�� �G��t5��T5�F�m+�o��&�o�<����53�$�0��%V�s���(�v�͞��#d��Y�a,����*��_ʸo�m���t���Xir7 �j�计M��!3�#F���T�����;s�,`r�ߒd�Ǆ=��9v��F��-QO��I�$�֬�HJX8{�M��\�O^��c�����m�#�PFCm�9���'�&�8A�g\T�=�����Dn�ywG�M���:2-�=�ʶ��\��|�]��V������w	N����e�QG��?��.h�_X^��$�Bkҍ�^��bM��X�������hC𵱹��=����-n�aYgJI�ʉ؟�v����y����������e�*]Q��b���ȅ-���[�U�f��5u����D�J5#1��;��m�+2E�(���S��P���T���21c{GC����{��{�q:��/���\�\]��]�1΀~x�p׍������<RB;��f���D�D�R��8!��n�ۣQ ��i���h�ʌ�K��uN���q|p���R�&j�y�uY

޶�O�p�8.H�	/�Ҭ��fsN�Ǟm�l��r|�{�ÛY2L���ƝJ���DЁ˃=S��(.��[�/�í{���Gᙵ���̭�ﾘ"p�"4��Ԣ )�5�!�8^�3�6^+!Y���p^�*-f�V�~YmHt���3��!��t��S���#Z5��\�^0G67���~�ٿ�75y�U��Õ��	S��
iw�(��v4-�{�ٻ7�S�^�6�u.�M�@	�L��|��ˊ_U��L�}��<�ʿ��u�CsÛ�n�/,�i`�t�{Xq7ր���q��&�W���Z!���B����̧��a;��������W୞f�QW�L��MB�Λ�-�݈���.p���(
�v�7����"�S�nB�#�9��ԁ�3�(mJ^fڷ�����9�4l8����~��.*�Y&�	��3e2�;��'F�f��jZD[�v��Qb���G/*�M׸vk̞Fd�c�A�D;���}�����h�|H"��B\ש�Ɇ��Q=6��\���,4MT��
!IՊ�?
� ��.ov���'�j����#����ܬ�<_��.�_z�Í3�XrM��h��h�յ��3�K>e�q�~1F��*�ת�v�_�p5��k
�"0������2ft�+�o�\7?�Թ�,�@t��L��$y+�L*#<�8��x C�=\��D]\��Bo#�x4��r�Xd�GfD���f�&h���3e�U�n��}��&��\�P���L��yU���� �
\��!D٧W�S����]�N�کó������U����������$��g�?�B��nj-� #H���h-	$��W�7��?�c0����Oe�(���R�x.B�5�g}��%�0\�৹��t���-ߣ�Q���dh��и��ʔ#�(T>2� �.�s����[��a_���N�:UZ�7�h���ar!aݍGҢ�{���`��!�2J�(�� l�E�K1�aQw��Z�1��[��s#G������E��
5�"z�֪��=��_�.��PCͿ�F֎�k�k������6����T��ϭ,9�g.f����E:1��@��/�LM���[�ʏ�Nᾤ��0^�$e?FN�d�K�;��F��N��$;�t���l�6����~W��@�8�� %S@̡ۧ25��M,��׬e��B.�e�^�ө������]4)+��,ӵkB������|hg�#�ۀ}֯���n�1qN����o0� �bm��O+w@Z*R������C)͘g�9��3L+�����`G�n�
�F	�'e�>���C|V����i�5�\�����bC��g:��-���q R��RUfJy/��*|]֚�����Q���6s^+;d�g��̞
H3��y#=����I�r��pp��mU^(�����/Q���8ېcf�wA3�����Koϔ�O����iryi�x21r�^ b�V�l���3[��|���C�W)Y"Y��Z291�m=XK�`b�Ew@*ܸ7�~�$�UU�=�|W8���n	���SC*)a��j�$���
�6z*٠% },}��9_�f�D7Nے��ڀ�� 8�u.�y�^�q$��N�>L��J�K[Em�MhE����[�z�'�.����M��^���7r_̨l����ZM�J�`�?�,�������I�b��(f�uY9P�����?�NMs�Z3� ���������9�O@���TeH��}�����Ŗb����3�k�GA�b�ˠ��9O?��i�B�&Yk�:����EM
w�l���zB_e���g�7�Ny�D���^sҢ
�e~x?�E��3S�Pr lמ�/��ݶ�*C��7���ɦ�k����qk��j�C�/����|r>j89w3W��2I0Pѕ�u�n�Գ�h�L���d�P����U	�[	2oߏ��+�-g�9uK��(��"?���i��U8�*s���v(�PU�=b�`P�Q��@a�cH����\ь+���|CѴ�/�?<*c;>�F��ڛ�>|�''&���8��K ��θ_4[��a���_7��M��i鋠���-hX()���ߋ�,(3Y��p�A�gv╓O�{a��l���T���g ��G�hB_�Jd����i��J�x�i����Z�.�*�mE�眄��a��E���P}x�y(�n�.�)�Q��ON�����8�n*J (�2(�}9�SOl���Zwߗt�� �8��(�wK÷��
���,G�K�N�b�S���j�|�wͳ�";����n�\��A��(�W�Q>Oļ��>�����J ��9����H�0���d���q�ʢ��K���F��LEy���(��%��Z:��Q��~^�D1�!����9��l��_ �dW���ӗ�U��(b��� )�uN�q>|���=��6_YG��9�:�!�a��,-�]q�˱�}X�po$I�^��t��pX���U4�U2������-��^6��z�I�9������`�/v� ?~�|ɿ�0!z� ����4�����0j��:Ka����F��yU-�e����[���Nh8�����)6�b	����8���]�|W4U�9Q~4GH�kǬ%�L������o���L3V�=Enښ;�_���5�<��퉩_�oG���-���	-Z�������eE��o�zc,}��Z�o�E�m�A$�6�RX�:�����0������a'3&Y���"���rЭt���^-��~Q�*^Q�s(k2���<�ڈj�	�#�6@ޱ݅�<�R�K�w��J10o<�[��������%�Z�RVvJx��r���ww�si� �~Wj��)��΂O�@�<؍��rD��_�Hi�?���03pH���ϸ�6d��uQJ.��{����,at]�u��L��~�*�sU0��eo���5f��?�+U�L�
��rF8��T~-.܅�Ӯ���H�N��0�9��s��cd�	����g��b���JA1Pp�P]��)z
���>\�yd�5�kXށ����L�i�,8Ϛ��8E�̓�AzE�u_�I���w,�>�k����V%��@�0���+���<�Lh�/�>��̩	�r�,�A�,�C3X:w�&T��/R�z+uy��5���NK�9�(����h\�����R����/oeA|>�t��c,�Q�#�ޥ�/�4��FQmW��[�����c�!)0��6:�n_~$v���v~�x6>��r�[B!�Sq��-��1���(u�6�� ~j*I�	wb�%J��2��܀,��ҵI��g��b⶚=n_T�Vj
�B�B�F{G���(��I!�[��I{p�ȵ��̛.�����g`;d��_�P�:�ߧ/�������KG2��y��3���_�N7���:"k���u�?�Fc9:�8�a�;�I0��8�>(���=ޡ=#�;(���V6��q�εtY����`!�87�rx��$[J�)f����i�$��M젍-%)X�q�L2V	Iם�>��{ư!V��)Aa�r�B{N�3����s�o�*+��>������v4X�t�G��
�s��&@�������!�E�#��"�&<ҽ��S� NB�T��eC�샍#��
���5'a��[�)6�Em����]������W�a���[�>vn1��D��g.�F�q�z:ʈ?ɷ7���Q�A=�Ї^Ur����S�z��{Zy�B�q��P��~g�D��ԧ�q�͂�iR0~x� Y� TūG��!��"B��Fv+~E��E�{�s�2-�wX�9��ʥ�^<O�v����p���d;�����́�.����A���z$�B6��z��c�^	�uN���`���g�Q���{��hr!LU>�TyXV7%t�������Q��WvO[Pm� A���ı�G;����jy3���G�a6B:��E��?b��\�y�r������������
N����^nRݳ/�MjÅ� n���8
�]x��W��n��j�M�O;�����N�D�>�lU@J�Ot�}幵�^���dN�����% �ʆ^](T �1��`������倩�#`�`���
�޶/��	�Ț���HR��8-ߧb">s�U��!υ�{���O<zlTN����$3O#���I��|9b�*��Q	r5���	