��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<�y'�I�z�OB�N��;M��������die")5��ª�w�r��XO�-����m�	�~����H�z�.#��;�s@j�.�eU���x�:
e^В�ouږy3:�#���/���6'�սc@��эgW>Fc�=|���)�i����c:�TF��zh�sh�
�(d����Yl;,��u�҃Z��MZ���\
���i����m'���j��퍹��^�b,(n_���:�3iA�qЄ	����],K0��qJ�8c3��aL����`�Z�k2|���7�R*���^��>��y'h�K���e;�Lp)K�`)'�ʧ`�:�햍B�7������P3��^']�\�����K��f7�E,�1Q)�oH�����x�KC�Q�Q�#R�ˑ���<dc������d��^�ːiB�����W�wf�p�T��I�nw��w;ۉ����|zT	���OѬ�U���GS48��p�	�x]ހ�z�F�286����|�����?��B���%�^jO�[�?U���k�#C�����+��?��K@�F�g>�f02X���4w����h�V9[A�l��xD��̠k�{�lX�q����F����9�^�$e-]3� 9��4,��Cp�l� ��l0�[h������cU����k��&�`��H��ᑖ��p���@�a4YHjr�p�����AJ�I<k*mN�2�W6v N3rǶ��}.�����^��PK��� ���\l0��j6I�D1pQw,��^ᑯn�&���`�y��Bn*ټZY�5/�QA���v�{��gm���w�m�ckN����c��7s
e2c�]�!�3:�����c*#��A����@x�(�;�Smb���e�B;����6ߥ7}��%x1���ēF.%m�w��?����ϭ��ք������6���}7���_K��;f����t9�������j�P^�K����\�sU`˗�/������9�b?b�	�m�����g���N�����e��)n����9���`��,���ӂ=-+S	��r�[�n�ȉׇD�nuȉ7�?G���	�L�zâ�T2�o��:���t��A/� ���[�YCz}b���w�`}TZTOK�g6��#����ϔ֌X�ܱg��(�xk�������']�-"��.;���b@��
㿨�x��w�-W�����)���kْ^E`�p���O���U��ٞ���j'��.F�������2+)���Av����%9V�#w��!��d�q�6��9Z]ͿJ��A�)/B���BI��,��w�&�>8��6��{�r�%cb�`��� �sg�G��щL�+(.]4�}q.od�YՑ���U�< k��	��-�Y�X_��ۉ"7�愷
��[$qd��w��b�i�Rt�q�챔�F*�ju<�u0u9Q��C����M�Ÿ�5��둲QyC�<Y�G�`�EPnc�'m+�S�,���;�����Fu��	w��m��6�}�%���!%u0��.6�B˛�y�qt�NL삄�P��Ŷ�)�����Yey��V�O�Dt�z���sڎ�S9�Nl
-`E7Ҍ�MO�۪%��KN��S7�2.���a~��4�v���f�W�~Oܗ�52_ɸ�z�������Y<�B����G�5}R���<멑�0�N�u��ٲ�����!����\����-)�0')�z\bv~_�d@��<5-X�sU��^���'Z����83�YE|2S]��2�.��f7"��'��I�%v�G��*�ڪA��@�����9�	~��N+^�_�͒��t̙P�}� ��6D�e�m�K���A'�_ fc��F���[ 
����n+�Ђ#�@���3Y��^`v}�vB���gi,�#K���h�!w`��D3An��ّK�K�%5�*�ܓ�x}���R:�}P(+TGjDCГ���f���` zz�T0�J����� ����Κ�B�?x�D��HD�H�ׄ�c����َ:c}���]칔n�,��z?�ßk�M$��}��_����:��q��?��7
�%��"��-ŷa
t�hO�FE�[����}���fta/��\�V�%�͖A(�7�hK���_�yܖ���P"�H6����V�Qr����ro�"�������a�ָpH%O��O
�0R�ڒ����i�)k43�f^F�W��t7�E����	�������rsW�Xk��>!_��k�s��k[X�5E�>��YEo�IYd�r��D3��b4D�W���)T¼~M��f36�ܑj�gDK�ok�l����9���G�n�O�k����@L�� 5��F�~9�;_gŠȀ��r��j��"����E�QPJ=jkD�%u�دڌ7mF�`Έ����jh�8���`�<���G{P��{;�RlEk?J7��H�)�n�M�t(*��43_|�EA� �R̵���`��J�r�{���򎨜 :��W�� ���U�KH*�(�t��jD=���.5���ac�dr����>��|@i�Ǌ�<�d�ЊIT�����l6�G'��4�,�5}L}�GCQH!��Q�8�e�]�}�kޗU�N�R�*�>@�c�;[�q�� <$6���tش܍�v�ۑW��\~�2��TU'�W5!Å�|��R���2�<t(����Bf�+�+�۳(f#��g��4Uz��p<�!K�leiYNr���!Es�.�1T���W~�Kd�����R���ȇ�.�=�M��~��M��$�(�aa�>z(�^��`��6V��0����"��[�9�0s�7�����(|S1� 	���B	���+�U�'2��{+��ƍ��>)�	 ��Q�=�{FG�����Q�J_�ݧ�˝���8�p���~r���u��e{۽ú�-@��D�Us9���S�u��d���!�^�:ľ�ݻ���h^ ��0�ut�vw��ܖ����v�]T��N���%�oprF���^��hV)á���|�����C9wͽ����ʺ�u��G�ZTb��n�d"j���F�ltr�a�VO�H�V?�@U��ºq ԧ�-�AG��	r��dg���K��|�/_��>�X���$�>p��f+ќ>) [�G���8���ʰ�_:��#s�U��̽o�¹ā��no6��|����X.XX�����(n?g[xtQ�
\���v��]G��b�������;Oæ�����}�z�R-y���f55���?H�pݸ�nh}t_C��6��gE���\���\�#��᠘w�:�J�`��3�M^q:��Y��)�o/�I���5+f��pQ��̗�N�`#M�}��l�g撤4ꋧ�i㵨�~vx����Q�Ȑ^�����U��꡾:��z�\F�v�K���?�`�t�(	���I`1��AƵ��T�����$�x��z���iH�h©��#�>l���|拺݉��xe��h��U��p�ڸ�RUP�~nq�K����}qc�o�j�a���+S�ݯ��,W'B���N���z�I�}���I+N�K������\b��2Y��}�I��g�^ޚ���;,���Q������BIk�]]��@�������Zu2[5;�%�\��p�2�,N"?V!F�Kar[#y�&3]Aٷ��ҖN���(E�$�@ o�>�K�1�6\R��D�c��=�tc� ��EK�_�]>����<!&O�'{-�u��_o���n�N�9�� �wcԶ��8�fGD)��i�&6���^E7_�ǎJ�t,�$g��Xʼ������u'�˚�铜��J`�[�E���͍E��,IT�����>B�v[�,#3�<eV�ⱋ�4o8а!���fH�_��}@�%��u��B��QS7S��1�Zy����tR%0���x ��i�,���Dw�ç��H �Y��:X��Sbx����\i�'�]�cG0`��i���-2�����F&N���d �=�L;T��s�@�B�*@WёQ�R��T0����C��0���`@}%:��I�%ͼ=���M�F�nX!��8���;.�]�X�IY�U�Z�a�����`�ɫ�W���'����U� ��/?(j�A�L=��e���qm�G��k9�{CV�'��F�肶fI���g�	���Uvv�.�� 64P� ��`-���;�)����/z[� o���ő�����I��j�U��l�f�^�����\|�w�";\����P�L�����wW��Wv��¿�M��{bo�;8�3)
��>#���qA0���m�%��GGI�P^?��)S��E�EK�sGݟT�����2GMz��P��󸞌W/���Y��7lLw��۰7φzS�O��^��y��çX�Pbv^-�j`��EK
�Y��RR�����������x��i-5����H�.gJ���g-k��e����*�� +�!|c�F+|��d�̷Y�I=���t�㷴�7��,��- �uEx.����|��2�I&�w���n�Gg2VD��Yզ�������Y"���>G_S���>�M��x���J��ǙUI5��q��qLW?��4!يA&d����x�&u�1�%���Tc��g��1Uz�'�5��"���A9ZaY��xC�!�3��}�^%.B���C��y��R`7�=_���.���]�?�78;|�NF:�� ���A´tTgW��v���E*g�I*��e��o��b����|�8��8�,3OH��3Χ%f�&[�����x�_W9��4��9�R��/�R���D�;��m��=�`�;ڝd=����:�>}Kn�^_M�n��N�	y�$��47|Sq�EF-��A�ы����O�6Üs���>jo�s��_�o�?F ����!�|#��XP�8ǂ>�� �5�4z���?I'�zw��IԽΚi�3!�dt��N�4�N��dړ�졆4�H�u�C\��Ӑ��4u�m���[������J����w'=G_FcB��a��y$>7!�%�#hE�گ��N�������~��9Ϸ�Qrў�f��c�	3C��l��i �]93�X��M"iN��Pf6 �!uWW=7OM�; �K��Z)��Z�6	U@`�����o��e;S�G���h��oҡ����^�'=�F%�!���o�Y�{��#F*(v��u^0�H���ND���5���G��H�Rxh0K��Ս�~4V�
�Z�q�a�A�Ջ�O�0�ʀ��2{��+�+#~��[?Y������̓]5UR�i�l����aM%U8�P=���9Ҍdl���+�X�Wlj�{��1kh�5|{<x��V��g�*$S-˻��s;R�sЦ��L�nci���Y*s�e�H$ޥ+}�@H5H�oA>WH���VM�o6�L>�WKw{��d-hz�L���y�2Ô�����W���]����gMĂ�k�6vY��l^�t�.4���r���X�|s@	�l��Ձ���E�멧��<s�F�`N[�:�A�/L!c����l�T"4z�<|aB݄�V��C�Z_m"g����:�d��^,ei�{x���:�9�Z-����Iu�6]0�?&�����mAq���I���Ɯ��Aմ똿�E��%�$���Y�!��͏��DF��Qi�)�(���
��G��7V�F窋B��X\A��&''����QR�T|(��&r!�}:�NR����lE�~�Q7�D �&���A%�O3��s�y���wq����ׇ�$L %'.��l ��w�q�O^u�g�y��[�=8�����?�ZTd�Qx����EH(l�B/�>��`9��^�K+6���d�?�l�.�m�%���)�.r�-�#�hxGk;�5�<�L����a�ϸl�������N/Ĺ��%�L9e����V�;;ݽf�Q��p����dw�\/����G����	���N�n~\�w�����@L�2���-��)�Պ��|ܸ=�b��+�;�H�F/��Ed��*���n�)ź8�:Y�w?��o��c/���oz��θ+���h�9)n�-xFd�z���҃!��#BA�q�@�U�<+�u%�~��G�I��<�씃p��s���jŀ�z��U�:�4���z4X��s��dp�!�ςb�[x�u^>=�X���z^����\u�;4�j1������*s�O���,���0�5DR}�Ri��4�e�<u�W�%;�c�*�7��V�C��A
͓���t��;b�3��
N�Rxz�9���&f���Y��������ƥ{�����}0V2��@4
�~�a6$����C���2����N��/���EѰ�̯��P�Uv�2�S]���(�	y��"ǊK��c>H���6��4��G������{����L��'�B�$�O[���{��2�Lw���� �yQ�&�[��Rx�����mU�d�){�v
��ߑK�W��RɖmnGy����R�0�g5�r�������,8��f�J��(i���\��NU]���8��,��g�����y�����i��\�X,:�L��̀?r��`[Qbs�E��@��h��RP7yn*� e7�{�T�@x���)N�Yꈁ�m䴜X�[ _���$@��er��� [%��n׫!��n�F-ċ�9)]/� �x̠��Z�I��ϸ�#�^�Y�j"C�x3�`��%Zh�[���a��!�i�ٚ��3\�O�F���������q\�ܨ�����H>�k�i\���u�2H�Ĭ�Zzs��C[\R������c
.�ǳ�54�up,8��pxf+���*Cu��9q̼Cv�AO�O�
��J�m��޶�.��Ø�i�ϘЮ��(�H�p��2���|�q.���,^3&�7�'~yPf��\:�v�0l�	ܴFߎ#2ٕZ�pH�䎙qW`�kXY��LMp�'��,�q���E��؜k�<�̞���;l�!�^�&��|qr�kG���@3-�6ʲ;��G�n�d�7�.��-��� ���*K3_j�� x x'��7�oJs_R�<x�	SX_���H��9�Myl��%�9�F�P����ڷ��!��N:�>�U,С��� @-W���}����+4����7$��^Kqn���:� �1-8���Enu;�F��臛b"��8E�M˥w��(�O�p+r5s̪��5�Q�̓W>��ߟ�֩�Y� �Ak�D�`+�o�F^�&�s���U�z\�![������[D	w���/�����V����\�u��@4Q�>]cj���텉ٽ����bWY�p�����5�3�I�h������$P�`�f��5�*Wn?���4ũ��W�������pC �v%`�=��̔�N2~�f��.����Y�ƕ���:ߗL��F�K���J���H��}Aw��ʁ�PJ:��8,vC�:��c�3��&1�H�!�92���P�bj���Y��u7LJ�EI�ؐ>�ln5ʅ�*"5��@�1��LI9��d8$�f=L�̇D���۰EJ�%7}^ɻ�M�f���� 8<��z�x�����M�C�����l(���=��9�G%g�vPua8�8l�v3
;G�-��H,t&��ϻ+=\�Fr8<%�ū`�M��;���11���g�1|�,/Zo���O�&a�(�b+�r��C���`�(�O�*��~��ld�o.�Wy��w��J���ϝ�Ͳx
�}^��J�hj���#a��П�&�q#���9�mp�ǐ��V���n��U�2����d��A=�0��tB�~�gV��'�;Hl��]�7��b�h�W���ЎVE"0 ��x�K(��(O-�R:@�l��M#����w��<��'�(h�b�M鑷�se!U�t3.��\������!��|�48��OZ�@�Ȇ�5$ք���ޢ�%��<�a�'���dD5�SĽ峜�x�f�k˓G�+��9C���(�MZ����8�������<8{){k\��vx�����]PItS|i,.	�(m?X×����I�<�]����𛪠�w=�D����yT~�g�}N���Z����UkJTQ%�:%�Z�ı�-�.?0�X�˧R,�sig{}-����l��s>���t���ȳ��XM�O6£�� �J�J
���3�=-ApYRsݰ!�w��wK3���D� ���_)
 ֘�)���s�!1��93����G4sN���P��������v��.q���B3g�9�,�4k�������]Q�׀��Y ��mxq﷙�C0ۼ_���BLq�𼋠�ړlR��e���`�)1)>!V� Io�]�\_/�7.��������T�5rݠ��4�Yڟ@Xy��Q�`�+8ڕw1i3������������p �`���]Z��%Q�sh"�@d��<���fڳ@��dyӷv�cd:
�G&bn�w�x��n���W�A'�V�v��5mX�D�-G�f��JGUʧ��	�m��בּ������*'���&FG��"T;��U<���Ef��N�O�e�*ϭ�"��"�&��[��]}_��4,�G-�)����Qm�����>��R�4�I4O�oU<&I��1���@�U-��3P<m���������7"��Gd���>���H`�#� O������b`/H���Y�]5����ø�)�6b�#ۍrV��$�3JuO�p�ڧ����_�O'�X�k��_4��E\F% �D*�U�5�w���`�N������;��1�XO��nT#�}Sq��{�3��[�8��������ȋ�*�^o�[�mjбWb4.��}��`�H׋L�v�@���t���/2��&>v��( b֯��}�	�M{*{��y�w|~��~���x,�Q�˲����r�_ZP�J=��H���Bh�Qq(�>>���A�xI��c>CS}t��>Y6�!���ɂ����y3���]���j�ٻo�D�S�g���Meo�<`���SL�$'�%����x]���ظ��F��2��ʄ�������Mw"�@χ�j��1o�q�a���݆�V���ߔR���*��g�$��`N��Xo࡙4�X�Z�'�<z���'�K�'����	��Oj���y�N�]���T�.�\�N�)xM
�0h^��y2����@N4z�؉���7���b�0V�6=���u/ˎ3�� n�N���f��-'����Z��O[M��#Y x�����9�V|j9M�^�)�F�Jz�*����K��P�B����Mr��Cu�0V)U<ʨ��˦~�QjkȦ��P�������||繞L[��2�
�hj��3�B��q�(=rRg���
�,9F���D:����2-AeS�����/8 �A�b�/}-ryB�*����*_���m��N����m`'�[~���G����<Ѷ8x��Dm�'�[��� �n��2b���*�0�����fdL�$�ɓ���X�	R<wM�����y�HN܈Ҿ�n�����av*����{L\F�A5]rQ5�ŋSi͝�� ��3loYC<ʡ�^�1��S�O��w�>�*c ��,3ߔ�5�U� ՙ�A5=n5T
�k���Fֵ,��l�	�C�ā��Î2�J
g�D�8�!$�� ��Jr���I�g캄ș����Ma�b�w�C���Mݼbz:m�"�L��MOf3��~5�'�D���b6ձ�3�;���q�=S��ᙹ͉����s�ͩ�{� ϫ��&��i��H�S��hd_�L�F��v�5��64���'.=6;7{V���=���"������Ʃ	� 	-D���|����R�G�R͞��'��4�z<oE��F�Oj[��u�v�&/��$�HH���^�*ΰ4F���~��ںUgB�ڏ��n�g�!eS?6�b�`�d�ݖ[��n�,���W�{���	I���0���*��.pb���cI:�:�x��rc-����W!)Fc�BN7�q��8JΑk#b+x�$��/�R���	�ldtNyU"���(^|4�U�h��iʵ�=:�$�Ky��o��I �o-�V�V7��s�Y{�����f�<k��vWf9�[�d�LH���v�lט"M��6q���Ǡ��@T��OslO"����c5XC���96Z�0�ە��5��'��VȈ�C�"�l<V�w�����j��(�;�t����8�	�����2����r��a��>[�?+і��T���?�L�7C&kK�ʷ�l�*v�$���ݭ��j'z��\D�ƃ��J�c�Q����&n�9$���ړ+6�J��y��9S��RWb�����6 C[+�$u%XӜ��.�I�bl<2ᚆ|�Qo�]����l�f����8��͎|Kɲ��cȄ�%%�~�xj5BJ���C7��t������=�\21�����g��Y�QKn�����)�u�A	��[��-XFYտG��[��U7����1s�z�A��o���f�7�4�����j
~�����W������w��Ĕ���:����Й�O���>��~�?B�w����"6�����<Z?�[�*OW��>Ǿ�[�������o����B�$9��F� � "ɥ��d�J���]Z���� �Q�K9P��p�]�������?�`^�{�;��'����($�<D���J����h�`70��� �*����O����SPN7�/�C{���2�Hـ�����|O��쀰�L�IZr�R�|�-�E��=Dc;�*����p�E�o+gG|�A���=9b������$j{a�o��,i���^$��děS�a�5۴��~��UH��b�`D�t�DR8��m�(�s�N�5*o4�Zs���7V�"�5R�%��
Z��g�����l��Y�	���Rxp\�o����6��e���;�B}�R2���t��M]�V�N�M��r&�;n�\+?:��]�4����7Zg%泧7��0Ezg�6�rvk�}@������py�*��)m��f-�E�N6Ă�U�I3�Ο wWH��H=Q�*{�OG�u%������9F	a��izW��EѲ!�d����PƧ�Kz� ܆��w�I9S-}�8��ms@��ۄ*�y�6D��QI/�(��a�`?�*�����֊#_K���w�}�&��~�Y ���![Q�R��&q~i�k�㲌aKL�Q���v=*u�/7s-t����s|XB�:�lOgǄ�Ң���%��(��a������E�����>���Ԍ���(g:pG�{ҚD��
�r�>�oD�(	/��/n�4Aſ�G�0���肪V�(���q4v�M�ߝ�ۃ���m^ ٧�\��ϱJ����'��������І0���� ���PVt�U�Ԏ��Vl�`�iX���g.�,F)k�c�T�KI4~(��A�ѽ���JJOŮ-����<$�<�Y�j�2A�t!�`"GV��u�F&��J-�j�~߽�b4��ǉ�#��V֣^ſ���0��y�r_65P�K\��Ul�!�?1��3k��X�>��o"j��y�&��,����� �/�;,����%���~�)Qm7� �%��0��dU#�w�A�������?c����=_��@�_��a��kM� ^ ��GDV-J`�6Q���cK�·��s���a�MU�{��U �K����������A�F�n�3���8},:�2��]׍+ �")��M��˙�,�}��:��A ����:�_�'4����d��6R�H��C'�62q�"�k`��&��5��a��%�]��{�=�]u�
�v$��늢����;�B�
B��>-�������|�@Q����fO�H��y�r�N4�c4��x�G��9�${.f�#���`Y��;�����X�%Q�I"�"��%�\k��i%�Ը���'ȰO��y+���})��(�4��k*%@)Ls"�d:��������s�*4��>��A���P��\�q�wƽQ�"����B�� qD�"?�j5����J��KGUK1?��K���c3�#b��O{=u��N�\s�����{�_�uS�͵o)��.����z�D,����(�^'��`&H���Ǆ+R=M�z^�:�������||��e�Z��-�iؑ&�$�8��m[�Nmpf�Jc�,�Ҡ4�T���>qU-�"�CdO�ݕ2���^n��
t%T��B��F����W��%�꺃+=�A6�Qa��:���k9T��a���0a���*�7ysVoΨ�o��9��^)�S@}�x�]�*+�Au��ޯ7RI�����[��TM�+�M�^�m���� �3�T�N�Nj�#Ne���1/�6N���#�G!�T����S��t����_�
����f5�����Gj�G�
%��K�e N��y�z< �z���4����9?k����BlA����c�"��1�u�0H����p1k����������˥��!��\_�O�!��Kgj$=�[�+1����8�(6�Ƥ��Tq��L���Uҥ���uVu2�!�2��{a���lt0�²a;V,��ۨ��e'��Z8F��P�̗2T:�����zi���F�sY��JSq0��X`�����8=�Z�_à,7�ON���u-߾��fѠ-y�p*���X��3Ipx�R������n	{�Z�X��h�>�yigf톌ߠ5�� ~o����hV+���y�*g�8G���7]�/R�Ic�N(Ch�