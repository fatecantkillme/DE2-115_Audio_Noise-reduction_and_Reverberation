��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf��4Oᐢ��\����Ⱥ�UҚY]u��'%E���i�_s�v�؜�.A5�w]��o�8K��V\s��(cf�D#CA�h���^����ډwS�����o#���V�Ћ$�1 �2Yz��7t�K�������� [�+��%qm�0��C����S1 ���.��sKzp6���F�L���,e���IB\�k�,��v�Ŕ&���  �{ ����l�Q�!��� ��mU�&���N�X)�?�~ՒJ|�jM6�V�Z~ӾQ��
[_&;Ham�!}�x��p8T����Ҹ�j�����_�r��bԼ2H����@��q��+�WTA4`�����|j����6�b�}]�ea9>C���*sޝ
�N���*1��?����[�ρ.yF@!�*�� ���mφ�Y��:����"(UԚl@-U�z�v�±Kq.tȘO�q�/5N2)XB��3������-W�U���'C�~���A}�N�l�MBk������(��XpZ�;�C�ڔ�R�n�q�/)ida^-;�EU�#���q�F��f�U+�1�B۟,ʇ��֏����/�3i@�j>+2�&"�\�"�Հe�VX�3)Z�M�k�m�]1y�0��Z�	��M0�	H��兠���ue��Q�l�zC]�z_����	���{�%'�m��$cK�.�^E\/�k�eu6Ѹk4B�"#aȑ"AE1n�.Y�P���������p�b�þ-�������fݦ�F�@řD�=E��;���;t���\��̷�rl�D�/�E�G����@MA`[���vOv��A�B���c�{p�,�o}ȭ^t��u�t��i�&���޴U|���6�7՜9UF�D�+��1\�7;�F�@����֯y��D#��j��SgM���I �G�����MTb��>`���> {�\�z%��c�T����Ls�֯�������L��t�Y<2!tX1�����Da5*~d�/I�#0���Bg�=]A��������Cй*�P�S��I��!��$e׆���ā�ʳ����@R���׉>JP����K�fs�%>��T��Tg5Wk}}�%1	_�����uX�Iܵ�q�B�/��;���5��vA-���${�R<J������ǌ2�t҃��e\0��*�"w��uʘ�,�ahj���SuZ�����`.�.X�ר��#鎘] 	��=�<����խ��<��ɝbr�x��T)��$��灑�,ߋ�6�B��c�#OC]]3��4A�N���V�*]�b���.�c���`�3�3Q���
ްߣ��R��}:M]3�-��6�ݜ�0�
C��\K��v�،7QP���/�Y�^�ģ׀�.��~Ż����1��ww��XY)e�$�7�hQ�0��t��Qϛ���2�72��3��h�M4t��'v��nz<;8��L�������O��������P#-$e�=I)! �6��lՙ�.ٺ:��7nr8�Y�>D?b�]�jXW�� ~$�xk�";U�b,B��<�j%@Z,܎��!ʢD~di�N�-����aD%���Jm������te�0K(�����rHz�֩w	œ0�=�Y�}t� !E��$�.[C�Fϟ�0��J��_p����V��ݏ��`ݘ�K�`��=Os�!@�91y:��ư+ ]�#s�4lc2Dhd��s�UC8s�m|q���_s��@���ݷ�BC��v^��`�4G�2o���J���*}ƿ첤K�j얨F��x�r_�aMq�Z��HM�Pڑ	�'6j���F�nϑ�eI`�3S]"6�Ta�c����\�z�a^�qh [AY�;F�hm�KP��q�M�$Q|վ<ޮ��J�O2Ho`��=���C��Ɩ��.�@���"π�U�1�C.#	��fm�|rY����f�] ��£z*�SI.u��
�Y$�}��)`R�j�B�ЀBZ�`�O[�3�M?y�!�����Jq�t��}M&��~�C;�J�#��U��^�'r�8y���7���&��wĜw���r(�u@tޟp� �n�!��Z�(|�[�<�Q��N<Q6�3)��q	1����c�{lD�-7=q����1CJpP���n�~O��УctVc�m����1�I��~��܋씐L*�&{E�s�Ed�r�.�Z��R#O=q~ιY�1:�^9�󸌓ۣ�ux���۫����e��=RT�ij��^T�1���[�M��c/���2�ۧ��D-'Y4�c��vh��Iv�Ʀ��|��|�e`@�.bo���(�`O�\�Mہ��PM�G�`�	)b�$⚹���Z��T�r��'�����rKɞ}�b#�d�q���:_����M��������Fqqu݁l$� ��T�.+��-�̍`g]_��7K�b��}5T91	�jWp�ܠ���u��M&yݠ��4��)�?�����.��?��]!���F��D�j��EUG�N(Nj--��9�V��#��ܧT����������y_5O��#!�w"�:���K=��͘�U�Sp/s`�B��0���.�'�\
D�W�IkN��D�Yk�	V��F,zU���!�4)�� �L�ܛX���h�ɸ5kI��c��7e>��l	��[�;��[���X�U�	ᛐ��~���Γe��Z�՞XdV�Fa��=�Mǅ�o9�-�jU࡫�b��>;���H�S���_�2��k#�;��@!�Z�@�)�R(�@�4��=���%ί��t5y6-nAr~�b~��x��Y9�a	�*~Wcϟ�[A��jun~r-M��r�>��r�MF�n���d�B9PFh'*�n�	��(���'�^�A�V��F�����_�g��~�S]�}�5\Uk�>.����KX��FD{�nD�\�~%.��C{����'�:/iV���9��#ӆs5��Α_s:A��/�P�V*�یM�S����`�k����)5-*}6�"�ι��.��D	��|(I"8�S%�^SK^/S�'�j�����n�.�OQb�E�i}3�n��-���i(1F>Kb����ϧ8 *e�ԝW�!·�E.�ŉJ�:�	N����-���]z�Z��*aD��(䋖��t2�e������$��1�iH�f��[�yqM'�6K�겹��;8h}u����,@&ޫtm����XQ��j���i�ط\�f���5�,&.aKoU�՟���a���f�͒`B���[ � ���1��3u{��8<,��� #�R�k�Uȭ���g�Ѹk��k�F<��3����&ay������إ>�_*��D^���R9�Z�$�`B�H�Ӌ��	'p��-���Ô��C����NX�OW�>�ÑT�����<fI-�X��I1a�8V�ҥ.v��� }�7O`n�B�d|h����Kk_G/^RT*ɾ#���틗��װ�n��x=��0v�-IuW�������;>�6
��-�~����ǏCGU�\�#�;y-����A��:L�>]Dq��ÆΆ�Q���������ך"g�ak@{Gs(��X�+O5n��B}�x��Rx!L����p��F���ݩ����6�N����.�J�&�8�G	ж�w^�i��@�j�����Z3\C� ����b�]�7)��`�H*^�W��0uvo���α�ү�yGi���V��ôD.��ZL>�t>w��c��Q4v�H6�!�!�%P;xٴͶu�ס�qGm}�n	r(}�v��u��n܊�z�O/I���ﾊ���خ��n�@p�|��5Ք���!Ĺڇ0A+�Զ�y&�D�ޟ`�U�!�}H�Н0f�z;O�>VPM���Q|�l>S7;�yO:�ة!:`.��\7f'3��(X���;� 3sa���0X	�q���l���H:���Y���s��ON�(:	�]�6e.��+�V-[���	][ �_�B�Ũ��t#	�1ph;W�Yzm�\�Ӊ��EMe�ް8����G-M|Ux��W����of��J1A7�3�IV��qXve�ʺT�0��t~o�����z��;;�$��=2��"�?U�cA*�7s�
CT���)2�~?2�
�)��@jU���9�I�A~|�Oh�c����V[I�����M��Ʒ�7���Bm�O��"e�f�F�{o���s�Q6Ύ�H�w�%�i�)�b��?��l{}���e��R�I'1���J`�6(�Z�TGְDǂX�!�g~`�O����c�Z�3�e�����!�^Q���D���JzA�I�JOSM_�o
v�;Z^M����"zrY<:KI�g�C�j%d�M��?a,��B*��V�wӑ�X�ty�	�)4�Cd��D��@�����bvcM�q2k�Ժ5Ro�s�1�hqF���x�YGxQ*����$�
�~X��Vz�$E�G��	����w�\x��Tz�	j��49I����&���Ӝ��������v�v�X��}��
d�cQ�>��ޤw/M���P����E���wW�� ��nsg_�z��g�}�� 楛e�iH��3�n����g�J{1Z0q����G���������;(x�YpV�x�!z0xZ�е~��l��1���65�������&鳈=�D���S3��(�� @��HCkr��
��A�!WwU��(��:@��~Aa��iݰ�ڵz�"3�
 ʷl{�&i��Ѫx�����u@E�1R�m�;z�4�'�X}��D��N[��m*�N!$�<ň��g&�6��z��V-E�CH�� ^v����m���lbA��}�7[��ǯgru���>�b��q9�D��r,�V��n�F��ɏ+&��������wD�Ǡ��E���0�
.�����,s�g�@������	��*v��$;�e��XG0]
��ǆ-�a��-e��q����<UEh�V|��kؙ�0]j�Tt� ����)��N�L���;ߢ~|D��EYO���&{�NY���1?�k(�|J=���N{4t(��;6#E��.\X��E}IzHH*���B����9h��}�pR�ـȯnΤ�jk����GZl�	�f������v�S/��<��5�M
��\п.�[�na�=�� s�'����:��iF�c�q��B���sF�u�h|O�����5D2���U�}�]���dJ�q���г���5pٞ�n�X�+Ϋ �Wq�l�Qs�T�y_�d@-#qj�Gd��Yr�|p=×Ƀŉ#��qg���@��X�8���F)Y��v�b	xtL�������k�ւ�d�g���������L��4��lm��t����W>1����$�i&,�����N���E"d�-�? �]��]MB��*ogG�ʓ��:��>G� {� p6�o8='E?�\XFWl�1�Fm�=�����H��[�����d�cD�#���i�`�5<@��-<Qa�ի�0	k%�wK8��Vy}R'��1KHP|��0o�0kY!���hy�J�����M��	b�"�oU��@�F�]۳ʽ�J����V|v��b�	��
�"�e��P}�D��n ��f^V����wr���+Cz�.gO��V�,r���Kyۺ���dPxnc��
�D"p��	���d�YK��� م!�5WS��0r3t{���Y8���f	�~11.���fa�%M�d�P�BU1��|�1��)�K�z	�� ���!p�j�`��x��@�s�P���M�u���P$�/���jRk
�p��r�2Ҫ�a}�>Z��	ܜ��Qf�*ѩl�"?O��{?>ȏߓC�_D����;�ƈ����%.+�<�g��f�^f1]��oՐ6$��An���[����ɚ^ FS*V��O��^���t�#p�B8Բv�h`ͱ�{w��ӓ&�o.� ����A/n����4E����Iy��Å
5��#���l3�9��B3wz��kX� �Q��7�w��?�B��qp�}���e��T�ƹ=�)m)����EP��Х ���\�k�Sb1dP���׳�#3�`GU����}�0��$���(���F5K���r��a`B�=[��?V;$�U�+!:O}��j	�3٪�~`�\�2
��ur�2!`[_\�1���iՌ�kH��T�&)Ү�ߋ�b��i�{���vP�@�XQ3��ފ�գf���y"J��r��q{�d��u^g&�K��+�H���N?%��8�G�Q�t���Lg��塢T��)H P��V�g3�`gQ.<"��t��@^�8�������x��χ��8��>5������j	����B��M�U{,w��,�PzL���J�:���I��;p�8���Rᦒo]�q�~���0�ju����vZE84�O�g��k���z�'�B�"Fḯ�����cy�0�*�n0���@�/�7E��Z���l� +���cm��u#i�ˡ�3z���̖��;Kx�1�w�Ƨ~�PT~��[U�l�}��7~EA�u������Bd9�,�˶�Ɛ��������!�h����T;���+�L �}��,�*@����E�?H�٘'��\U��P���iUt��2�0�+4c�P��J ��{�u9�oy���;|A�&Y����|����r&�S�N�,0������\�|�����b녺�fRZ�J4(��?�5ه0��+�͹Ᾰ�*�]���E}7V88gF�!!.����Z[�.o��|+r����Տ`q(��j6�����P8I�HJ��쟱))���$uzs$��}�)�x0�M�LM	�� ��7�e�rQ:j��Ctp<��`�z��P�r,x��ǝ�l@�9�/cW�gą^g�UVJ���� cI����2�+Zxl�R|�J�7o�vk`� #վ��m�>F�p�AS5i[��Q8&8��V-��>s�Y��}�x��8�+OI��}s��pfk�l�gbT>��̱�{�k�fHzݡ�g6C��~&�9u�|*� {_��b���Hxr��2,0�`W��}M�e�O��=�?B�^+�-�G�av�#�j�������,�}q��Xږ�̤t�ΘA�FD�vjc��+q���oL�����ֿ�n@+���0��t��MY�H�'-w�Ҧy	�yA[� ��i��ZF؃��h͸ZL���������anm��&��N6ܾ_t�O�KB�^��fߨ� 	$jǧ?�w�|U?��P�����)�4w�%�80aHʪ�r�D?��w�%aS]XW?m#��C"@[`��c$����/�i�!�S"r�2� ���4��5<���XJ�cBT��݄=��n��r�
�{@H���c�v?S$�@��;�O\�,]k��/ڐ����tE����˶��+�۰���뙢L��z�7 C��W����ĩh)���!����u)�嚰6�V���(W�(Wz�ת�������D�추��d��u(��m��D��9�����xS�:Sڂ/���pŕ��Ï��\���u���.���0�l������]��^��xw��@�
�C����	�oD!I�,͜F���~%�ao�B�DpR*�e9��Sӓ�|�۪*g��?���C@5��&ǈ�р�|�Y!���k�/s`��Ϣ�1���e_h<��u�pK��6��{e��i;�.�.ۈ#;	�cd�c� ��i �����Q}�~�WѬ�Њ��
3��zǧpgo!"/�!�����0�/� �ӻ$�%%t�S���B�4;-3��mU�	��������9�;��p�)��	�����#��q����a�I�kN������Zl�e�b;n���gn���K��U���Y�� x؉��r����E�iEhX{�	f������F>��[ۺB���*��8c�����Ͷ��G#�4�ꕃ�Sg+@�!��7��ɚL�҇Z�UzdkV�Ka��.g�U�rC�6j��m>��n��
�ye���� i ��u�'3��hU�_���Nm��]J��x������Vբ�Sb� ���{-����u�w����/2���aƗFڡ��2aCi���@a��j�B���!q�?�k����`�`V��lƶ/�g���+5���P�y�<�2 @���w(��1��|��-��&ؚO��Os�W5r�u�ǭ6�V9�F�r���v| n�jC�?�� ^�NI7d�FZ����=�M�fX��	L�%I���'��c�w�)�x}Ƚ\�3��8!�������ZB+���Q �w%zg�924���U+�c�~��z:_��!��,2�Җ���f�я�ꖛ��E)�m\�tu*�2ZN�k��������2�oX�=�a��Q�Z��B~�6�m �I�#�� x������~]1�*"�]�6nD�m�ĕ��F� %J��t���n�P� ѹ�_շ������Mh�1��c�P�"Msߡͨ���"ğ�|�Ui��5�(K#aʬ/��0�
���G���L�f�BQ$qw��aBÿ����&��>X"�UT,aD�@O͝:���d^�i��́����1+!*�pn<��B*����R�n�{�����^0,4(8�d�"mb�#��,\�r�<�O~�R8e���I���>~鐒��~�wP��S`�`�y���n�<�=�S�P�*H����/����hC�M�sFa������;U�oQ�2�tVr�<�e/�h!5T\�Aw��:�iu$��S��Vt�#���-��=�@V���V��l�aFS��5ߎK��$~F˛U�d�r�
��_>b��L�Y'��v^$X��ԑ��������Ű(��8I��Z�,:¹�ϑ��>�6�3�p�LA�?��9a힟�u	l�
��0B$39 pQ]�R���+����agm����S���h��t-�ʿ�Q�Rv�װ/a|��wV�+��=�5/��@��?�� �a�Gx������U����Ӆh�I�UD�M�${����ʩ�~��|aJۻ�C��s�,�^�� c��[L�l����y�ru1S��$� +��SBa�2����,k~��rƤ+,�L�Y�	����H��:L��b9���r�G�<�ڀ�{w%��B�v��? ����&��]��{.|%���(6��oePM�چ��r1W���d�aH�Y�EΗ��sq��Q1���C��)�hZ@��"�'���XA|���3&�����إ/�׫4�-M~�cZ���ɹ�g��MK7A\{|��r6Z�6<*`��HMϚ�,_�z�\�$�);7]CE��t�ה�w�y5��ʲ������i�;2�����@�WS��ɮ�?� 3��䢧��N����J���V�Ȇ�A
�y��*�z�s*���p��,8.?�D����y���F{�Ç��� PLU���W�� �������Gw�@`�=���4�������!�=���eR������"�]7*=���1�fڔ�eŴ�Qvv��6tQ�ȵ*ŭ���Q��0�Q���(�#4ςm�M6�WV�1Vk����h���yg/��Y�l_�d�&���=JB�SIG���t_x*A�z��1!c	_m�ӓ�si�Xr��f�c4�f���lCw{g{����8]V|��=~�t~"��碳5���<��/d����7<G�*-3Jb�*z�&g��:��P���Z�'�N�J_�K�ϗ�P�j�i���,p��Q�j��㑈X7��aW�敝Fj�eF��ƬR]��j@���5m��8����dK�B�C5��c�9nf[�HO�~~B��	���6���+G��?�������KG5{��n�B3x��\��?g�K7�\K�n�=�'����9:93����2q��V�'���]�Ng��H���gK�_@g	<s*Q���C�Z�h ��gi���	��N�^1e(*��0���Sn���0� x�F�����e#�ӓ���v���y�
fFǊ0l���.�ˀ܆ossk~��'Pc�q����;�z����Z�W�4u�6W9��n6���Xx8�2���
y+���u�dY|�,�
�h� ��'�����F�fQ
]q_b����5��ps���!C>����<���1��d)າ��!s4�`��i]�B�W� ��H��e)�jvu����.F��"��z�32����ɕ���~��,��񤐿�՘kB�I��(\�f��j������E�����Cg�U�vr�: U9<X΂u�<�C�A�u�V��qx)�	
WG�d���{��Uܷ�D)j�_�^��O���"6�I�p:�I(j�)8\��fɈz�ƃ�gB��`�����=T���b�&�7pUwmU����݅��U����:K��\!3������a(����K�P؍p.4�����\�m�ը�����F�"鷿�w�H�3�����;vM���w��Z/ �x}���soo<�(�џ�\Xh�)���lI�"�'M�R����[
N}0�Ϣ�����~��<3��h���'X�ޗ��	0���1M_j��"i��C��Iy�dH_W[�sO7��
��Sq�m��.�����M����G������-��,����ǀ�4W�.���ɺM���(�i�Y%>�H�L��{�8�o ֳQ�Ў�A>���x.��3c(��d)P�WS�D4�l�F���6��V*�c�>�ʨ^*s$"���{ 贊��B��F�~�qg3�i��#�!�3|Ɛ��_"�y��Sld�5c��䋂����H(�<��vF�7��6�}�z�}h�:3�6�ɛy��Y#��I9��/sI��]�c�1CkփpY�e=++j_�蝩j/+���O�ٿU��ЀWA�_�T3���UOL������Q���M2���[�7vc1�t
�_,��2f��b#UxU�F��j��r=�>#���ױ^A�_���a�B��nYv��M�-�bw�(���j�s��-������c�E�����~���WR5ܜ�80�2Y�ނ8�ܔ�B�Y��@{	�~��B�wD�c��ܔm��8��x�i�=A�����c<��W���|��Ԭ�#o�b��|'1˸��T� ���,��ƭho�\�^���ܰ-��V�♦f���ΖRף���W�Q��_��d� aG�(I�06��S7?g�8����u:� o�1ܲ��R)?ZHeߔ�8����bE�6�/�G����I�N��g�(��s\�q�ߐ�_���*IєN��W�u�[�c�z �j۶S��+%��J�WC����4��I����D%�V�Ĩ��S�Q�����6C�BVM��]���u��b�����I�H�O�U<�bY�)�z���G%���?L�Ֆ*q�3�����P)��?�$~�n���FP�q��NX�1Zh�ORDe�[L8$ �`ϒ�0~C������K�H�s���B�|$K��N1�90;�:���̕U8�b��S�Us%ʲ�;��p��6C4�1B�ڋ���:�{?���,:W�6%�5:�n�������p󸿱�u�5˽$Mb��˒��z��Pɂ��U-/ L[ �-N9�UaJ�����~��ǫ�r���Z���nR�P��96X����/�|�M��(΅;g�s�uo~�p��� [��b��s����GzJp���aSS���y���2�T�㾦���hK*�kK\T�����O��h�^!&�1�����r��q����rj��곥���� 7f��V���%�*��,��^&����Nn04_�wJnưꟅ&[\L��-���iS��}�Sov�aK*(uK���(��#
��gخ����j�JI������\�Z/�<G����o�P`�[�m/�l[����2����_	�%�-$ŴHU���33���S{��EGF���֊���]�ٶ�0��S
��p�ބ��5��s�ꦣ�#��M��S';�\�[޷�`a��K�%h�E�5��_ *ʳ�"T`����˳��{�=De��f���yKԎ���Xq5Y����[�!-��?&	z_���(�6�6��a��@὆�������S��E���WCl��{�:���.������ �|�{Zl<��.
R��Y���6���y�����i��H� �AV����Ρ����z��2_ZwM�η����+�^��4�آ�<���E=��uʦ��@3iP�	�V���P<U�A�}l�N�r:9h�ֳ�y����?'"�؉����_z!�5/�&GvK��D& �%�:���W) ɘ<+�y9``�6��2k!���9MTk�F[�~^�&+�ۜjyM?ˮ�����^�$��{�:�,�"� t_����eM�Œ@Q���E�<<�<1_$u;���՚�p���h��r���,-�W���k�>���A�^����4%DQ��r��g�X���dҐQ�̦si�e�)PV�F�\G�0�y'9p\|>�WDi5U�$���R�ïl��b��,�?��΋w�0�?�-�4#;���P�3�5f�h�)���2���xZPi����,��[n�v7��9�|HG3��XF^ۜ�CO��M#�$��&mj>�y}�[�9*��e?=��G����gT\ߋ��?�[o��ᘣ�c�2�뫠I��{n�	6�9�2�l��c�#C�@y|7D|:/�^~	#jT���	��#�7�ҙ$��{P��Ɗ_���-�������oN�T��VF@Rc�F�o��mJb|�^��%B_��C����j��� =�����)+�S�(���k[�	�a�����2�`���~����iQ"�"�X��O�pGL7�< ��Ͱ�G�A�&���n�T�|���4�ma�Щ��ɾ]��ɮ��"a�XK��R'#=)��)\��Md�1��ؤ��	>�sI3]�[��]��?[����� ��Yϓ�*�J�J%���۷9���	'��e[T�.�4@���0���to~�%�TJ!+J�^�q\y4��"���l�@�	剐�1�r8vw�b#�-�;4i�߽�Qq��5+R������Z�b�<�=�0V>��Qg�(�)&����߃ 3F����~7�	��Uk��.B�vz�V�8�����|Y����}\w�<��(��<.9�"lRA�}f<��Y��*6��ͱ_Gw�c�ӧ��#e��'��W�� �o����
����B�̆��t�c.ƽTT|��	�r�[�Kƫ���C���S!F��)��qh����A�!��9�&)PE�%�n&��-e�Jɖ�}8���6�C�o*5/�$����(\���=��@��ŊUc�(���Ϧc ��؆����#��7U �	�(�z����)��'G�a碼h�-ο��\x�}��cQ��C�ʽ�G�{��ui8A�?f|L`�Ѧ���Z��y=Ó��.;e<���!�� M��WJ~ʢ��X{��M&>�9���X:���z� �8�-��m�/䦾�X=�O��o����;@M��CY��XSۥ�� ��2�z���L㕆׸Z~� pl�o���a���/�C���,B��v0�����7�,'[��H���4C#��Z�G����{�G���9�R)I�[��M���*�m��"����-b��hHe�D���,�����qֹtd�Q�<
"r�0��+�̀�K��S~ح����t
�yu�����T������GCT���m$*Z �*o�I�Z�@j�Ʈ]7�%+G1���\����K���;'?H=5���0�q�gͶ�[pT '��be����+��A����'S�=�������1�D��a���^�G�Oܿ�5Э[�@��0�I�_L��`�G�Xf��S��X}�8�}����6o��C�λD�4�v��D�f�r8��FƢU��i'���LT�	�i3!M������qcuX����E���4�bN�R��:���N��0۳���Xh����3���^O��Fm:��Z��7o(?��WF�|2F
2:����<��: 7�6��|?(���L<K2K���h�������#'�3�yŦ��*##&�w�жQK�<�� ����^��2r��Le�Y{/F�3H^����i׊mM�p�_������>&�98��2�@_���w�;WkC&���
@�	���p�R���x�"z��fa��:���ψ�8�IFҫ\�&u��Y�a���͂�x^-KD���ڸ���}\
�ʣcc)u�Ў0賸$:�d?)�S� ��r�H<U�x�H�!��A���*6��]Ap2�M�z@��*ɞ��������_@x�ؒc1`3y�e�����s��k��OQ�`Ы���]�9[�=F�,X1�u3nJDߜ���Wn�r�(����==4�CN*Zq��������OcA��A��][���%&`Zf�w/`UƟ���7���BM?�����v�Q�x��%�T��w�sg/˓�E�<d�1V%�}�i'�~D~��{�eT:ߵ��FM�ˑ���U(},�3e\�@C�-��7�U��� �{`/�������9�>����c�`:D�w�9�pcMݜCD6
���Ɲ<��-��t�՘l�s�Y�ݍN��_�)�hI�#��L=����ya��<�*�m�b%�-l�Q��G��+"�Q���p��N�	h�?͖��q�;���Ir ���� �oWY���lv�S��J���
9�
���j�iTj�2��7t������gj��X����i�J�.ԓ�:OMOw���M29�z�+F�jT	,�v�
}��yc.D�II�"-n7�3�O$��D�8�2��Ԙ�B��Ph$%�8w��Ћ��\��"���N�@IVش�8�h��4�F\{�Dب[K�-���U)�چ�����p�x���F-�"�����U��ć��Z�q�D�{d�9� �h#q�9�H2�a�������D`[��I��d��{7�I�
7B쮥���;����e� ÓI5h?l����+��f�ذ�C���	���m��GJ��6/���ǎb��z�|[f�{�F�Շa1�<����tj�:_Fd��+t�Q�3VZ��9���W��F�����O��q,Q($io��b���iRI�K�M������w�J_�[��ܚ}蹌q�e�X�:�1��t f������?� �I�>�(-��x�50 �=��@n��/�b_����˻��u���
�N��ܽ-|��c���'��*4�;!���>�5�����~=���i��>�;ж6�'�|꽕�g�9N��8�/U֙�Ǳ��f����&�o��y8I7�xC� t�z�!D�|��M�n��J��Y(A�Z7�A�ȖJ-�Ha�O���s��'�j�}��#+7�>1��8�K^+�o��X~�Ö��@���j�Ir��^Zr��v ��CVm¼��ą��ϵ&���T�TחUҥd+�b����f�/��0?�rA2߈��[���#��5�X�\,�߹�����z�]���E����;�yf���|k����f���1M26p�?��}[�1+���%#\ֵ ��X:PHݴ�XY�PP�w-i�7}��t"�83p$��|�>����C��x���^�Y	�b����T����Sr
s�bB���ί�SR�-����0�X�Y�9��a�ɮ#����,Z6����oG�l�����f-4=G].� 4Eq�e���r�@��4�>P�;���1�Rt&>���i�8隥
"��B���WY�%��ej<;lr�Mێ�S<{S����԰8�y^[ �v�M�����OG<Ō? ���S���O�D��9��z6;��&�u��M��uj�T�%��Ҳc����*A�HR��e~��홴�f��ҡ搜?�9��C�?�|��.T[�O������.�)���j/0y�}Jsp��d��=;��C쐤�!��8!���W���X��A}9�c��s�"7�4a�C*,d��Pi���`���r���_�:���|J����0ݎ�[ȹ���t�߷�� �I�/��R�Cȝ%>^bPXV���n�g��&��d�+4�ļ�����/�(��UӀ�'�όqŎ;����QTF��S���\������NRb��畭���ԅ��޾-����4u�&�J�E��?3��ih��S��c�~t,"��X�z��Hɫ��:�#���c���	� MP�☑��u�k ��1�u�ἧ��Lr̻��+�g�@����Z�'`�+��lp	k>��hb C���E(�ꀄ�o�KQ�QSW�rv6�7춵J��_���St����uN������ot#�,:��3F��a�ag(n�W��5D�%Z	<���VEO�	T(�#�}���/���v֜	)c�|�����@��~B��MèG=Y�C*x�Y��Ir1ӄ��_���.R���^�ؠ�|����X�xz%P�Q] }∸���մ��vx[����F��Q��e�l��ɖ�$��cD,���eE�Dcr�KL?`���y� kѪ�fdhT�$�+Y�R�%�(f�
�
�^w�e�K=ma�U�޵R+���K!&D
�T$��6c%篔8	��+te/�ܶ���$��^cO�Q�?�3�bhw����%^IP)1m�\�!��1��K����J����Į�	��t�b�abVk��`�$��G>�B���V���-��S������Y�Ս�g����O�q�ot����R>E?���@Y�40v��E�o�m�{),_�_s\rz�Gg��e�8��X�D�m(B�`����-��bJaTj w��f�ʐle���c��Cg��R9t҆]�L��$�%����: �\Y���7C,���n<1�����na$I�ͯ��1֦�UC��{�I�p�T�GJ%T�?�V�;JvC7�i�)���25��L����Ӥ��;F;�.��U�$��RwZ�(��T���QlQ����P��ʒ����E�:D&jr	��p��ifz
ɤ���Q�ZC���FRM�����oI;w�+�<�7Fǟ�?��<J'���J>l��9UX�7\N�����>�Q�>�	����᭮�b���B�5�H�m�r�;( c��S&�9kc�ѪsB�\`����I�