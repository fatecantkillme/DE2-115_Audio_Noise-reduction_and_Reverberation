��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�8k�)9�k���J�f ۘEN�R��>�Ug:�&�1�����E[�Dm逗fh�~IWwI�1uN𙝿v}5�[2�'������d憐+i���al���gmҩ�ͧ�>�p����^m���\��T�5�̧��w`9��]B[��J�]����5������?_����%���l��� �b|zu��P��N�1;D�8o�f>����>���j\�!�P'�Lt�n�M	ճy�]��͔C�9���h}����V�'\	�6`�8�0���N�U�/��������UOur�2 �G�x���\�wgm������*����<k��]}��آ:���)-���o+�@Sm�j	 �Ӻ�T�Q;-�㕦��{R���8�4��H�*ħ7\*�ؚ���ˢ��p�v���Ӎ���l[����u%�����U�5��,���"%N�$ӻ������~eh[F!!l~W�mb�)���3Ф:9���͓�r��l�b�B7�1k�;�L@�$�{l��+��ϊI��Q�8��.�[݁�<5@�O��<q�z˨a� a�
�G�?�,��}>��m��=��F�[
�9���T��}����x����E��HV�B�5c�sv4��Hl_�k�g�ȷ����01t*�Ct���K�9�u�:������7�>RNs��t£.$�׭��f?/`�u��p��V�<U(����H���7���f-�?�{�����B+M�t�5P���Y�\�0/�)�HF�S��#!���+���/49�U'�R>�v	[��F�z^N�Q�i�b��;�����Q���g�py��+���j�i���}	V�B��k��nn�ТJj��ՠ1D�)y[���󟰥�>Ӟ:fu����m�~:�h��B����ᦀ9����E��.BU3�5�W�ARJ��h]�B D��c���� �.�=�kp�`�+>DSʭ[J��f ���⓵&�(���iV��M�I���o�W6��7��zc]!'5�3O�,ы|��r\S'�|�]��Y��3�f�@�z���hO�UJe�jH��v��L���4�8w�B�쾯����O��^zې��ԩ��A���}ϫ�jC<JG�>&�o�r^1F��:�0�\�K+*g
��*�8z�[��ݳ���OO⮜_Y�u�G&���Dkz${�:���P�h��8�� W���t�Wpi7������o�o��M*�Y��7H�4�;�k4i�pU���Тs�}b!\[�an��}gDo_�����
��:7'�]<F��&6l�1��]��HO��D3���ӟX���@�P����L�s7q���Kyo3���Yǧ0���Y�$W\9���k����PFE#.Wc?
���o�ه�j='�j�����s4�1�t_�?V�wo�!�Ts�"G'w~��\��'�����h��������� ���d�x<�GZ�8�H�^h��-ò9e�s�݉s���3�(��u� �s�2���pp\��
/���6�#�ہ��=��X�ȐN{�f
M<6�X������a�څmD�p�:Q�m8Qʑ���QO�dXW���+��H�ф�.�����Z���݁國u���e�8���	O쇚���������n��v��g���[�������M��!V���	f�N��M�zO�#[]!�i -�l�lZ�Dt����\�C��� �<�n(��t߿� �[#�)4���0�}8��*��6+ږ���6NFL��m��Kc�\`¹,�F<6�yH|�f���±��5�c-?���F�A��ȅ�Oe	�yxh��� 1l��(�r�"��1��⛞�Z�Fwns5�<G� X/�fk�D�J'��:F0��`7�����F��[�m����GLگ�XTI�<�9�C�:�BZ>=KvS�ӝ��N��K5_Т�
��x-��Nk��r����#�� B\up�r��pl��!L�9@��cC��^P����<K=�.1�B�ʦl�Ӭ�����x�j>Mq����IvBAM�>������}bN���be�MR8�[�o��p�1�SS��Y�6\���`;��h�Ed>
��wt��>N!S�oYKV})���eL̩��%� 2?ʝ0�>�G~��b��w;���\h�>_ t�?Kf�������O0�z��nin��G�u�^k�P�ێ)0�~��v�d_W�L=�Wm[�����O���Y�U1Hdf�vv�Oemh�ZiO*[�tD����Cu�W����F�_���������PY$n�緝/㴏��_��0'r�[]���w����Y�a��;Z��>�4֦��\W~�=��w�k�$%m��$#hE��Qf����S�����l�����7WM {0xM�#�fZ�N���h�4�F�31!�}���"���q�͕ ��2&$Xr�d�aHdf��K7m+>2ȶE�#�uj�����Qk}9u�yH؃d�_�E�q\��i�p!�S�!W���!�)�K"Qԅ�h�y�t�9C�^b"��+�ks�[jLj�S�(��7�m4����`�+�Y���ɰv@�>N����E؄ّ���d��))�{���6�q|~�E��]�e�J�����`�D{A��X ����j¤��]��ʁ���A�T@`�=�rsv�|�#�}&��`=���wǌ�,�:N�\y��0��Y�������c3�O���Y��+��߳�\�f�֖D�G���Q	Ӕ��m�� U�v������o��u@b�3?<!Ne�z����P��	�ذ�K��t�R?���5b㲌q	2�9PA�K
0�����S�y��ٝm�O[1��X�Vk8
2�_�6!���RfcapϹz3�C/&,�V���5�]�(����u��G4<��))?%�6��+zJn�t2����A���+1�r�h�P�vF֍I-1~Γ�&1�e���.:�յG�pS�<D�ǧT����8��>�r�JЪ�&�?�S#��^�VJߗ$}i��1X-Q����~1������\���ױ�X�R�����/��4��!X��=�I6���
�H<#H� �K�P��'ˀ�Q�6K{���k���!c��j�	!_�J<MQ2�6Aܥ���a����*D�H������I*�.pV1GaSuE�a�# K=2�����m�Fb8�y�PZ���Y D�qe	O�����vW}�Y�E�z���c�?��`+oi@�K��2�H��CI���P���˾Q6J��6�Jy'Nb��Ƶ�������U�<�a��3�F|�1何�y�:����_�HLU�čl��-�G1�q"!��"�ss�qθA��+ ]/�dMṴ�\�R>�4�{;�BG���;�,�J��MxZo�-�b����}��f�Ͳ����/Sd\��P��V0
}K�����*~:���N%���ၣ��Q�Ҏ��%�vX.U�<+p��-M.�|���W���x�� v}�r�� L��e�ll�(�z�io�
kC�	ǁ���*�,�%hK���@���&�o�3�
h<��o�/����e���4�;MoF��K��d��Pb�K�%��JE��B���b�@����f��_�t�aN��㽟9, S>J&���Zd_��*���yZ����eI��n���4�֔���
�L�7���O�ae�˓�{�?��%U�ف ���z��ol���j�+�P`]���ea9GV�vk6�3���Rў���[Ỉ��z��ջ�)�3���gx�F-o��]�g��1$f_�����k�a���SY���F/�LkT�?��9Z��#��AQ�%*F	�B�Q�Sׁ�ǖ/�5[=�i���@��H�mm�ے��=�U��"�n�].0Ν.��s,�A�OQ�A�"�g��r#��#���U�s�� *	���A����|<���4PC*\�S��cWso�c E���SJ�I�%|ɗт�2V�N��nt���D�i܋����jb`DzH��lAP��#a���Z�'��B['�^6_��I��]O�JX]�
B��9����=\E��K�ㇵH��fd�7yo�[t�����u�")��YV��N�6��H����	�����c�EIQ�T�Fu��kא��`�+M��2D���]�:dc���{`(�CM-~1�=�ЮU}�B�E��vs�OL�w��(ૻ�I��O#�V�Z&"�Mh��۶P�M/\�۔��,����'��v�#�P�LVŨt*�_��;�Pg�Eh��A>�kս��<��0 ��B��ֈ0g4��R���ND�U3�-��V��Y��KVۘ;�ק;Xۇ��&�S|{���b��|�C�G��%����}v�Ia&HU@�E��U����DMEG��.& /_�1|�`�=kĜ��D]Sԛ�1�f�	.����4���f�oK��Qk4���\�}R����9��D�ݦO�|.��#���TK�p�e�u���lFb��_Hj����4�Wh���hF+N�۴"T��(0s>��}g���#�[;��y���j�f��`u��洑�I���9����xh͊?~�e!�-H(��z1QQC��Xګ�FF�yztuu�'�q��/E��잰�;��J��@G�U���o&# ����N��7;����[K�Կr�w`�dţ����Z)�c�y:9���A?����Y�	�j+�i=-4 �B܁w���9� �CI���L��H�"VB}I\��p���қ\!�W����}f�o���8i.�`�@}������Ô��:u2��®F��&�hڻ|�:nS%�\�Uy�9/�w��\�����w��G�� ��Jq$�K�2>M�0�mG0M�/�c_!�ֽ��&n��O���(�7�Nbeec嬧��af�E^�EA��Rh�2�i�ǃ���7��k�`����{���;�-�%��n��Y��^�3��kv�_h4x��q�A���9 �oC6�"b� o/jN�<��6�)gEA�0,e83�ڍ�� �>�X(
{�<��!@El�Hc�8�j]c��a,3��Nœ:��.�>G'��3���ۜ�����ϑم����HV�*5�s8�w�LIt��$�'TQ�H�c���+��a�F�j��j����d�Y�>� ��z>�5�S	�$��f�k��T��	{"��<�䛈�쥛XOTsʨk���s�A��Z(�wit��X���8��yQ�f/v��f���\�V/�R
�� 2�"��J�w[73��{{��p5��֒N`�/W�H�.N�R\qDE�I���e�����dԪ�a ލ�K�o�����/	Z�C9��Ɓ���f��ǃ8�	 ��n=�DA��O�!�:����Ug��*�4�kcƃ�Bb��C�F�N@�\�q�጗��Ƙ�(��}��x���i@5����ǵ��//
��1�ꫯ)�w?���TE��J�Vm]2���,�i΁	���u%Z#W9��w��B��,��q����>�+�] (��50٤A\hG*X��l�"�)�^|������I�/(�	/m0�QZ��a���ip�"��¼�떯6����n�`��t��Dn����a7�{���q��a&�r���y�Ґr�8@���2P�J(�����^����*����B�^F���ܟ������R>��9�/�ʒ������n�L��L��û�?�c�J&4��ω��&2�9O�� �*Tw�g޴7^��?�G�%�ohIL��;��}�H�����h�N���G$�(��n�w3�`�w�g�K��;P)Fw�&�� �&�0���v�Ewu%���3J!h�t�g���
O���5*�A:��)\9�
�3�~��r�E��V .�����VGN�Wea�����'��Zz;��mRMZg���8�g\����
��"`�Xq*��n*�.@�䋓N�p%�M��ش٪:�F��N_^�M�Mˏ�6�B4�C)c���	�?ȎJ�? =e�j���ɘ�ښ�GH��: ��?��Na� �N[=�G���ү/y���4G>9�r�˸o&���a�	:pq� ���de�����73j��n����Q�&�5��n79O���}T
/�Ɏ ����x����i���wL\��F\�x5ň����y�ݫ�2�%D��r��x%�Y|�G�/�%�����Ȳd!Fgk�N|���7+����b���E����s��b4�]�߿��J�����yc�R�;���.:��R���QLcq�0�K����7�)�A8Z�ߋ�1Crk'���Lؔk�d�`
�{ٕ13�`�3(
F�Ӆn~��5��=9]������8۽��3���?�`� ��1�W�Ȏ��C~���)G�V�̤z?O�`Le?��e�!5��C(V��(�	�e��X��a�-��zv���U7z�nhq�VSq����Y�E9v�H)�(9�4�G�sTmCv�1���� ���m:�	��(�(�0����vZ������L�k�By�Z˅����8W��vUSK����#�3��Cɇe�O0ǞEP)_r-�������c|�W�B_��Ly2W����d�i�T�MLu�8��U�A��R�2,��y�TNuv�ۜ�gJσ�3���N��y@-�G����?*bѵa�x�b�%��j۟�L��RWG�鯁�ݐ���D\�xF��S��C�������}:�I?Q����*�)RBd�Vx��vR�Yw�S0�yi��i��|H?2���+H��)b��@nS|�-��!)⟨�OG���|Rv�}��!��A�6��߭��P�.���y�(uc�G#���W(
ܺ縠�a�j���
�5
u�J+os���?�8�����ɵ�]�i�
 �/ d[2���H��|�A*1 �[���»�=uk1�>�� ��WxS������I�]�Ғ�$�^���>�<��xi�j�&���,Gs����-�H*�w�"`��f���?�u���l�Tc*����^6�D�3jd=w��@g�h%$͗⎾R	���>V����x��RI����&��E	i7qX�wG�jƃ����'t�d�ǐ�9yB�/S��"Z��wQ Iu�w���m�=(�N�~��,�i[��DjM@e�;.�Z���r�h6%���/	����L�e}��s /�n�c�r�(�0�qe��QH���ɦ�|��EJ�A�4+K; �t)�盳L�ZaB�\����;�6���×ȗ�-Ӏ���+�`&�Ca��O�Q��_�7�`k%%6�wΩ�)q˽��x�t��H���#̌��3>C�
�<~�g߸
6�a݄�7NN������\��2G
U���ew7n��H)X����tM���_?*�+���{<�����}s9�:�Ǻa�M�v�5a^�{��,5�̨e3S��kBЁ�j6M�ZR6ث�ڔ5�.�i.AolB��@�F��|�c�)�\���t���=��P�<���N 8!g���P���\T$)6;��o��1���5}� u*>��֯}(�SA/���b$.�>+�r��yX��$Ty{�~HW�:�.6�E�~�Mٺ3<�~Օ~/:��H#n|?~����6Q��.EG��,��xY�ʹ���������]&�%������G2�/!Aa2���;):Y^Rח:�V�I�-p��W.�T[uIp�+���Fe���a2?�Ḯ���vf��:�
��z���f�϶�|�ڕ 5�'\f��΢����B�(ů�r��q(<!��Q�w�;��F#]2F`�N��F�B�@ٰ�v\VS$Yy��/�������}>Y��q��3��!���(���n�L�e˞<��{Ln��,4��  �y�L�[�� yk���	���ȁ[����Sݸ �D��:<��$�������DU@�R�&�7��Ị���2E67� .�G�ں��H��%��n��T'D�Y�W��u�j�[H�����/�������*���i��/�K�k�wɴ����7�;?z3��S�%"�b�eB$SWG�s�i�3�:��=�|G5Hxs[�φ�ˉ�>�߇a��0eR��sv��6������?�8��n�'Ѐ�~	�H�X��:����P��-I��jT��d�
r�03|Y�V�0ԕ5	���bU9ɟ:r$�� ��R���M~i� ���a�a���2�F%t�Jor�q!��cюc���Y�JX����+�F�I�YM��h/�d.u�4nfK�X�GO���U��c�ց����wW�mr�g�Kz��jj�M��7�z�6��	�Cb��>��N쨡%{
����b�=w+��e@�Ɵ�0_�V��KW�'�����WtB�cq �ϡi�S��� ].]UV̻W���L6���,Sxo�+c�>�瀧�,�Zg��_J:h3��(d��thE�;�}O��$�g˨dv�Z&F��Z�;l%���O�V�ҰJ�Y���nw��h�d @�|����e�N����t��d ��9S
~���j�6l =�o�t��4'mhG�ςh_k�̳ga�>�MbO�D��P�a};N���>�����,��·�-��>�94r�����<��?;�;>�4W������u��4�ؕr|i&sRV���k��*�}B�NXt��,yeL��+�9z��e�-,��(�敍��d�prE��`�ǒ�5�}�05^�/��`����`��o^�6�i%�V�����_�v��E�%�N1㋷��*�8'�빐�,]�'�c_���.&u9�#�ټv�M�r9�Y	��q��X�n�e�����}Y�$��P�m:���/���5���<�#u4�}�̘�P�,�#���Ji�O�{d�������:���"*٬&M��&qY�Ȕ�������E���p#�����TJ�����%`.�����ߺ���z�$3�	�0���XUT�a�VZ��- 1?B		m̆h�m�$��S���+g��D����+O�&��B�"U�N|V[�����	W�h�'����ֶ�=�*v��i��x��~����~@��ƕ�׶t\�Rvi	(��Q��<�>DĒi����/G�H���*��
`�v�)6�YB�@QCA*�%���.�tUm���̍yaZ�r���@Դp����K��� �r�R&��(0��1L@LH��;mB�»\��KXC�	�"w8�w�6&y;B����dr�\�p'_4I���Qs\����4�A<錗GKŕB�zl�2E
_G%�!ܺh��]��:�jt�YADX�z���,���W��7]��W@C-�;31�Fg"ob�����	C��J���3���
�#؊R.��V���!�r��c���|��!�&L��d �k���@�O�fE]-�4n	�A��Dl�P�xZ/?M�u��<e]� �o�}��k�u��ҁ,#K�k�n�>5/Lh��0���{�&Z����I@0j��lE���׿X�!^��T�a:JUa���[���ݼV*u��H檡׬c!~$Eө9��yᓩ޷cF� a���6/Rxw��M/k��}�Hx`�?g&n��M�`�.9L���V8'�?�����|���X}e�>1��6\I2�n$��J	�D����s7=�1e3�]T��_�N�<HC����2�������ʋ�\�B�O��x	0�3k�3�3<�َ�.�0���C��0����;�Qxy�`MY�ˡ|�ۈҞz߅Ge>��\�q�@�X�� &۳K{��-BZ\�Y a�����j@���X�N��gC�]�����\��4��/��'�}��R<n��u����"�?����N���`y+���)�6#�D��#�ٺ���հ8�'``��s�xc��u�������Ɗ ��0a"������a
��\���&��������d�H~���S�2�B�k-��"�~��}���p8Fi��ٿ+������V|z�]=��ެ�Ĺ�� ���st�|W�]��SN�%�;	m�e ܫ�j艦��O�T'~�I����]�KH���g�G�A!�	�@+ �[��R��������nQvx�ʟss��|^��N-�gѣ!��:�@WL��t����X�]6:>vF��و��Zw���Z���U*�jq�'�i�.JL�A
�ٯ��MZ�g�d��0�_o�s�u;��tΦ�<H*����ڻߗL�(�޷��"�.Π1���*C?�t���"v��-�YR�=��\�.6o���w�m�{
�5}(������w�6%�o�xO
��_���2c������1�����暥�䜶��2Kf.�X��?y�8L%��<>�g%�c�+��H;ݿL�ء'[c`d=�s�n����Z�"F�����X�����۔��a^��^��O�R�X1���ZO|�����)�M�?��DE(����]9_���2��NYZ0��
�F�\�J�ݮ�H���T*H5�f�u���`(A�N�9H�Z��6��R��}6�7��*χ��������؀9J��+�װ����.T5 ��2���H�C��8�bȹ7�=��q�ݑ"y<s�Zq�P���W'�F��wh�)�bvf���~�=��@���=t7��Ȋ��K���m	I��b�|��G�[D�o��g�q�9�C�.s�|����H/,�{y�"��h�n�<�8��}i��Coĺ�$�3��Q�$\)���&����v��2���hzs^f���Q�FD3���Va:[I�,��'c̷�#���K�����A;���~��7g32�� FN��8O�O0Y��"�2~mߨ�Q!�y�3wq�V��a����Cx]~'SO�Nz��v$7p����s��M���]
�Q��Cə�=�;v��1�K8���A����7��:��|��F�64�YהUš%��~�V��cǒ{-�n����eU�ET�a����SC�ej�>Ə\��dr�-܌�	�\��E�;�VG��n�ø�$�[y�Jbe���2ķ�+���}�?�����JA�U���}f���[�sңR:�ows�U�N���� G�����lKO��W��/���6<($O���F@�W����+;�/�I�P�  ��������P�oe��w���"���$y�|r��h�04�P���7w�`��c*/De�:h:C+~�����"m��*�`.�(F�R�����! ;�'�"�]���6Ԯ��
��_�ٜe�3��ơ����>���I�Vˏ�媩��t���?��<��*Q���"�vh�����,O ɞ�$� ��U��G�,Z�m���bZ;Ƿ���������6�|*t��p���b����{�Xk�jį:�M"Mҵ��EH����#�<	1�쭲���=�[��~��˔�!Zm��Y�����"੏��\�����D�	Yyn�>�N���"�Xϯ��Ћ 
��G�;h-?��as<(�C��7R7atD�}Oj�>�cS��}�l]	
�D9�A_��;�CPx�r�r�?��g��+k�f��4T�A�t ͡H�(��/�)�L��WA���=�t��i3~"����>��`�pP� d�D��¹mt[�B�^�(\.��eI�|2�J�;�M�佟!�����":m�7���m~T	���Ό�F"R�������Jх�1�~����!V'���gB��J9��"���\��f�6�/n���Y��G$n���V�;:��@"o���~��A�ogF�Y'Vv&[�ܟnc��w���V�z��A��9��@��Q�o�L�F�M7�i��,a��w��54�ʝ�T������\
��`_��e��3	��V.��z�
�9Os��m���D
����P���Dp�9�D]��x�����qK�	��ގ�+9Zn2ˋ]�r��F{k��e<�G=}����e������	��B�j��C��Ns�%��e�B�����������n�Io��|��"Gn����x�ݚ!-\M�j�xM?`_UnH@��L%о�\�ǣH���Rr�<oy�����JP;k%�#���-�{����O��h�8��{���F�u�6/�6�=lĢ��-X@%Ӥ���t�?Jl�bt�+@��mqE��`���c���qu:^�{�d�&��7�).S,���LS��|���B�R��A�)cGe	�o����Y�Rm��y �Wؤ.�&�k��JB�zx9����G��S�����@I���g��m�D$QZ���ZT�pZQ[j �ν+�+5z�2ޞ��D�'2��� r��?"�wܜ�E��Ȏ�~�h!����x�^UC�`E6����������OE:TT�J<
�����Y��8{��D0t�1����e Z��@��(���fe8{�k���z����_:|+G7�Vk���D;�=�C3֐>�&����'B,\������i5�6?�z6MbO���,@ԭj|�k7l;DV/S�J�3���tȘ"E�6C����,����H2H�})���f,8ԥ���D�P`zve6\�����,�
n:�
��W�{�����Lbӵ��3l�_�A"�5��]<Ldr:�p���S�O�|c�+�vT���[*eQί�>�OϹ�pb;�+��%�q�A>��& p��_�d�؃�):s�U*�9�a�f\�����Km��������Ȩ�W��Y��.
�ԝ�D�J��Fb�i�+�5A��t�o�nR�Ey�_m�Q�w���0�)+��/?����a�
�D?�By�dD���0��HqS��8�+
,��W1Ao�	�P]��L�s�O���=r�S�扗ʊ9�&�}�H�D�烦[��#ɳk�ʙ,m!3�2��w p7�xB���<�Cx̀62P8�~������s�5X�-�ƱhT:@�A�E�yjJ,Y*�[	���l��- G;J���]�����fPĜ�����P��,ȸ���p2��.Ҏ�1���������y�/�K1Vw�^,�1
�P�Q���Ġ��Z���I��Rh?_ø�ց���0�-M�Zp-��w�ʊ��i2�[�����%�:oW�o�FU���g�J��-ݴ�h,�B9��c�Uy��=�o��S��6�?'�����%s2���W��k���5�	u���	K�d� g+����9��S<�/��8���Sï��U����#7����Up��^��ar��d>f��p�b:6f�A��/�h��mz#���o=K��!p�p`�!�ԗV��1d!y�F9n=2�M����IT�f@\��d�'$��݃>ڦ�< �n��gu�Vû��x��0�>�xFRd������7J���Dբ����A�\�!\$5�U�&&(:�5�唨�6��Y{\1R4`;<~vcV]j��;ל"d�&��[[-�b��܁�>�q�C {��p�1ct_��VS���F"�
�U$\�0,�:�Ô���c�l�g��K&�@V�g�����x�9�x�&��MN�Y�X�P68� ���Zg�AR��s�͖v�<R=w;�">-�K�;d�����Sxd�ٛ�VL84��Hm�}L�y�(��޺Ml��G�D�>��*$���7S�V�5��ސ+�	���԰��*�uI�t�n������.�a﨩� ����*It�Y��qܦ^���:"v�q����z�lw0����X�`�f�5N��.�^7L�	f�u>�P�,rc�<v/��O�w)�����%�?.+R�J���"���9��X�����gsƤ���iM���!V��f>��G��O����T,Jr�ٛ�[-����˺8:�k���k�7oR�3A��M.�&�i,�q_9,���C+��Uo�Y+�Nlk3�`���1����l�1�Z��q�8ӂ�����D��f��!�J�+%B%S5颐���@��z����(��ώt�����y=�b��ɉ�r�<9~B�63���X8^�п�>K��"8��fDc�n>ÇV��	b��Y���BТ�4�	��&����dc�g"�9�F�B�
����z4�Y�1~ߺ��A��ޞ�����a��c�d��بkybm]�����Ş�q2�mLdH�`\��uNA�!ai�l!m8���J t�s�A���p)RS�j��Ob��2;���'�(�>4D���������Ud3�w��n����5B�zt�e�<�~�y�(1��=�X��|,6�/�d{�TO�njQX�}�UZ�v��G:�{�����-�W@��"e�fS�Gـ����mt��C������"O���xg��z��p�p���l���@W�e��p�c4Y�	R��Av6+�2�ý�we;[=<� ��^�B��ٽ%���k8#��qwrtw19z�q�V�̩���v����R� /!1 �����S���!j�y�*.%T��>o@*�만��*9?D�Ԗ��Ԉ��B�+|[��4�	S/2�+���*���U''�n�,�db��o��(�|s�k����f�SotK��� ^K��Sj`�L8���.���V
X�5l#awM}���u���OD�B&�k�޶~���|�:�J�rN�,G�
kEq�s���ӭ)�9kff�k-"��r[�@��_ʰYj&�E��j���*3s�KHU%�Vv�����¾d6pG�0�]�Dg�k��;�`����ҹ��PR2!�a����}�r�g��OX�ٕx��u��\�=�p�N�<��Ŗ�R4KL�,JL$��[���U�2O=(�d��?����k�T��Q�EJ�N_����u��xbE[�[\0��y���Gƌm�n�)r�~:�������-w�|��9J�J��֍%�x�;���BD�ݠ�DU�m�̷V��I:���I�i=���&�r�"y2�צ��b���S�@�TrJ,���T��Gb^��p�f����������4���c�~�'���)n_/靛�QH���q%|p��8��5�	>�'�`�0na�oXh��j�3� �M���s������9�\2�����G�k	R�<,)��t�c�(F&d�[+��5�e)z��.���MZ
Au�Z�&��^� j�L�Wre
L�j����%���G.OOgZ[~_�(��2?`�1�\��J�J���D�������J3�v	ˁ�­��W���=	�
'�������[�x�_p�J4�-L��Nt�ė@���Y������@���.�y�8�$�N�:�6VJ8��iU��智@����1���9�,M�TĮR�L�Т�w�ZD�i�_��]}�>�j++�8�y
2�)dYS6�4����D���Y����� ������d������&�_����b,����(�j�j��з ����[���`)k�5k��S��'���N�%�9��,;Um������fYqn���x��o�i��&+j�䏯d�K���cc�����:)������ia����y���_�ɵ|4v�|�"Gb�I�UHzӥ�=j�L*J5v���P���v'�<ȵ�m�=�D�:#�h%xde��f��じ��S�qT��L�����k���`�ky�P��:Y�y��.\�И@:Kn�9T��Ā`���rU�t銘>�F?��ag�4o���3���	|�:]Z������5����y �[���=���w1�O�$�+;ծW� �pj*�1��r b��Oت�Ej~�k�C�po�W��AT�n]���MU�y%rՆ��f�y��_�b�����s���w�h��c��W�n���b�kO=�uo�hC����+���^������>�^�N�Sg�3#� eU����d�cY��Q���\-�1�fby�*��iL��3�)�%���p=�����B��4kц.�2�hV�Rg��3p$s�*l�M�[~Nv������6{z7�s����o�^���qI�Z�1;�8W:y4��������pmW�(��!��nz=���& l2ܨ�z^z)�'���K�'GF�H����@;~�K���>�Dfg���4U]�1�.����x3-a�aX⦸j���'�WgdO	��" ���%l�FB�*�J�R��z�r"������J���i5��	�D��3�O"Ό�����I@��i����֪N7�oG:�%��,u�!<�E�:x�E��)��,�ή��|�_�ɡ�=��w�> �M�#��i�\Bt��5��f�K
B�4MS\���5��B�tv�䝜0T,��V:u��t���� Ժv>�z�%���59�>���D�t�]V�K��W'���MFPk4A������o@�-����(���4|�5oZ�^��c,j�3Φ%�7��Mobgd}�?�u�lԱ��	-�p��J�l?z��Xg9c*������&�bq�$8�P��X�����f�bU!2d��m3��^#����?��+ѭ�m���̤u�l`yA!$�Ʀi��^o���*ZM���[2�^����v��w��»Sm��	9�۸m�&����r��9 Vl�Qw\�=��`x<��ʧ�]a��A,d���C�4�ݵ�(�wzo�QziZG�6y*ay��� ����̆`��(c@��N	��r�4���>f��n6^��CNN/���k����Ʌ*���|�)��k�o��]']9�bv�%�ȃ�)D��]��OQĻ�"j_��.ԏE�ɺ.>K�Xp���/�F�i�z��dh:��'Pp��j	���.��ۗ���l4�4iŅT���&�����\ǿ@UO�{ D�!	�B+��'����A�,��X�����#_�>����k��,�����(O#�����AX��S�W����ڼ��+��Y���w�;��p8 f�IO�� �J�QS�1؎W�>!<�Ϡ������kd���U����.�:��C#�☾��)�����k�8 ,��y���}B�
-�	��L�z��h��Eyg�]����8��)5�����}��o�l-C����">����(N� V��`7 t�̻p q�@wV:L�����m}`y_.箏�#0Ò�KEEĊ��K���wҒmb&^�(\��"S�'�u�S����6�w���K����v�mΠ���Np��\��Ͷ�m�n]M��Y^�@��u���u�w�;����)&/�Z���(p8���I��|���i�XB
+��"�QOȑ��ɝ?
�LV�8@F��9��C�R(dui��x��F��͡����0�N���ut,�91kJ�Bqv�	͸�۝�}uD�b�h�)���}����OW�e�[��\i�K}{�i���7ص5�H!aaL��<12����J���w,$<x�⚛�7%��y�Љ<��P�l�|� �ĳ����Tf��A�����;��^@"ǙoJx/ږ�8�U,�M�����%mJ!�'X���"'�,���Q�$s�f�#��b}\��y;���n1�p�݄a�~ _�Z��vm��.q��:���]��C�[�f˾�l%�;���sگ�����lx3m1$���D_�K�I?s��1?�w�}&�3PKط�N�,4�E%y#��T�ĢX���_��)0~Л��*p܃ �w?���lN��ԑ����f<�AK;��p�K�ج�J3����!=D���wA�q���"%��ֶfҝ��=��a��P�ȵ�</Xq|�ݻlW�i���Ɲr�x�)F�]�H���]}�#e��y�ǡt��L~�*|5S�DQ�5g�⹊"�.�h��[Iݻs ��~G����=�~,/�o3��7�3��e�H�nB�Jb[w'�&ns}΃nK�H�+�q��<2�$��l��e�*��`��:�c�\А{�f%	_�GEM��Lg�*�ބ,� Ws>]o��M�㈑���%P�{�S��dV$�� 82F���k�
�P�~���J�{`A)�e�k.����"��͙7�nX���p�|AN�OdO7>fA���	���8XR�1��������4MR�OI7�Q}��T@�HM���Ě1��Ht��Փ
}��F�B���N����[w���^�[�w¸����K�Yt��~s#Ca��~��z��{�	�����J.���'��VN�vǪ�|�ѥ8�q�ۛ��z��M��,=��).x�5q?����
�5I��	L�
c"�j�[���f�DԖ>��V1�sl�ˏ���3�`�񛉣�E�z�A.�m[��m]����N*)�R�ʟ����$}q�<��c!�%��Q��$��N�TG
�9�,�:����I&�Kꌁ��UR<��f�.�zYЙ��o�6[�(�jǼZz��!>> ��t)���,;*�M��'N� �؈���
D���|���΋U#�R"@�����ڝ2&��͇��
�op6���Y���e�Ye7�3EF�xO�c�_��^����ZS�G���e�j)x�������Ŕu�L旗��Hמk�'c8W�b*��ϵ���@�bXJWzd�,,���a7�J��?�_w�!����/eEל;���U�EL^w��ې�����v�=��xj�M��.���Ҽ!�����u��x�A�f�N��]\W�� ���b�0l�`�{�xr�%� ���Ͼˠ�T����1��*� 4��k�Z5��I���2pߨ������v|X�B5��y�ӓ��~�������,�W�{�w͝p����-�	��-Y���1	��5�Z���̄KF��\��+1���t�0oR0s���\����@8ߧ�	���m#B;��*w~�ٗ��N��zf�_�?�^f�QӸ����\�e�"9�_mC/jКV�U�Q/�pІ�N�ߣ0R�ϥd�,f����Kr�!�]4��+��j�4�u�C�Dx�6�1!hs�Jq�F�~���[��g�&p�ԫXZ{觖�.�	�&���ţ����2�i5�&0f޿�j�NLR4�9<���v��W�h�R"�#�<�X�Xj9auSc0���b�F1WV�5�⬚`�H�Çh����	:k�U-�FKXЙ/BO��3@�j�V�2H��h�'?��|�'Տ����b]�2gӋ�f�|��x���Z�=�.W�S�Z�d�a��#$>�5e���M@o���Z�����"B�J��[_{eb��d[���LY�� �Z��.5J�E8�f���Ѯ,Y#�0v�A�aA՜�SZ���!������ăBn���OD�Ը�x�������K��T6��*�y�1*���1!]�����F�����&�ʩ��٥E��^�Z��k��K�5h0��b���Bb�w���U�=nq��r9�D�� eEc�u�k[qWif$�ZЅ��D�8�ə_�w-�,�k$��F�@)�*E������W
>��(Qv�{��'e��
2K ���c�U�
�1�5s<w�d�K�e6�z�:t�����5����(�C@(N���U�&��;�2;�p�?a��t�:���'='��t"�b��Յ���ƙ������]��� ��S< �����D�`]j����z��\(�F�惀� ����'䆨H� ez��W�y��m �����\��7�*�1�T@��#!e޸��@~��c�P�(:��:���z��hN'azFqjbx������Of�|3����]Z��jH�/��Q[-<�2���}5N9�?50,��b[�g��#P�����ը�8&�D.�ʴ
�Ͱ�%ba".%�����H������,��p��f�/}WG�����(8�׹~�4�CP�^������k�IR9���/҂ot����R~�Nz{��vF�����ׇ�O������e�H�?���vi}���u�ss��OC�a'��]x���N4g�F��w6F��:=���������Bf�G��1/1��UW	�;��/t c^x2��,b��^�V�޹"P�q��u��w����[������O�4[�)�ϪJ��;��K�/ Q�n8%���R=m���6���h�Ѿ ad+C1��O!3��?�z]G !�*������!�I�Dx�Fc.�(z���� ���8#�w�#,e����OW�eu ����_�&���$L64�VX�&�?���-����W"�P��{���)4&�\#�#݋su�����RХ��K��j�@���V\0�[bHލ��	#��^~�~B(f�K�?���C�!ʥ��is�+�h�^yғ�YM֌�+�7W;�_\�n��ՒO�a�g��~��k�@.� 
i��p�l��ʓa�\d��*|)���[M��KX�6��73��>�m/�ADgi�e��M6��R�>��U�|�Uc���/���������v�k�̨�@����_F���3�f����y'ÿ��{盘b0����,6�a��
��?!(��ѳO�Y&�h֏|4�BƲ�j�;��b\v.����#Μ�'%%v��9ʹ�ހ�N��i���nډ�+<���F�����XI�?yză�|�p ^�ts#�����6��J��`_]�� ��z =��H�W+�S������6��%�/e"c���A0Q4[��C)�F��=��X�������������UĭQ�b����>܅����Ո��[6) �[�{'y.^봩����O��;��b���P���g�k)�V8}$GŒ������dg�!.}F�Q~�X<���*B� )զ�oxI�a��������U�U�VѤ����9O1�S�Q�֫�-b����;1���}�f�1K�h�����;��$r��B\Б�\��Mw�������H��J�Mx}��f#��9�K�:����'i��s�d����c��u)���o7 9��VJM�����_!�1	����� #����������[Bh{�ސLx�"�IhL�~35:�	��Im�,���V����#�Q�1=|�蛶�u��������ʭ�'ѻ7`N�	�����j���F���\IBĈ�3o{�x`������d}�9G��*"�z���-]��6=�h��=p��`�r��u���n��N3�q���\G�9�sL>��ۥ��WZ�l&��y��?W4�-�0n� ��vSу!d����2��YU�Z&>Q j�U���=�c��"���z/h�a�~�:^R-��&���o,�j/��9J�r=mZ��6Z/��b�6)gp�n �'
�k�f`> Z1��iЋ�#W{�q$e��)ʊ�yEٺq�Z��ߐo��i׵��?���-�G�Ь|@�G"�,n�����E 3�X����܍nCd~v8���>0jvx<��r�4L�,�p:�^�@�c=o�F(q�bU��l�Q�\���'�%�84o�a�X)��~����#��an��l4]U���Q�f(��YG*,�B�|��Z�ٛ�PJ�� ���KX�H�}�6rX�If��pV�H?���VᩏJ6�S�?rwFl��cIJ�w���}	�?����w- ��$`,M�ɷ����O�I��$����r�vH���B^�!����·$�Ju֔6�jc�&
eG��k�bz�G[�ޑSS2s�-�9cBX�i�ޣ�Y����A�9F9
����{��0�~�1U���5@���M4_�����%�H�w�r~�� ��������C+:��K�����,[H�U�?��fHx,`I����e���Ah�@�O/r9&(����ԑY����k�����d�<��s���O��̃�4�C�i��l�jm��ѣN����?Ѱ��ndhr �M�)>��F&�N-�^z���[:����8�0q�B��-��a��:����>�)����l�Q�X�hP����|x�ef�5>��`���<j�������P.D�ɣy �V3�@�U������$�s�f�#�?eoVr���<���:�j9McG�&�dks��Py%�����e�u�t<�7~7���Q�O�]��9LH2D���2�U�T���2T�/j7���fA\)�@��qo����M�K�߱�e�$?�Z�u"P{��[R�r���)�t�-(��ڥ���+����`4�f�d0}��[�h���?�X�j����:��.��t�p��L-���0S�Zڮ�O���p��}cJg<
,Wf�7N9�݇��mb������G/y|�3��u��@=H\��W����,��9�a�
���#���E��E�jS7C�f��*�����@���)����vO�[�U6[�q��r4��:x� �X�-*�5���r����8<�~��$��u�s
,�H/r�n���S>9��l�#���cmG�q�&d�7�7m��N�Ê��;%�\�`*1n哢�}BټH������99���gK��
��:��K�k���A����/�3,� +��x�|���:��B����������-z|O��P��L��1�v�N�ƚC{� ��拍��i��7 1���l?�W�̡��A�����1�)]S�J�S�3��}��p�Z���i��˶��!	���/��s�e��>� v�:�w�[��=�gg����
�*L:�(&��O�Q�N��~�1EE^2���YR���JH��U�1�,<,'zK�l�T��-�1 �!��1,�*����nʐ� ޽��xpX%�*;C��;��-��t(+d	��q�4h��<�TҶ?�1��z���[���\���y\�*[��l1��t��;<W-������65�¥Y���g6Ppx_��X���+�C�� ��슻�tR����ya���h��-���mW1;�U�&�ѣ�68������#�1 �.iwe�?ZMH��W-`y��\5�?���ڰY��@%Ȍ�)�%�'��T�JV]V���܁��wj_�c���IU�B�,Vp���G�G�N��}m߫�<���ݫ�Ʒ���ǯUU��c��!�G푽fS��@�l3
{�G�d�{M�Tܫx�փ�.V��w���!���$);�>�u�dA�[H���X�>̲��"g�K���
��l	~/�m4������@r����VQ.�CG��^��c�F�%�0�s%%��A��1,:0s���G<��|��Rib(Pg��M�e��`����|=�9"<9|Q��L�~�z�:�=|LL(���ҁ��QF�֐֚�Y}r5��=TS�x��16��:PM��[��V!L��+��$��9`_@��XV�s�&�0���þ���T���=3��qmN�����l����ϊo�p��\,�؏
��w�0G �?~��f��E�	�f��!�o�խ� '7wr���&kKF�(V�����Cq���� �/���@P�{�M�5 ����5�H}6M���,e�`��	H��+�iR�q�Y�#j��n�+@/<f�BA!����Ij����6*Y�j�I���u����t?��.�:AV�,�݅u;^6Ҳ*;�0�a"GC��c���M����ky��v��_^��fx�Z���,ׂ<D�;����
#8E�E��Sa�S�L���`�w�����O�q{����ɌD�[��¦z�,�&F(�����Ӱ�b�k^�]�M1.�A�MeU���`|FBT�ۧ#�n|�9kEO&}j�1P�9 �E󋽥ɂ���ʽa��V������Kry���Ȧs�L�v7�Q��I�nD�
��6��ϪJ^��I�Q^*X]���-�ތӣ;��0�շ̦pd�M0̩������o}��;n4Lj��Loh��b*�~�ϖ�	}�)�G ��D���y��O��L��>��kD�b��gj��p�&ǌ�S^����mC��N)�ΕUATx�.T�nR������.�S,Jw1�J�g�uT�Q�W���YrPPZ̟SYO�j�Kz���8k$�j'f&X�Y����L^.���m�!�{;2WW���^��H�w5 �A"FRrI}z���R`q���%Cn;`���;K/�a�����}n�V	��Ǭ�\Yˈ�������[����
 `���>$�t�Q!@��D�l��=��b?Í�o��j�_t�8m��5�����Y �-;ܫ�X�2_�bpOH��"ـ��� �V�A���`���V�M�]��J'Ϩ7��T��E�1Ss��R�#�����$���V7O/~�2��͒��[3%ה�򞽟�:!j������~�[~��}K�	m�jڭr�ÿ��Y�]9��;�d3h ���m���s�#U6SG�^����G�G���X
��%�?xv;�1A���l?#���4�{6,H�����{�l��4ܥ;}���g�n��;_O�����V�J�\|����GsK�#X}�zv���+Ѷ�V�[�xw*�Tj#^�U�o�D�  ��,���r� 2'A���ńY']b>���JQ�5WW?`s�aq�m��$U��(E9��$�D��N����Ő]A�A�ɨW�@.�-P���uQ��r�(�ߟ�jF� :��;f��V��ל�������b��ӜM쬪�m\_�(���o��XVTU^�L�Q���JX�{gi�,��5�A�&�����v^�G��	v�5λ��=�,=��q|E��K��`�s�f��`�<U,j���]"{\�t���lo�p�Ξ0��U(�Z}���(�\�=+x�p��փ�#�U�̿+��O�T|�o;'� ��b1I�`
�u���H=�	����A�zM��6QQ�5��'2�)��o/q�7w��u�/����;������iC���I�\P�.���g!k�px}�g��o?����/��5B�X~#�����G�(�a�A�扌}m���]A��T�W�ǂ���V���2�;$LH����-8��.�&B�-��a"�2�j����5N�F�P�-��#�����i��)@\���fp�7?���ؒ���tJ��� >�B�3�iU���ҧ���6���_M��VW�"��%�2�� R�����q���$G)���U�j�8�:������³�~�,1n�\�$��٫��0He+Zb-�Y��:���	��ے���̅�����i�A���.�u�9�-z������3Q����a\��2g�T�?Zk\�׎�A��,��& +|���,
�s�_���e��$�Z�#H���/xu2�1*��$/�dc)Z�I*�/�!k���6u?��Ԃ�U�Y����j}A2z/7q�v�ʞ�;9U�V�u�x��tό��sdIyhRv�,:�5���%��������Q�i�`���@}�|����L���0��Q���s�ep"��BeJH��[����v��ө��}/ߠa](1'�|xޭt�2 �����Te�7�Y�J�S���W�T�agۮ��!���Ug�4lc�1���k	�)���'p]Y���:3;�R�K��qZ[P-Q#y%����Ó2�������D�{��{ۧ�����=�7U�ǯť/<B�������Xj/D��P��,���ݖY�b��*F#m�An
h6l�|4PJu�wo��[�H2v9��o�9!����\-9 ?@U��&l�}ƛ��t������./�L	;� �E&�X3kgʶX�����z;��%�U%j�|�ƈ����K����=�T�AVÀ3#bsg9�؟�Դ�ƴ��"��G�8�P�	�6����`ꔮ(����c����� ��-C��\��dϲ��MFm�0I�_ۛ+xe��`#D��_�)�[���ۘ�M��q���s��-��߰��}���ҕt�S��<�Z���jB���n���Mu�IIiU�}3[��ʺ��Z��.�X)����$*�f�m�M�0q�_
��r���3�8��ц6�d��l]�6+�)�¼�6�&50�G*J��Jb��F-y޸\т	 �Ok��#���г"����?���dq�z	�-vcH5@8$w ����q�ҧ�_��'��õ��D�\�T�� ���~�ms�/ U����M��P1?)N�85�H�Kh]�0��[N2��K���9ɃPB<,���
I,�1��Q�^J�������� �r.�|�����(J�d��oH��:f���U$O�srv�b�h41����'B��Z�C��e
Iq��z�ΰS�Q���0_{@�o�>h�V�ѣ�b6+�����q%����1��6���>ׂ^b�q�T+��_L���K�˯g�h�#D=m�vѼv���j���I��N3H]��x���0�証��V#H�C�E�[n�#���>F�?#Al�o�����`���t�\^�Sj �e�2�FP٢�e�T�!�i��Ȭ�6�O��S?I���	�K���.
2|���v�������;@�4�5�7�*�/��]�/�wN9��gB=�&�Ew™U,�hJ[�K�tj�W�
��m�1 t�Me{U�0�]h�cC��s��������W>�A��xjG��F�ѠS(�2�M���A��tQv��������C����e@Ao�x��ʍ�e!��i�h��~[��ާ��8C��z�����g��y#�lur��avx-'��<y|��{�"-H�٫7o����r�Cr=\��;� m�>Wv���x�iYY��6���ԗ�c�FwƯB+c�����uje)I�{ �x��	C�5��������z[�C紑���3�&���*��@�r1�q�+�IboT�2�p���>&��4�:�M���&z��~��x�4���������NH�������$�>c)jNK�L!�!;nJ�z��]]7��>s�*�垚!�1�R~�*��q�7|^�:��F���I��~��� A�����'?4��u#q%��'Ũ��] AY�xhJ��U(�"K�Lh��a9��"���l��?��|B�$����#�L�}�Ta�KQ����>�"��9�����	�<O�ժ���}�����,eC7:�ˊ��}
$Fl�e�mD�B˫��$4w���R�c��{Y�[��/Q'�%��izw�@iX읰3RE��T���'X�`r2��<͸]v7 o-�#�2p��VS�<��c�^��#<���D�B������,>�'����-�E]4锘,:�[v<sM|�����w�d���h)+�[Ņ]�����a�s���̓�0}!�by�.?�Zޗ�+���
l<u���B�"�ڃ���"Yr@IA��(1�-r�S(b
��^��D��qEz��b�n�*�*9�j�)~-r.&Y��l����\{��2�nHKw1��'v�r>J�R�e�ٍ�A�������9�IT���A"yt"&g1��!�{L�Nr��a��p=/2qv�����orv �����Y�zr�{�~�rV�3��~˟oo��a�S�����%!nE��BG%۩�}�`�RAylc�P\3w��y�%8�h,Zh�-[T/��}�.��ڜ�@(@��Mm�	M�N��K�R���C_��x���sg¥s�N72�K�#��W��Y�`\�xEv�h_�q=���+�@���+bl7M���I#���&
wvQ�*7ݱ�y��'�A<�����C�م�-[�P��8�e�ӳ/0[��������m䙫ڣ��N֫�ԋ��.$a��[y���K17D+�k�
$�ܨ�_,Fl�cA�~[0C�cҵ�*
E�|38)��O7���m7"��O���Y�?�D�:���$J��8�>~�|�d�ɢ�n���Hh���%�$4�qp0����m�Z��P�	��z��*a;жD£:�b���p\�O��S�a��ځ�Rt�9p�(P"ڛ������tHbĴ�OS�"N�}�Y�K�s
q��'Û��C��f��Q�4)e!��]���%�>;Z�${~�q�m�(������V�XE��vd����@��4Ǽu������_c�o,�V�A|3��*_��`����Mi���,2 ��Qy�f~����O=�!���;�z��M����MO/o�{�Y��.��F���vJs�kC��P²�7x�M�J#M�����r�	� �p��/aE�vy{Hk����ܤ�[Ǒ�A����z
�e�{�>�; �[�SP|o�Օ�d�U6H�Ǧ�'�	�"�\gRF{3�9>19/&� 6���Th ���a��5��A, �!�N�P���i?$@=�Y�1o�ﾭh��nP��d�8��@��rJ,�5-��M�蜕�%����q_��7E�}C�tw�RD���[c�#Hu�Kf8�TR������^]A�Ȋ�e�h�'�{c��]00Ӡ��\G��Ѱ���K�Mznd	���^��N�9 /s��XR�&�A����֙��m��)������@��@n
Z\69�O3~5�N�͐ W����d�v�>�,����w�*@a��J��/���T����l��_���V�/����/�؉���y�k�����k�_ɴ�t�'܍�*�f�5�h�2�:f���e��P�C3�
�K��2<�{oMm�}jY���<|pA�=-��u��(�f�X��d�S������FNo��K/@JA��Ml��!�����2Ӿ���N�6Fͧ?�yb(�TAOfr��5!&n�i�_��P/J%۽�D����άb�w,�8�a/��b����0�P��s�~&���e:�� `}B�`�w�'O�ހΥ1��H�!�c��SCV�7�X�1�<y5~Qb:�>2*���v���S)SeJ���e��ƥqQ(�5�1@������i�,8[��P鴬/p�-]���*a���s��6�hx�\:أ��s	ؒ��D@ n_1!���C���9��I�x����j�K�|IP��v�����=���YcD���5�m��y��_.�{�(o�����#Q2h	ط����|���+S��+A�<�#ܗ��L�-��SűF��1Xg���z�]��/��`�ؒ�y2)lUK�,�͝�q6��w�G�KE���$�v0(d"��*a��r>��ya浾�7�a14�B<`]J̎��I܆4�oAm'�[���r��� ��S�$F'@zٖ+�">G����1)zE93m�bn��%���*����՟�x��M�`M��ʙ��^�?k��7#��v�ֱ�Y���yB.��\����I�SWhU�P+p�%0��DU�xzq>�i9�6�'������[��U�nR�	�7ê2:��_n���D���e�� 2��T0!׫x�	D��-(�qeߵ���^������:�B��4��jg�Ńp�h�XtɺcB/���§�Yh��u���١�֓�s�R�m�2-m��'Y�N��������@��O��wR����6���NNI�ğ(� y˵�k��E����9��m.p
��I`3ʫ$�oSd�����a_����`�?�ܐu��+S�����C��.t��A#�l����ͺ%MբE<t�#׼Θ)�}YyΓ���UF���*
T��ù�j�J׻/j!z
s�a��4R;�)j|�I�!~�L��I�̦vJ�Ӟ�>l�M�a7�o�υ-����3��,�wqL��o�ruI� ��'�*����F��c��jM``B�|��5��4��5s�͕Q9�U���w�j��\;�U�vz0��bp� **�
���)�=�~�n�"R��E���XB�U��;�I�����S�!�9艹�c�.�Ӗ��)���˵�`�Àm�$��!�G���-��hd��̎E�v��^�����-;JU�9�r^�d�U��ɥ�p��k�@���r�����D/�co�����Z��N�U|{g�|��Q,B���Ҏ�OV��R��<Pq���PA�H���J|����i�:��T�H@��00zb���w5굾��u��i�ӜQ�c;�������_���q�4�.I���<��.����%�6�N{ �� �n�Ж3���-w���P�R�m��FϜN߲w���hl̈V�ow��uY{�� d���B0�KdT�5h���gt;����I$�4����^�F�|����_$�t�R~�I��1���X �� ��w	�E�6��2��Ӛ�@�,���TH�(�h�;{b�}):�k���"2.�4P�Vy$M�.��B�,T�G�v51ǳB�*AR�7�q���x6(�mD���%�)cv:%,�����a�=���
��+�*� W�jjd���p�����EBG1���E77�ɟ�B6��P$>�'*�pO\�.$�*�����|�%x�s`bgg�td4u�2~�/`�O�Kg|n]�Z�3^�N)�����a�(+�o��\/a���?Q������:�i�������x8E��ݑ���,���p�YY���ȹc�n~城 �����
�cA`r~�9n�aq\��ou���w�\;���#���l����9������bg;����x�K�v���|�)]ϲ�H-�K��!�^S�E��+�tQ:�S+#?��Sl�~��R2�]Jn��J w���q#hJy�!o����E�q�8i���Vo��%UR6M	�z�~Zy�~7+�<R�|XH}[e@����[��czO�>?[E�"GD� w-2����4�� _q�sD�б�c7�[��x��C��S��%l L��G��be6��T6(�F��a2�a�H�c�x�8@���Ⱥ��#���2����[;�A�3?�`���taΨ�euNf��3� 4�c1#5�gX����9���Y��X԰�y��T�E�i+2�T�1Oĩr�
	P"�.s�+�Uܙ�R��ƞkW�#�U�zR�����(G��~N`�YV�ǵ�2N���%��8�?c�u7� �^��E�	��x�ۼY�eת"�0[(ۮ��$G��m5�<�z:��:6�j�?l�Cti��QQ�6�%�$�$���}R�$�x�X;	�J�ps�����\mW������*C~�Q���I?�tf��?d�C9�Rƾ�V#5f/XX��َ��+���(`��*�)n��G�����VW ���7��E>���lB���y|h#q��cg�-1�>#uVz\�A�5��E����pՎv�k�g�m�-��C�s^����~'�N����\�Pzۡ�5��L#�ks���g�V�[`O_f���3M��)E�@F��n���e�����&R�Q�����iu F�MWRŰ��P���6' �$�h�~6��v_��D=!�!��ϓ�,y)	��Uۉ�עD��>�U�㮄k�Q��#Ӂ�!-BѦ<���U�{F�G�}�Ƃ1\��s��X��_��+`)Zt}�?#�����r�f�6�*(�C -n\�[˔�%d9�W,��r�N0�����І��9�|����o9�ST�	Pv7����h 0Ú��!iȣ8��̱e���]Pu�s_>f��3����	k`N�#LO/�#.T��{u����4���b���}�~SW�(��=]\C�"�(xѹ��e�� <�h�J�i�u���ܨ�����XϽ�Tq �;��T��_���g1�CZ.�q�eϯ��'��$���ڧ�R��c3�d��
�5w�@9��@��U_ۂ1�1���4'�+�?1�e[��g��Z�����wQΝ��q멏m����Њ�;�ƀ�<��<���c�*��*��Ҧ��}$���k3�qMr�e�ޣĝ)n��,a��e�Ku?���s���(�A��x��#5e.L{�� �%�2���!��p��zM�.(Vk��rh�[~{�����LME�I�+�����Nx?��n��C*��(���
okEd(���: ����K
���N�#��T�^�k3�B�j��ů�I���ՙbd ��қ�< ��g@����K�_M*&�(S�m|"�óg� ��T�kX���Ɩz��w���k�7�Ĺ2G&�Q��{�!��6�v�Vv�a�8̰Y��5�1�K�����9�:��I� �$�/۫p|'٫�����:�ߟ�5�#�~K,,Ԣ�b��.ݿP���8�5�FzU�����f��X�  E��Q|u|�L�l��I���a]�\����JP�FqJ�壪���ʥ�M��{��K�����QA'��,�h�heZg��C>�D�g��=q��8���t�����+,v(�ɴJx�ᣇ��]d˨����s����D$"�N0fQ��>D4�\�q�A(�fV���	�Nc�9�,��/�mF��/έ�$�rUC�'�1�| �8���$cy���V�U9 ��yt�Ҁ=DE	;�����
U�3g���Sc8�x��/g2��?tB=�m-�]�h|H�X�<�`a�L���x2��XS¿<ؾ�5Xlݮ�9
	��-�<�+q�E5R!Z��y��+.���w>����M���B�ol�=j����0�u����%�����"y��	wa�7q��O@4�ی҃j�Cu:���'C�So����R<���¾9e���4���;��2Ƀ+�;bI�2Տ��#p~0?�\�-�P��jB+���ַ�4��y�sต*޿Y�r^��͋ڏ�?�^����js[\$���ě���A<�Tv)����UQ5�uh�Ԁ��=��7^9�{�3�,!C��������'�����G}�0m9}Y�����0�ʤ�EZڍH�陼5�L�#��%�nS���(%�>5�!��3�����Mb	��`M��O Û[k���)TW�97ۦ�bi����9k��bn��̨ۉ�-�c�B��.~�9؅5֫ ����`��u��1��
�-h�z�3��@;k�S�����^<��ʫ,�� ����]8���Θpe
�Zީ�"�P;yaɫ��lO��*�4^:	E�*��L+.݃@�'�o@n��t���
�+3S�7����q��{�_�Vc�_&DQ����7����<t��d~uʸx���-���F#�6D�f�S�%+t��n�0?���JR{xҪ��M4��-�����U=͓�bUE��O��$�rg{:J~�Xe!|�B������/��H�8��4���w)��D�����|MyZ&�F)�ۿ�2��*�zq���Y�_�1��=Gp�/��\Ӄ9980,0VP��*�g
Z��çQ���3B78���"���	�V�/����k;��[�����ek%�Z��E�u1�s�|š�yȲ�?lp�>�(��71~�Y_�q?����Q��Xq��}"�:�(m'�$��K].FWW�4��5�H�� ��Li0IK��-Bq�1�f\��5�փ�?�`n4��T�)�Jؾ�J7�Oii��M����2�M0���������#�3?��k3ǁB��4C�������hۑpNS��2��v�q�E����w��!��8��n;��Q�O�]�]������0�*��3���/e�Ǌ�aVog��MA��MxD���^���:��jf��y�ͅ'�M���1+:_��|�M�q�s���+�$X�:�L�p�dv�5R��``��H��Ii~�'�F|��5�(Vq	`��۶�-�¬\���p�����Z� h�6}��O���8/M@�C�ʌ�|�r������oQ������F8A�M����q��-���]��X?bUX{����4�:xA��:�`܌ll�����D2yٌ����4��b�w����߁4���M��8��Q]��p���hq�%��p�i�+�{����ǘ.?"����d:����Av��]�u��է�w ��g�s�L7�`�,�w6@��a��bTئ��	z�p�M#�bJy��`�����%ua}�=���۩U��ce��������#R[}�Yi�sJ6�$��"03�<��=m�o��vUT_�Aav�g�u8x���������Q�*yh�}3�~��:[Ѕ��A�Ժ���F�{���6�nvǢ��� >@��|�c����&%�Y%�<�|*��j$�1�	�&ŏJ�$o�ohb����)(�v`�4��U��e��.���N�{�,i���؃�r��gA��`��ܡ�}����@���_���_yc�;�g��|�I�hH�P5��PY�=���BE��l6I�N��y��M���i~�&�N�������������'
�݌I�P��`��I��T���U (p?P������NVS�.Zc9�	�$�Kׂ��L�<�{�{��Z#���P�OL,S����rsp5�ܷMT9�4��F��ϴ���gen� �����v��[��y��3)e�{X0��b,��`����x7�܉7]$�g�"��eL/�}�Ps$.t.�X��CEĄS;�8S�q�����V��w#��nˆ�+x�e�Ba�̴z!�}��?A��:���;N7�����ƶM	=�`yM�	̡�2�I		L��b����S�ь4�_�P�{�)G-kn:�T��A$�CЉq�C�y�V^� �(��q���:��Z�
�7������w �} ��VpT
ʧ������>�3t��)U\m�1<�b�К��&�7Hz�����Z��f�0h�H����l��Ո ���v��|_�+P
�R�#)��v�>a�Ն�\ۇ��n�wx˜�6��D�K�c��b�RɅ���`���B���E 
��d��zV�(×����g�
}�>gRZk���_p0~Eٴ���g��H��K��z��#�x=٨^��n��:iRrf���G_���1�q��0SȎa�/؋�OH��>/��Ѐ,�w	9�nsF�M��[�m���؋:h)�@��z�#o��C摒��F-N9��F�&�!H��d�,�o�Z*d�����]^>8�;~D���Y5�X��|W �h�{x���L���ӃCE�Dk��6���㚰ʈ�.K�g���`�5�JF��HT"�-�&}r�;����x�ÕRo��/�G�JY|����2�7�O�&�j�����H�+8����_6��َ�%���_t�>�H��1�¥77�ɶ{����cn�kLR�4z��߸�73��������覍fQb�͆AѻV�����ìV��M8ٍ�4#)f�
�5]gfp���m֊�^�=^b4��N�D��P�7����E�,b�y�����q��a��O�yb@#�I�'p���ٚ�N�z���1��r'����0���k�%'��	�"[ڡ���Y
+��
o߬�����U�r���G���5z���H>�R� �2I1�M���y)_%ug�W���� `$��(9��F��.�r��f�1t{:���@�7D�Q՛jl�L;���㩹�*��r�̲@ ��N2I̿QŞZ\ޠ�����0yuR�}E�K�ڌ{�FY���%��;���E�J���R�}���h%�ܙ�ٜ�j����C?��I<�c~�D�~r(��~��-U�(\{�ӊ1�3G;�D��H�����{���p� ����G��^�nɼ�ue�o6Ev{�!��T�EF2�!zSY�
�_"1��N.�z�<�T��1����磸Qu�[�|J�0E�J̓&�~�z�w�:��a�]�3�T�t���d0��Azl��-�T`-k�ճ���,m:�:<�@��E�5��SԪTr9�r9
���5q�K�4�ھ[s*M��bh�0���b�
�
� +P�1��Ά\_ak�[�H�vL��i�J� &`7��G�T/[��c�c}U�<����Y�2Wy&����<�K�2��	W����e4+�wxe��M6i��Z2�Q,��&v�[��1	�TK)�|;�	gn����ʒD�|�����P�V�حZ�A��CW +m �t+RT�݂�����7�9!��
��l��U9�~������Zf�Ex��paK�(j��&�|t+�����#f�����"Vgd�ڭ�ϛz��pd;�7)�k(���*���W|�d֖�ZJT�L3.O����\8�Bp�J�y�y�1���\�'6�V�e�旺����W�!���Zf,�J'��g�� @����p{��1.(��n��8�|CD&S��,+��%0]�$Gj��N�&�Ĝ�XQW��X�P)�V+���{�y��4��zв��ġ�-j�epz�`J	p>�n�i�SJ�����5*xS��.��잠�h0tF&�%oVU�T�țQ�x�6	�.�4�yd�]/N��P5}C-JxC8�6�k.�g�|}Ũ�a����z�������Ygn��1)���oIC>��k�E*Q]�p���p�{Izr���*����e}�@#�"��r��Y�]͹7�/�M3��,�8_�r�& �A���<==ȷ ���������̺�);N<vV��t���(�iҍV�Nb�G~���}�܉%��IX���|��J�;���C�Ҍ�lu�K'�ٿ;�%��ID��
���y�Z���������Vgz���Ȗ��Ts��u	�I��B��&:	���1��͢�Z�Dm*�(�`D�)��F��EikZ��V�m�G��Z�YO۽]�`��gw�F�F���R�Bj_$Tv�"sA4�LR�e�@�h�#Gpi�ȏV�x����EKt\��}�9��;ϝ8�=�������Xv?4������E�4�D
e��/��X߀��w3��&6#c�.���!񣶨.&���e㞈s�a��B�EÏ"�b�`�NP��������!�	5���qJ�2�������%�"
׆о	'�_;�V�������Ʃ9�Nd�[OJ�� �B���C���za�LV�Ǉ �X�F��e� ���I�]�xu�g]S�L��C��֠a=��9d��s(� �G:M	O�~yd�����<���y�?�BG�?U��ᏂP������m6ڐ��k����&���쭍�6�
_u�O^������,��щ1��� ����g_�ag�z�W8.���z���8�%��l��� �揎V��LN �~��#&��0���/Q����*s/�c]�� �u	_�f���^l)�8�Ks=�~�$:�����}���'nb򹇄*��ô��0z!����UF6Y�53%Z���
ˏ$�e �#s�}�7'�`U��+���.����z{Dpֱp�4lVp����fd$��mf	�<�i���[����-�E��ҫ�r��ܛ���Q"����� +�|G���(��v!�[vqf܀3�͑�,�¥}a��������I�h_�ew0\v�Q��3)�"$�S@�K�+�ώ8h��>h�b���� ⯁i"��]Z=}쐿�-������2"#i��`����|���s+N�c���l�io���JU�&����뫝u���������:k�M���11S4�U8-֭�U��ɝ�m=Ta��0T[ѣ�꿑N�:����X��F�0M����Ԇ8.X��}ݥKځዴ��{�a϶"b;��7���4�!冨����N��1bu���lt�4=L�i�ת�<iq5����9�ͳ�J���x !�I�v���:J��t/����zmDs��4�iW3�a����+L#6u<��9���[����%��Ls�2����y�ŧ���������c�p0��̕�!��ʪc�g�c�KCʊ�Q�u����ǐ��X ��O�>��n�GG\�)���W�zT�B��s���{:��G�����3�[�`�Q͜���{B#�݄����4�*�;N�,�k+�<Du���`��C~O���;pJ�zAQ�W�"�D�E�?-!��Fix�4a�T�U�jN��Zm��/_ZѺ�0�I�q�s�Ʈ��y5��|/M��؜˽�=�o,�1O.�$�1���`P��,pZ1_K��n����k�)���e�Ol_��ܤbW�/�6�
爀y��o~�X��},ɡ��Q��D,OSi)Te��y��/Sv�{D� ��<��_Z�G��r��28�Qr�2/��<4��g`伱���O�-LW��]�G�)f�t"W{��;4�k��_�����tT-����F���T��!C�8�j��)�}��V�ȱq���`��=ƿ#]�"�	�9����'��:Ip�i<�	�h���Bv�����q�_�^{�������u:h�<ӊE�8���;�n❄F�f2��3�K�z=�t��if�H]y�D��ۭ/�IfE���✮qU����AFֈ@�y����/���{��R���냇����q���>+�}�k�Tͷ��]:��Y0�V;����UѢ��$i�y��SK>����(xJw@�@_�o����FP�����*�����z2��N1�6`�]�q��È��ml.�>)��G����`*�e�4Y~�7��@lE0�2��ƛc' =���2t-:s��I���M�{�r�/�ư2j���h*$�/s�c�X���(+MS�u�@�Uܫ��=�����A+��}g��ݦC���d���賙V��Rw�A�.E��"/)ײ+���9�ã@1T�5Th�._�'�H��75C�3ܼ�P0g��u���}�[��Kh��r�
929�� ���qn�����ep�@K���3�����7X���r�5�I�+�e@�ۍ����h�7��ī5����U�<M��a�7��lj�Cə����C"�q��6Z=�|8'ׂUѲ��񃙕�1<�.P�谏��!��M�T�mp.Z�x��L�ǸO3�a'?j3�&2��;}�68�����ă�O��1PQ�C�ނ�y�!)�W���1��5C�Q��3Dbz��u�9�A���e��%<¿�:"t���h)��&�𓟹rb��Ł-MP�P�HPOb O)c2�<����`�1��5P;
��&��bt�*:��P~����t�I����)h
�@�
K��Ä���{�!\HC%mл�*J���EC���/��5���Ř/.��q�M[��g�PM���fD�`n�8�/��,��o���q�{��<��g�:d:�-ÅՅG�oI��]U.�n`��W���w�]!�(<.cOVc��V�Ė3S� tg{A��}l@�ЭS��vi�+�A����tǦ7K��@k�Ff��+,"����a����UQ��j���>�F?7��~�S�,R;���<�	H_C4��%hu&��==C�(�g��
�-+����z�q:�S�vE��
O~D�8ݬ�k��=�`�ZvfH#�U����C�8�$����o��E�2G�� ���a����}�V�1�'��F�0�m)f���`[8K��vd��/�)
$�*V&����hs�\�%&��Z��4L�^�����N.��l�W�h�v4{��ɐ��S�Ԏ�� ��ޫz"(J*�t'�5��o��3{�p^M�S���A�`��|L�?Z;����_��������36Y��f�A��[�"��p�z�k�L��s�`Odz�J��n��JD���g$�_.���&�sG�z�n=�����F���1B�D�y���=��٫Oq�vF�Q|߅�ֺ�����������y�I�AN޳vRU)�*��%�����āK�0���,?h̦������מs�o�-�=���ϭ1H�h����|O�����R��y�K(��O	W�5�>u��Pt��U8.��t.��g�g���?4�&ф>�+���V(���a$�#yk�(�"r��~��.y�Zq$[�<66o��|~�/�J���p>%�{���ER,�AF%UE���~��4=�A0�IH���<@���n��NxH�ͮ���30�rn���h�s��Kf�m}�ǜv�kNi�$�{�C�B��#�cE�9o*����:-l1����Kn�	�z�2�Np�%�E�^��^��v��"6c�2����p�F�=��&�!\㆐#�v�:���	�rzi?�י���\���ޠЖ��&�m�("A	�	A6y�4�IΠ��Dh� }G��F�1��D0�)�;4Z
OR���F�z����">�dĥ  Sk�'\N�2g=��|7�Vut��%�?\�q+=�8��T�	�Z��C}
���L�K^N����ng�UG���:�����᪉�t_YJe��.j��b�w1���kd�IBh��
4�G�xB�q`�k��4{��SgP^�Ahڛ�z�r���*b���"}0��B�A`�{do4���:���ѬyE�Z!�$�Gl��r����},�B�F��q����3z�ϴ�xV�I��6��'+*��񔬔���},���4u��u.xk��B-���U^R�I�?]��[��O�ӀZYi��
��
/N��T��%��6�k�G؜�)�^|1���4��|�w�9
���]�5�6�A�p+�'2SC��	��S�K(�����(����T��x1A�Jiu��a��%�K�s��{�D(�X.$�FqЪ+�\��ڦ(����8s;��_0��%���]���ɚ�s2d�FO=r�)S[u�����|Tʰ���"�t��z#/�3�O^�;�R��S^�\X������S��Py��p�|���sh��|4�6���t��l��t>�!M�b�r*�0ق�Kjn���f+��D��)�~S@G�b ���u#l9��x�F���9��~����O��B�͵źRzQb2�Ѧ?�W s�9a��(9R����X�Cb8������{�$�!$@ߡq�1�rWSU�\�Z@kg��[q	�G������\��9j�^����W�;q,X��#�6��B�ԯ�[p�rQ��r��v�b+���(QsI�gc��������o5�L�;�W	xy���:a��}��q��+��w&G#�+>���nI��YZ7:)ȥ���e��:�	f�'D]��V0�K�5ھ��#D$��\��=VL,�rJ���&S��e�q��6ݷ�:���Y�&u�6�@$�?j�}Kc���[�~Œ�me��GP���WK'�dv��=DB����F8R��ע��qz0;}��^�*��\�I�X񯾙u���"�樼~���ĄB=���{
}$%� ">d
h�'��hɣ�H�.�w����e��e�Ni��v����Z	j��"��Ak�fȏ��ڒ�!��k�o{�Ŀ�	�'zD�h״�D�)�Jj�W���-�ι"Zڜ�L��2k��@t�x7i�T�<�*۝gF�/_�v�,�*]c�?�(��M;���\=�ew�I>ݰ����~ i���{�O���#�S�=v����$R��ܧ��l
x#�
�aI�L���GO��%��nq�
�����p!����,�H����*�
+Tax��:�v9q3�bӽ�"t� ���M/3��w^��8C��5ʀ�ps�BN1�?���єCA�;Ł�]�JxR��2���lݺ�G�
5�<�1���x��qWr��Owx�*�7�!�3�Sg��u��2�3���5�1�����i�q�S�C����9�K����6]4��PqBd�*���	��q]����-�B#�_���鵁�W� ,3�.:�ȼr�Q�����6PK[����/��E���w��9؛b�=ɝ_�q[d4烨c��܍Do]�%]� 5����>Qu8�"�C�y�������0Z Y��$w�k��GƆ�dP��RŔ��8����'#y���&3.���*���i�3���"�I�jQ����,9��A@�<OŞ�@l�L�R�
\ʀp�RJ^�5ݿ��|{��9��[��IS\Ȑ.0P�)�s�;c���QN�t�E�����ڍ5?�q]uǍ�ί��{��637�#��To�fӳ�t"ߜ)'/�d	�o��AQ�1sm)�>�lէ�@�uE�������8�b���!��K�Ե��P�*� ��pH�0��`9�j�z\��U,ZX�͵_��Vj��P�g���T���\U�k�� �PK�rnr�
�����==s3������������}x�=u]]����Y�XoΚ���u �{�0� ΋�F!�s��k��'%D6C(��P$�m�P)]T���)+�:`��OUbJS�-��5ۉ�'�7Y�����B���z�r.��Q�'L}��N�#"�A�&I~�>w��v�|���9�N�1݄M���[r�@�gմD��֒+�?�Ŭ����|�q��9k�����2�~Ak��<�Y5V*-_�St�>H����v��gf���BF�_io���3�
�N�z���g����cr�/��p�;�
-u���o��
B�n���ָ0���hv�����j�H&y	���ˏHs�'��u�)��-��.�^*�R�񿂙
��G��;6�:�Bm_Y�q|���ŐI��a����+2yy� ]�R:\�-�g�d���&��L(�{e�!�]謩9iO��]0~��B����*��Nݤ[��;��}�Sm`Υ����L��=��6���`@䍱h���2��h+p#Y�?J>�r�z(?��+�n�QJ��b��L�KAs�w�̙��N�r,�)Ʋ֬���'Wlz��se���8s�j�%�x���h���
#��o ��L��:���b�5x�]b&AhW���C��g�E�.=ׁmѕ<(%��ȶ�QSE��:�!���Ըv����>	�)�=b}��@R5�uƇ�}W�L�(>�">��Y�3nh����"|��c�i._��XC"�ܛjDtP!��綏��	>�E�C|�9.�=G�W�ТI|�Nt�z`��
J2�JS�����y��� fg��p_d����p�㹻s��)�[g��7��m���S�L�a�)6�(ק"�nu­Œ����;�fu���>�a%DSS�'� 9�9��E�4���gΘ�3��1�s^<c��r������>����#�j���zY�i�jN�~0h<��C�/7��Pa+j�y6�~����f�F�o!�����Іe����³��j�~BK8�J�X�I�C ���đZ� I��}D�Z�^��xC� ��ù��շf�J14�Ϊ�2�%ߡR�qC�S�|�}�"A>�ZG<�~i��i[�ӝOH��ۥ{+�*c!�R�ؿh\�:a-�����"�I#�7�r]o,��v��
/�]�ͥKWtн�CuM�:�F&Wv=�=FSƓ&�A�*���^̾un2?��2Ki ��T.	�\k�?d���"0�Cv7������y>�J�1?�ϻ��X�vs������i@�Tu���Y%Z�~��e�T�W�eR'�A6�]�Λ>�I��uw!x��F��$N��_N�Rpc�>��H,�`V��!�4�{��}��P� ��K_6�\��!k���J\���<XE�K��t�n�M��/{�D$f�BE�@3fi�������bb���{����巉ީVx����ʰ�����k/4��C0o��8�D+Рx�ZI�Q���v�t���9Q�hշJ�&���P��o*�ԧ��R��2�	���Q�.�ɗ�����&)�|SU/��<	/�fs��m�
E��0
��%}�jZ�w�SEl[?�({s���O\����f�N𧖤"�����E������R��@��~������.1"��n�_t-k����"���ǡ4�#k��]�U������Px5�����?��N>����Qڐ�Á�J�7�4~BQ3&ӻ������r��s��	�Lɦ��|��^����j�j᛻'��2��2�}�����E���eY�R�?�=��2�����
�'������k	:e'o��{�AH�DjQ�jAV:�u&��4/���J����^��4m�e+�̢$�xii<���%��B�_
�(`�<�/��Q���B��d������Atg?����J��͒�y+�ҵ3 ���ǽݼ^���J��˅��#Q^[��9��p�fj$�o���"���;�}�R �:
�h` ��!�e���#�#�@J������a��Z#�����lPWC
� �'�����*��0zv�>�r��x�]K��3Dٺ��V���͇�ܓO���:ݗ%��j�@���|5�oo�e�p�ZI{������Y�ٲ��V�������
X$9���SD>Aji����ۏc�gyo��Y�LPGt���މ��Ɲ�yc� 'B��XNM�[T�G:P��Q�v�C������]�P�i}vd�X
_C����d�J�X���$�Ny�j��:S<��e��G���z� �pmm�Q�V$;݇6���$#����hA{��$⇐`�/wB�r�rE)����ǝ��Qzp��d�x<��Lra�T����WU���1���]0�vb��?4h��}1�{��?Vo�a�Oj��� =�Z��$N�����x�������(�)���h����6��x�$H�f&�/^aØ���!9"E�tŪ�U����}�nhIBu��<p%���=��]`M��u�e��*�DH����.qԷ����@���}+����:�&����D'�������e�Ó2!f�V�{}Y��6�l�
^�	�;X����H��;z��J_=�MAL1�<5=PJ�
�O��� �X��i���%�������e����� �T��9��iEl�ݒ��X|��6�B��)�{���k�!�����-�4����d;�T�-]L%�j��kgGf-J����O�{�@`u�Fo�8b��HF�c������jH4�s�,��yR\��לg�]|Q�F���z��u-��&%ߘc�_Z��!���L:��%�j�\��?eG��>���R;[n0��ˎiϔ�ba�T�1���G��$�wH(���.	��(/Ő�v��8����@|g�Nv�wh�����1����%a��[�؀����5r{W��Ջ�_�e�:�j���;����.Cj/��%So�zF��]���J��� S&I�������������e&p_��ζ	:���x�+��-i�9GrL�M���\[��1��nB�璇w�������?"���r*>N���?{�:6�{��g��CD�İ�?Á�AWe7�1� ���+�g�jk�Q� ��8:�������^X,0}r��Q�Q��ͧQ7^�.*�wFp�@����4�-�g��O�v;�����@������N�DuU�@���+��-~y
D�rZ�
�
�b� �k����~��o����������Q�z~�q�<W�.-���(�� �C��zWh�ʛ-�/'��
�@�|�$t�Zi�;Y	�p2�M??�T�܅���I3�X�Umg/�����p��H~�=��C�2��/b������+]��W�7�m��Z&�<�H��h�C�cu|��o]�K\lP�6�05��A�ׇ��N��!\�E�%�@?�h�� �a*�h�����RI��Lw�	��=0p��j�34�T.A!�S�L$_���<'M�y����3���@�F�����8�HD�H��������;��W�)�W����Pe�y j���a��M�4�YlcS��I �#h�)��E��"Ս�G)���x�*����mh��GI)�Z7���o���(9�WS|m|�pK?;��RzZ9�X�f�HS�+�#S/��4��o��P�f�~��9���>ˁ^x�_!���ܜ�˯D���8�:�`\����N"N�B����z�m�W�Ӳ�G�\��S����Fi��_�Q�7S�I��*��;�L'����/ @��U+2�D�R)l`��puh�85K?(���b��1��C�>��F�	n��wӵ�>�Ç�ҁ5א,�T�d"���'�a���+b�![�6!/�	v~]M�y	Dw��V�2bM��'�RG�Vk�G��ǩb>����ؙQ8�%��>Z4ܧ�'��,��s�B|Oɀ��cȽv��iWy��;o(s�1�t��!����n4b�RJ�w{t���Rs"��e��@�����!��S{Mti�N�(��]����ゕ�t�F$�kF �KN�u��m���ϳ����+,�Aڂ�ᡍ`eJP~tK��I�lӀM�}� )�SM����v/�k�R#%�I���U�(Ȓ��������z�J�!��Jj����%F�K|��5�)=�|�h��e�-^�G`��Me/g_g��!vCG#��z���Ȼ����s����c�&(G*uhu`B� ��m�� 	�c�eѫ3uV�R��~9
���)������J'X�����G$I��9�;�'�R1P���-7�D�5��һ�/mq-��!�H_�k� mu	]�_~қ�<�4�ϣ�B���M�(��I����'p���H�{8����( a��z�iݠ�ԝ��i�����k��f��������A����Eaa��BgI)t�UL>�n#��6""�?A�Sy"��^�b�Y�I|ʍ��
����` �A��:��zLx���V!s���<�	S�*\{?�!&����_8Ov���l'�m%�?����;s����Hl����k+���$��x8��㜵-�Ӎ��~<����O�tO�C���ˋ�!)�5H�g��67�Uݕ�6�{�,���MY�]k��֑X�"�����w�ׂ}D\3�J��#��
F� ů����	�W0�B��6U�S�c[��j[�%�R�f�I+�".X"� N�����Kub��c���X[�����z����ICf���0㕙���*f��pz��Ӯ��t�.\���Ғ���P{I˱����^�YӸ4ͯ����q_Cbc�<�b��I3
��w��?�w�n�Q��\�����B^�GQ��AE?���p~��Z�q���2�Q�Ԏ���i�;��LK8�;d�Z�=�Sq�b@H��:��A!�3��z�Kg�������P'�lRD(VF�o�\�_�5�<����@<�׌�錦�M��>Q*��h1�����T��6N����Y�/C]�����oք\�أ�!�&��\�D�S(�m����N==�]�L���C?�K9�L�<0/n�&�0O<(N���{O�?�\��MƎ۝�0��f�cb�a3ر �&��^V)�o��1f�	*h2��2x�1��:�o>�;=�c��juL����E~[!:z����d�KF��>@�LLEw�*-��)7W�J�9��q��p��U�1Ȣs�	�v%a�Xt_rꙸ��F3��O�"��?��KC�@�F&+��
��v.t����ç�*n�q;�V�����U&N�������T\6cҵ�9�Ъ%�|t�Y���q9@@XEiK�sZ��F�z�O<f5�ҧ��c��r�>��l���8ى��D�X�;�O1J�;��o�VL�\~3C��F���y;ۯ��������ڪm�k������?\��VH��c63gj�޺z�\�4\�J��4YY�)�Jw�r{��8�l��
��G۶�E�����\�_���.~sѓ���8?����%�ɀ��W��� _
�s��.n���VAA�!m��Lb:9xR;x�z��T���%���W�6,�+l��� ��
�y�g"�����T��ѱ�S��:����OUl��
������E���c��6�&�Ε��a	#s��H�O�~dL�r�|�@���Y�S���[:qa���o�E�u��ͳ:R��((�?��G��:`A�ED��D_��R�:�s�A��d �7���U	8��,�K����j(Int�.i�o�J���P�!�ʦ��U������wb�p�k�������D�+�����*�1���ZN�8k?j�Z�RY�'��х�۶ݵ�j|Ej����l�'��yD֦'���R2�jԟ�@��I�i��Q��xK�بPC�4D���V��]W�\���O(�f1���$[{���\�������B�o�o��5�����d4N�i�5�[l5G[w}��?�TOX�6��}ɽ�jT��"S��%�T�V_���f#}��9^o�Y�n����������L@����<I-*�o�ݑ��@�g��Q,�B��ܬ%X����aҩ^Zj��E���c�du��[��
���.������j%�U�zg	���J��Eݎ������1�>�^7��w�K��}�h�wȮyg����r�ދq!�֚!�v�"�RT�<5���6|�D7�ҡ���)Y~+B;�'azWoXڡ�6�֕��;���-�#H?���YZ���UR��]H� ��D��o�Lc���3i�J��R{h��S��6q���P��a��u�`���u�:�����׶nߵ��|�>��d�-��9,�&����$��n����j�h�^��\ۙ�I{�M`���Xv����!�	o?8&y|���G���p�"ח�RI�n# �ֹD�����O(B���ʌ�nUE�����e����y���{�}י�K��3�����Tm�R �ݧe>�2z���~�G�M������)�^��w��es:*HlJ5$o�z�C�fG��$��]����Di��k��7M�'�S5�e6o�^��j��0�v(��_���T�רz����r��V��=<9��GC �5@��d,������ܻ��Q���ybp��#����/E@�н��&Ӊ���lp�&�`?z�/XU�VE��R&��E�.��f'M�[GBu��c��n����mm���U1^��Xvg�O'�F�rc��*�3�W`�-�饞汼ZjL�3����'�ʭ��87!s�N�K��M˵_�`<�sú����8�w:��lS��#��A�`\�F@�ڞ����am�A��GX�P/���Y�Hͦ�K.�%�h�i���,w�KY3J���-~�"����h�1�Ŗa�k�k�Vq9�7��u=	�ܑR���?6\���*:�S|����G`�iڻ�>!>�{Av-C�J[S��k,�����F"Hh������=��8�@�J�;5�%*��0�1<k5���2�y��v�<d�zj<�͇p4t���!����G��u�_U�O4S��FX�^���|�%�W�|�Gr�9U�g�7�)$Nl�mMd�/�En�ʅ�=h��=�*��uGowN���~�k����-�'�ڸ�DM6F�_�b�wp��ͧ��N���(�Ŕz��&���N�>A��ԟ����w@IY�~���Uo�d�$�Q�O�Tm������9 Hy';� 8JY���I�J��{Aʱ)���ȗ�[��[�w�0P�����,
d�y�z|0�}@��Mb)���/�6 ?���,�Au,�D��,���9ȓ�WE�2M4�R*7���F��~�IF��0v�9Zh�ZLv�3�O�}4�Ϝ�=��Q�aDm�r�. ��P���%���R�������Qݡ0'����E;c�E�����y;���>̦'��z�UD�懬M}��۟���1�pa{�,y4�'�O�}'���,l�6,zف����wؿ���;Dx�vɳ���눵�ᙄ1�=�tMFq�ɺ��]���J¡����s2�3��۰����S�V�fw�R(�H���/:n�a! g(b"�g����3��M�C�;|,[�"cu������Բ˧z��jd��w ���V�t�ϭ�8�F*f��1T�M�ď��Í`�l}o��34�tL��C��Ap���w���;��վ�*�o!�th����V}�Ȋ��j\�B��Lf4X�a�ƝM������ጇ��Z��b�����@^tt��ۣ�&B��>��oP>��_N��y75��sW����[��Q�b}s�4��(/����4���t�cq�F:��0���f ����q'�_�}�
���s	��5şL(D痡�<�z�4ofK� q�xn#��wJ���7=$W��h�U��7�@6QSP\hXV�!϶���{�1fwX�Ɗ����Yh�b�����r�m�Un<�[�P�G�~����Un�e�P�e��SE��-X�U��|��c�����&t���'��@��FkS,�/���|��|������ʉ���(yV���	tk��G$����[_؃��?��1�/�^#'7��J8 �PVKw1+�0��-r��]]g�$�6�g�wOҷbv>u�9�� i1"+����F���@���,-��Z���(��.�M0>�)�݊��l����o�$�O�}���Pg����G1��������KA�vv��K�z��� �Gh���͋sy�I�x҆h�Kx�#1&����^Q��N]j�e��z�0�35~p��=�ʮ�/Ed�����u���_��)������Th���X#����Ď
|��R��\��?u��Ư��UUxdW儳6.I;R~Iȧ*kJvnC��%lw9+�G'� �XQ6F ����5ӘخK�^
�-�!�Do��k cŷ����H�ESa��9gp�}���H¹ �iM��5h�
�s�m7��4*�.�7�s��Ξ�|��U�s%��?���.{mADP�w��(�
��<7�l޸��ѯ�X��i�(8�,*�gy�η��X�iw��T��1 4rC���G�?�� `)K\����?t�2޶�7�V�����>z��Af|�EF���׋�x�kh�DI�P���m�z�����kT�D�I�wg�}$��Ɂ��Zc�@�9��.@\����R�Q�	B|�~il>�K���� o�"����9�m�@4x&Xu�K|*��䃔xȃ��06t�cr�u�(���uA(I�\a��k{=f�G�g�0�N�XXp�ޠD��i��K�����Fn�v���:}�y`��>E�~B>�
�7�@����9��������f��+>��7!���!i!�]w��~� ��@��$��Ή����F��$��t��Z���ϕ�@��RT��8Dj��꪿�b������A�fbP�=�����/���եC�5��7�A�]Ѝ�Ω�a���{�m�-�� ��W@SsA�=.椅>�R��e Ӻrm��8dV��-��2[/�P�ɏ�o،5u��Y�=3
fr������-<�T�x�&7�( |b� =�&�u)�+�玃2}���-� �=��;�|�zk
QV�L;f���S��@2~���r��=��2�꠆�"+�t�B����\mf��Q�&�I@�Jst�hM��5CV�b��`��@���hN�X�K�y��c9���ֽ�;�re�X�H�R��ɸ��B4�P���ە��'Nw���ߣ1tdh��_)��y>]l':�N���C:�&[i>�-G"��558pׅ_��+���G��qT1e�p�nWm��v�(׌f�$#Ѯ�(i>9����7oAC0Y�!N�t�ŀHeB��v��_�rn%-���8�����u��F؉�� �v��Vg_<w���n��P}��F��;� n�P�<y�_4	;�G�\���-�-�B� �L��N�)Sy��ۙ8í����{���T�-���ҍ"��J��B�tqWrw~������0���Y�h��C��4�oh�i��c*[1[���P��-�YN�<��JH��Yy�6��p($�xaTAP���mO��d��0; W�g�
���ǺFGTd�w��� ������2�������pf+S�̝?<)[���;y܃l���]�s�l�=����G
i�3���Oκۈ}]E�'�a��h�ⱴ*� ���2��\f]QRq �[&��3W_�?�i���.z��<u�X���k}	���e��ͻ3M��Ң���� ��8G�ƶ��W���ٻ�B�;2@� ���)%W=�O�����@$��~2����D-66~7����EK�/��	?'�1�&���r4�ܝ�lb��+���;&c�M�,٘��cT���~,�<:�sZA�W����4�sg~ȅ���(�|�����kT�LӔ�μ��A���CO���b��"$��@��4�϶R��s#�k/�0G�Q02�n�����x|��"����ض���f�֘x�$��G����u}0^c���7L��-���$�u�D�Ʌ*h��{��~�� �#�Av_�$BZ����*�B�^5J��K|�2��."�2k#�i�!�(��<. �YQ�<y�OTG�g0<�3=��\��v���֤Џ���j7�S��O���!��̀�jT~��_#���Π�Y�na�[D0P��"�e@Ú�#4_2c[ ��f��V3���<��ҴQ9)����|��S!���B���stL��74t���Ç̍t�ʸ��� 80�'&�˹��z,Bԁ�4%<" C�-�Dܭl��a\-���9^��
�NXP(?�L��}��}����d�6�H����Df��QƗ�ʸ�o��[��8�`���ݒ:�/Xz4�(2$m�&��NaL�K����7��`�کn{�U�E��I�H9����t�hN�p��C�Ӈk�!�Y�"j�|a�~��r�|'-�%���pS^���=Im�B����`RX;י�#	~��Q����.�����:���JfE�ֱ���<?�����/��py}�RR>G����AeM�ڵ���"v߬�.�s�>��9��F�%t�(9�81�����;.J��O&�V���ZL�_l;j��Tr<}�z�x�� ��N���!��i��v��ѐ���?����8������៽��~�O,�����Ъg���v`�&��Ku(;8���	e���Iǚ����&���������r�����T	H8;gu�M�6�W�Ҍr��t a�y΍UN��c��Q���~5D>o��a.�3>B�Az+����+�5^n=q�B���ؿo��V���e�]<�gu��j��=ވ�N!&�D:��2��o~���� ���	eSKא��\��J!�.{���<6�����-�̔"H�(�f������gS�.��^����N�g�兝����q�h��j���Z,��!k���U�f_k��^��.Fh��u�vsKlq>���)i��wH���&ĸ�!���(�S0�3[F�j�(�;�"��7���2�?m�2���\Vw��Y��;[��+�H��[�{)�u���x��h`1�c����N����$.�G�~�W��m?=^����]��=0^�ES2^�� �� ��]MM�+��������r�+�}���*9�5�]�O��r\��L6�����آG�o^�ǖө���p�\��/�����쀙3=w��_��}���Z{��W�"m'fԉE��]3�ژf �2�6�u�}Տ�y�i2��ge�$�Z�H�"#��Q)�����d�6>�MB��T��D�4�/���$b�@�Ѵ.��	~��\Zv"����~�Ҥ[aѳ݂�TD���L�a�hz�fr58ʇ+Ǟ�p���)Ĉ7����j'Q�& ����0�z�?�Č#��A����7�u)���oa_�����P�W��)8kw�b^NZB	o+v͹ǝ��p�9���'k���A"D&��}S��>�_+��\
��}���t1��=�1x�j�5Po�_��S���̔!�Xh��|/�w8�T�~���5�R�J��?(���Ĥ��v(S9�M	��o9gA%�T,Ȳr^�ZgC��b��Z\ ���S.!���;W� ��5e�Z���>��>���r��i0S4���c����3Tq8�~��$���O�أ��//�dEn��a���S�=�p���[H+r�XƳ�F~X$���(p˺�v�i�"J����R н��T4V2�ZO�{}Y� �+ )w�^�ؑxϙ��mc�*�>{�1^ii��7$F�,R�7�XƄ=�b��쵫Y��D��;U�-E�a3��}��'�/xR�P�@�Uo&ovlfN��2�~Itn�ޝā<�%|,�1X���l�$͛]���@l�0B�i��n�+AZR�-�6؜���UO��ӭq �_o;�����?�_��"�Lh^"ei`���3��R��F)�VT'�C�8HY��Q��T8ד3V�������%��vN��wM�v�
Fh��HQ�����@�����s,�r�e����Jv�c���8��
篦�l��W��2��){!�1����,�����N�w(^��OJ�-1uR�6�r���X��6�}��+&�b��El	�he���3ߖ� �P�.����W�|Gj/+h�l��q���N��x�`i5��F��e�S����4�l�GL�/����2�:ֽY����u��Wf�/�.)W��Yz>��J��2��HBY��a�o�^xB|iGE�U�$P��ȣ=��Q?1�_V_���](O���,�W���i���p/5UC>���]
~=)S����.-�҉R�w��/�yPἫ?��)��*�ヷ~��_��Ud���ߴ�m3�Uz.�vs�+�4EF��$"�f�W�g�Z����I{��K^?kb�W�ιz���ϭY}��]<�W`qǊLA�M㆙��g�G��5�hN�e8˰Ӡ��I+���$<Ҁ%����{ו#�~AN0|Ą��b{ܿ�-����!E���?�����uz��_����'��ٻ%��8J�H �>��s{[�̘m\���Ʋ��п((�_Tz�86Ϟc���a�w���N��`P�'�H
���i�o�d��'��ֲC�ˈH����n>���u���B�N��*��>j_,�Z/�K-y�1N,�>-5�0�5Uo��$��ug�G �]�_Yf�p�%%��^���O��iwTtm�\��gT��f�1,����\�>��2��ɭR����]gG]`
��t0r���&5�n*��n٣U��}DY`��8R��"_Cb{e��u�����f���_V~�`L7���.e9J�bS�� k;����#짯��5^3�Hnэ��N���5;|���<�K�<�b��}��kۏ9AG�te�㤯���|�&HL���~������&x�bg��Vڣ�8Ά�W�0\�U�Ԃ�bA�ǰM��>>6�mi~���67�� �i�v�cR��/���<c6M���0h|�� ?�������{��=w�U�Vz}�8t35�m�ܺ!�ٜ .Zc���MZ��MO�9��S�q�+瀇5������գ0lo���Y��S-����!rdN�^���]d(�;���~��Il�e]�d�daTw6��C4Y��\�u��E!���Czo�Ь� ���D����j��A^�=3��-˥"��C��Z}���`oj0�0�e�FA
V�AL���׬���tnL9�A��P�ج�x��T�%�M�����_�2ݻ98ss^/������L	à�r�9�_�x'���;ڃ�0\1,�z��1����[�|>����7	�fn��C��Oo�Y���(^����X�I�<��C�b=�T��]�<�]&�B�3�V��T�2.��gf)!X���6I>1A�����X_���1���)A�H6��i���Yi�W���g�o�4 17�/-�B�����%�=�%�`��>�kg�k}r�A��,|K�B�S^�C�����_t����r�o��1��7��&��vW�y3��pA/��J���z������P��ʨ����l/�� ��z���gx�j��ۼxj��p��rT* �u�!����P��ե�l/?���o��^�m�X�ͣ�^����Q^*|BR@)]�����v�O1�)��Կ��L�-�)m��;<��]<��U���0����>�J�����p���4X�I`z(k�\9䊍7.&�ށh��K'ImKS�۲]��4�yK��G�i�9#�)��:eG�� i?LEb�8��wbE�m_� Kt!u�4�}�(h��$B��z��z5���O��(�f�H�Q���~[yG+��#�u]�/�6 ��,j��r%��C�*�|5On�m�ۓ�
& ��wHu����ϙV��MC~:/�ܩ{������Εbd��bo�~���Z��cн�]��4dɐ����󍇗����6_��D���tx';3���F��J��	�C�B�k�:�Ƞ�����;q���k�.a8F+�qr�	N2U�^.��U��J�Twf��z����^j��n&@_�?��h<�q�;�7�9B�	Q�h���4�Wo3�XD��� �l�#� 4�c�M�����~ )�f�Y"�`	�}��M���ŕ��<�	92ƮəV�O���Q�TJўc����#��Z2� ��i����\}��Um���e��:���~&�f��Ő��c�fોL��^w��I~�S0"���{����Pp���%�+���cti#�
,������S�`�/�N4�3�Hr|��L���Â�Hҷ������MA	J3V��(���6u�HU� H� 
�M��z�AT`�Z��DaR�32?�?�lv� �n]��C%0�e~_��c�.��='ec��{g���\6�|�Iu^��]:�f|�a������Xm�+G�q��]���2\-ݜi���j�t��ȴgkBz&e�T̼���c���~z6~�0��������r����<{���vs'� �V�02 �K�
��Q�p��m���L����L���Sfl.��x*���	���te3�"M���?b�$#�(��ۍ�����[�@9�ޓ`���ޠU��I��dh���|L�f[���đ
+��>\��ìx+^��@�����s�Y=��՟��(�9}ڛ�܃���G��x6��L�a2�j��*+!<����w%�m��'�E��>!�����;o�\U��VDʆ8@z��7�KKtO�뜤g��Ydq
��4�Kt>�cj�9��w5�eE�&���;��Cv�咅�)Qkucy��;jAEھ�\�]�	�3�w�1߭�����t�@�2F�9��{��_qմ��ԲlE������"�>]}���
Q�V�Rs֒��t��z̏}�"euS��s����A��h���dw]�V��5}|��P$1۾��RV���B$/ ��7�#�w��}�4O���oR��L6�X�E�C�'s�C�̝pMM0v����N<��Tc����3����)�A���>�Q������hَ���Z�T���yi��fAO���Г����:hO�򥻭N�w`�R�{�(K����}�c���ZV?��S�nZ���(_M,o/�v�����%��` ȴQ���4���P0�����Vo	RN8��:�����!4�Yd�f?M�I˽�J?膜9�1����]�y�{.y6������H+�X3�����k��W�1���"���@ ��������G�
�����FL���8>�5�`%4���`��OTD�h�%�D�۱�%���Ds�3e�S5�����R�0Wɲ�AEch<����F<��f��y˭$����.dl�DU���}����$�����|�ZQƀ.1j�?��.Oc��l�$�����JLF�������S��?ž�`���g�29�h̑�vߊ���uU���XU�U�(g<�
�"tz~}�3���lܩ���w)\�GФR8�YC䁺�������'���1��M`�dX#�L& �7�bo��
���$T��.#�0P�|Cň���Sw�'�hK��U����K�M��t��'(�h ����h�J�-�����0����{:��`�3��Q``�-�)U�����$��S��oeC�C���t�Κ]u�z�����G@�tz镕ûpgT��o����>C�(]o�-���J�c�β	0*bUx� x���R�t�^p�+��:���r��n
֌��A1�KjuscU��p��{�8-�'�zC)�f���] |Hi�!6Y,uK�^��N��XX�d�OdktSOsB�@6��1�@�um#������K�o%�\�Y�".��$%�ܱ�;�W���=vY1�Q�{�B���������$zPI/���`ͩr�,8���cq�3U� ��<*
�K�� �U�:��!�!#־�"9����s�~�22F�
$�h�8�#;1-^�AH�"����� {��m��r ��\��ߴ]�y`v�f}���tx�叡r���"뾍/���;�R�j-�`0������2�v�*�qZ��?�M��M��!�Z���M�.<v?��\�}q��2H��<L	�!�t�)���?q*�y��E��xh�Ź-2�K�=��/�� $6�4�����LT��j6��Ȭ�8��Z�;��;��uS�_�����)Y�흗�}�;lrb!�=V$��;a[v�y�d���:!]���	4M��|Ƽ���-����K��)�,W��! S�M:�77�~�_�DMJbt����@�40��aV ��Z������pO%�п)Z��|�y��p�-GɅn�GB+�h1�;YmLE����Ŋf���.s'�����C=��J^*G,�?�9�x���GL}�\>�f�7�9��Ǎ;���h�V�z�{�ƕ��D���G9<���?>XM�)�#��m�x~5���U����F�������NBD���K%vn��l�h��63�R��Ył�|
Z�8)�<]C��i�'����`=x���ܘ��w��a@��&z����^K�''}��?���#�#����J�l�y���|"L�莜�Ý�/�W������,N�CΑ�? 4%wW�T�a�}�ވ
-mմ�q�������ȴ�B�~Q�ֲ���ʠKJ�D9�Q�.Y�çɍ� 1�pԂѮ͸2,mnJY�p�v_���"�/%zR���4�Ȯ��)�nB�]�m6A��h����7��7x��Z<��Ե巿L5p��*��)7O~,[�0��!B"���3	�TnC�dL�J+?�s"�/9l�P�$�y ;[�E���[�K�g����H���b�GR���
�f'�3�|m�+���5a�K�PЄH6hR����bRfG�������ղe�����C\�'��7C$��+K���I�ীC�AZ-���c8F�9�)3&!�:��O{ƄEf���j����ډ��ds���i����1g���� 7?����qe��L��'�ʲ�ۨ���ѷ"a '�V����� �G�L�.B^��VA2wj����ƽc�@�MA�K�~%v=%��6X�F��Ήtp&N��fĈ�!
�u���6��h�4qK��^8�<��q9/ß8���nA��LcB%��A��L i����AAߓ`Դ���	�Co 4�i�uI�\�ؒ�<��7�y0�\ݎ��6]Iѝ�:$��p���N�&���¿�A�ܪ몆�T���o�`��*�{�L�mS/�p5A*0s�my�n�-�U�
�G��\2@.I˜)zS���u�ϫi�g�Y]()��˜eO�~��� "�����Y	�_x�6��-&����s��@"5k�U�b�q���9�[FZ"!�1��h� �B������V�e�?G��� 㙊M�$�a�,����V0D�+�м^���fa��+�|D��Z��_�S�Ô'�UM���0W$)QBqB�-��{�Z��_Ut����'��]��`青Y�߈���F�Xܶ�?��i.���Ρ����<���G�B�t Oh�1)�7�,�%e\�)Ҕ���#�:��'h�f��\&�A���ٰ��xë�1��d�O�?�<=�=�'�'��0�4�`V�`��H6I� �VB�m��)�7������'�f�|̺���3��/H�eٳ��&v������{�e�v�#U��Uȍ۟n�+p�����L�6`�Nwվ2&j0�O����'d�û]]�����e����H���u��G�~�n��L`	LI�Mb!wlB��4U߉=���`�Kd�J�;'Z�v8��ʤ=I �/��(g=��;E�}n-~.��U�b�(K<Z~��&����KO����5ͥ��S@8T������MF}'*;9y	�9�/N4��d<m�
ă6Κ_�7���� ֆw`��,�-B[b�TZz�N�v�Ocϩ @����N>FECs+��#ª��t�!^d�E [�L�r����<��D|����Dƻ��;7FxNd���ᚪ}�f��	5e`Ү�?�~L0g8C�j��q�F�a��&�R`��
(�j�QB�.��,�����3Hy*�~c��,�<�ҥ��/�/��z"͊� ����]�=i����Uoh{���2��̕��P�E�7��#�����_���<p�2�Jg�������;�2F�s_�h&T�������i��=S�wL⵴�Tץ���9�K�쑰)��Fr������f^Jh�IB��Y���8�=�U��=�{�_UXm\��3��BS���R�|�fGʤ[���j���c�F@��L�V�y�z��:Fn�L�G�4��S��4#�j�_-�q^��x�(�҈<q�������3�8`:���c�������Y�M�]���7X��µ�%BU���'�#Њ�](��m�Ţ�v����B>�r�d��j2��a�D��@f5얃�Y%���P�u괸m�[h��<���y;�G����Z�z8x���|:��:�T����ta�F%)�/b���bP'��A�'�(���lS������Xy���I�
�"�m��C�\��&���	2�"�SmT���+K*�������@1�jȅW�;><��QWDs ����s�L
�3��4(0�0%�G �_�N ���4�!n�ݵ�=���ߜ�[3֖�M�K�c���lvse�>��
��tH���֑�@��K�P�?yK�\r�ka�옂�Q�ȸy��=�v'��BK���.�Ȉ�*����s�SȂ��gz/Q8�#�R�"�{�峟,r�@?��v�M̟���@�	h�3�qT$��{g��E&a9%��`���Hڗ�-G%G�:���O��c�2�g)@�3bMt2DtB��7�$���D5�L'��T"b��r�z��#�d<FZ�WM�Ri��~�9\�V#(�� �����
l��* P�Ͼm�J����Tp�~nT�1�.<g�CGB������6B�Pa)k5:�9���5�Y��u��`e}�S��i,MOx}��H����ƒ�n7��5�z�w=�3�0��$��y���ֱU���L|b$7�[$S��\�g�hE�E7PpF�U8<b�D���R���� ��\=9=;������j �tNMV�0��\\uP��RY�Z��`h����0-��bh�T�%�Gsh��b�&mm�US��Ԓ��},u6MލW~lFj�c]��h9��(�Ci{�&��1|�2$IU��ק�[O�z���^v��E����ٰ�K�պ��ɗ6���G�>;Ґ�7;�Y/�X�:[�� ��W�K2�|F���8��ݾѪ��K�6v_m79�3R�gB%$/��a�:"ٺ�O$�pf}(�L�^4+��CT.��D�i��y��8`L�)�*V��)��+yw��`�c���[�*�QW��ZJZ�b���f���x��Z��Emظ2߯xi�S��K��n�C�e��9z�{�Y������G�Z�������Os&����ۀ�E`d���[�s�ͱ,N�")EƜf�E�����;����*3�6/�0<M��͈̓�d�M퓧��#��	#�O�j�ƆLd�b:3��7�KW���'O~�G�A�����Wu��L����pZ�v��Rc��J>C��>`����D�����m��P��@,���!�]���7���*-�Y�Zv�'��"�5��ꅭ\�!ҁ(��I��3�r��� ��kA�z��%W�^z��;� pnA�-}���y#鯑S�4����6cE�g�ɗ�w��� ��!�63 `�?9�\mŰ�;^�Q�i@Jv�躹	^�2&v.���@g�|	��Wg.��l=�Zޏ %�r�E�"��N�>ŭsK��ƕ�q�S3���|�$)����"O�Rs�2Bb!�N��B��"h�|��l��(c��'&V���E��D�,h�3/��5F�l���������ѹRK^l�u%6�Z�!io2��$h��*�s�����~_V\�2ۮ�͜����H��hQ=��D���1Te��r~�\���c�8\�ux~��%���d���L�͋:ј;\�ɜ�7�`��Y�_N=�W��%����V��h��ř�^z�1ft�b?reŕ�v�-l.84m�S(��'H�=}��.䣸?M��<��J��?I���i��'6� �Ty��G������h%@��ܔ�~��#�E��CӬ��c�(��Ɩ�jNs���`����&�]��~���g	�T�jV�7����Te����.�>k�D�۾9�v�g&�P����V8��:�b�0%�2���}���.c�r�t�����Q�_��~�b8KHi��^�"��X	�F>�t��+�8�t���8��Z�)��[{:�*��E!��;�zOC��?4��Q��"9a�-�����p��1����1Qm���.yf�@�"��pz�^�l���P@�{}�3Ĉ�����uX�d1��my$�L|��Z��4ݵu!��c�K����2$�7����,��l4	��*@7ɞ}�B,�\е�8�*�|`�|.Ǹ����5cG�OT����A��F�UA���,�-G�>O�~:�YN������R5q<r�Hbp˾��5f
�d�>�����*��ö�/���M�Nr$_̕�]�y�k+�f�ZC��?�S�"]�`��k��N���ӹ��"�9��q�Zch�d��#�2Zg�>ȩ�u���"h1C����4�S�oJ���O|�XWߘ��dwǶP�F3'���0�#�¥���*;��G���Cy�=<��1�J�cq������ ;�śJ����z��n�ϓ���:���T\p�WK:x�Ｚ#s���)/���l��"j;������aԖ.�$XJ�Ǣ"�Ӱ��<�,COQR�h�k�;�Dȓ�;�udo� G��N`��-��'���,א< ����	a�G�֛'���?�M!a#���bs�c����g��9��CW�ʫ�ECL��s��l[R_'S1؁ߓMvr�L]<	w6�>���E�MX�vf�/����z�ː���p��ʕۉ�؝�[6f��P�Kz�hqcc������$f!�G(��_$�%�N��o�s�����Ƙ�j��w����E~�Y~ F_TL�L�AJ�-򿬮&{�J���7���{i����|��x�����<�B�4N
��嗲ufz
���W� sM'��%�����!",�ر̒�"	;���6&K����Zv�ܣ#Bc��7\���=Fe&܉��s�8�)��]yS���iCΪ%-��q?[��$��P��ST_Uy�P1.�:I1G[mΜ�Y�����e^������AY�����,0�F���b�¤0T�h�L�Ѿ��.�|�P��Ͳ۔���fR	?�⊳�T��e0��(�A=˵�%���o�Z�4��������F��f4{��O1�f[����U9����jg�����l���"�RU +���6�1�{���Zp�v}z鰩�})e�M�<��h[J�o�q�vPM|o�B�������QS����[s8�W��2����D�r6�G�g>WUu=�m� �,�qRX'̚@�g���&&����þ`i�W.k5������IR.gA���X2.y�cCC]�Y�Ց��!t"��&"�A2�>�����*�n^5n��)Rr47����a8�<]��x��/Iӱ���D�[����2�>���Մ�t�7<k�w�˗d���^$6�b�u���F�&�3S}��FR0c�H� �YP�W��	��[�2�o�p���~I;cV���h��,?�s��?�fʬ�I(<��\�\a֟�)5�dY��J�q1t��>y���"�x�9Bt��Q�=��e��q�F��� ?���`o�B��0��E���˦����!�^G��U�S�&|���g�&��_���Y���D�M�Fц��_�{1��jSH�-oI�f�,���_�ᾷX�1Hl��>����Rl���o�%�*��.�^����No�_l�tҸ���W�}�� /߲��O�G5>K*L�a��k0\���R۾U~զÏ|̯��"�W����N q��R,u|L�+eA��v��Q�Y�l5{3Y�s@�ۛ��u�1����pI�^}�t���\�@��cO�V��;����4�+ ���R�%R�ku�HkU#؍jq���w��7����7�.g�[r����M��/��|�;� w�+��Žc�����I�'?��H�!2�t�n��>Wh0-0&ځ������َ{�]cB��s��y�96�>�$��T�(^���E3��N��������� CW<ǌ�.�E�؃h%�ł�ϯl\8�J�ܑ��=	,��vS�M��N�����{��+� kvJ��ew�P`[�Zr�u�8���1�����(ߚ��P�����F���u�7��_V�s�`ޑZ��WX
�X�2S��A!��=ac��{�]?vPu�g���̟��Jb\����b��{��qZI�1�}��Vy
A������;�`z~�_Kf6�X�N��Cf�L��	~��v�@�`Y]��Wo>�u��mO+�'f�G�W'(�!RaQg+�0�nM��PD}�՚ۋ��x�n�>�14��*�}�~4?�`׫��z.�@\�-�~i+֕1Q�%��~�={@��jM�@����^�p�1��NW6
��W���e|H�p<u�>!%��/�1@?��瞍,�,�[��M��A޾ �l>��{�#cKB���z�#��O=�/�8��e�zvL�`c�P�
<X���K��B�D
ѣ-�I��o@�eM��r�!��BjXv� 1(2 ���o���lԣ�1Rtm����C�S�e;���8�� K"��6p1@¤ ��'�$Az	ҔTK#���Fő�%����S<��"��N�b=ѹ��Ky!�U�tH�K�J�		Ap�K�e�7�h63�8�et`�T�s6���Oh9�x�!�-��vW�U���7-����댦#�@��T�}�p "k��.���\u����uY��GCY]� }9� 8WS�%:/A��`'�Y���'�����|�̀P��_\u+���5i>���&�ý��Nl��0���p��"�����<����-�����4�� ��.�P�"�`�а�ܶ~��Y�X�����ZnO��m�4����|��|Q_z���*�B���ן\��X�$��-.���+���.��f�V���9Qh��~3��&iX0��}�h���|�}<\htl���Ph%����s诌�-�[�\�s�Ї���L�O���w�8�u<�>�V�Z��M�%�9m��쮨��WU�:�B��S�K�I���Y�c""�}����+���mOLK�ۢ�$��f1-�6�:�#v��/�9՛5�404&"�__p�	���:�7�2Q���Z㴋�2%RQGn�,D ��Aj���I�P!�JzmXr�Ž9���u��0�q���䭍��&b����S���7 �y:9V��O��i\���0��6�q�r�C;�z2m�9133�pF�;e[J5�ёF�Zhr��"�ZcmA~�༚�G�l?�a�۰Q��m|�N��S�)����c_�؝0�k�v����u(��M[֗�S	��̈�$r�e��7����>@	��M*i���6���qb�"˼,'�#<��sRx`������jX���t�ʭ�H���X�Q��#��*�eya%r�dS��r�9݉Q�yp�E�������D��҈Ң��W�p��c���Jp�s�]���5�{y���e�m��'JΚ#%
�lx�nћt�<C#.7h���UT�A����4�ˢ­#�Y"1�)Ud�c,,�e�O[-[�g��$~m�\Bc.�a[U�{/���O»T�Ab��͒g�R�f䶍T�M�*<Mk2����8���!���y�N��wA�%��S�V^����3e:�2�RU� N:7��]���	��[g���m�9:���_�E�.�?p�v~_����@c�������vA�G����q������D1�f6zA���K,7Π�=#,%p.���^�F��N�b?-p�i5*:kD�)��2���β��bI-0i.C�Wչb�C>�MX��N�����|���J7n�M�9���MQ�,�kV�A����d��ړ� 9���s���M�ry�mK\��� �M�Ϣ�}�Ş���?�}{���wPGu�@2��v&��0��<{=T�&�Tx�`�o(�T��;hbEd��0���3�F��8�5.��o���q�.�,z��������M0Qq1��Q�HA�-��V�1;z,vl����B��e���F��ǯ���]�����*t���ϖy ���G�X��K�2U#)*G�A}�{	p�TT�S*Fk��z�/7�om)I �J`�����\�ڼ�����! �T\�kX)3�����ҿP���Y� c���j�>�5=~`"A�H�*0��O���m$��J�S��*�@���t�	};,����Sv�C�R_�_9�$Ę.�$~&�d+�ΰK�@n��AP�Ȫ�eR=�F�N\4�-R_����td$��Lz�W�\	����$����'�N�;|�Aa�ke�P�\�z�ݧ���bFӴ%4�R��.$��k(���i��� B���g��ca��d�����ҵ�~���e����2��pSw������,$;#�|��S� R\��d�_�������7&�bݾ:�E�`��A�Q�Mϑk��m���OlS�B/g��>n��m�\�Q���(F��?z� �v���/G~Fsb|�i=x�*[�4۫�۹�D&`��m5���.�B�O�.�����1R.ͧ�_JIfJ5ak��>�qU��{�q�AR,����/��ܰ���R��<^�7�h��g5ǭp�Z�����r�'	$Q*��Ж7��I� �K���i9��F�; >]�%�[澭����8Y�����&W=.�b�3T�`(HgO�DL!���z$ݏ��G�ҙ1���i�U�#���~=jCC�� ��&�U4T�^���L @�}1^��3�io"{�{��8�s�J��{���"�
��Ll�,�3çK_(��^{�e��S���(C�����`\b:�\"�C1S�Ʃ�E�8�u�L*a�5}t8Rɨ2�p>c�Ʀu(�ꊋ���C�,Ȑ_�a�m.9��>(��������L*;��3�mhKz��1("�堫�A	���E��*V�z���c� ���\m��]/i0��O��j�\�!!��ĉ�Ǯ���L���i�-C����=���{a"P9{�=�������f݆�y�g4#�sn�ל���R&݅�d�(�̘��P��8O���P'ơ(�.A�π,���R4[���VYyQI�qoi�t���ux�9Y"�|}[�'"<�k��}M-��a4�����C��x2�o�v�8�V��� ♵�%x��x�'e�NH`H�%O��Y���
��ڛ�����������o2�~�vΟi$�t���#[.;}ɏ�Y̝�����ǎ�¬�{n���
�@W����M��>���U�Ql��8V:>��]�y�jyx����^_��
(,6�Pb�����i��Ze�(���'!�����JOuY�u���MԻ�~"D��T�lNs�6��P�����z��ie���V濕���X�u:b��-�c�='����!d�Vn��(�1�O�7=8aw���h#�\9+&-�ABWqH�8;��ű���ŭ|V�]�H$<�в�[Q e�~�+��ߩ��Lr�%��jB�N�VU;�(���9�#uW��ƿQ!�9���?�L�!yl�ېI�Ō���W�\v��C�
S�@����Bz�u��V�#tܟ���|�'�����5B���V�1}�݄��� ������vԗ���[����c~��q9F�;&h��/A?���3� q����5��ܘT�]���bC�*�k����R�N��T7<��ξ�zD����ؖ���? �2l�+�R'���I�+F�څ�Iu>�-�w����,I{�W��0Zw�8����YEzV�#U5%�
?8����SQ˕�`G��%m��"�ty��dV��v�o�A>�T�ێ���z�[x%H�&�1�w*T�K���x�d�>���f��b���CM��ge�X�hp�C�[+�-��K���hgUVVbhՓ��o�����lS6�dv��C��c�^<�n ��5��(�W�ȝ��A8�T�xW�{dZ+��U��o�m-̉!��s�N�m{� øhj��+5n���'��⤲�x�P�<iP�^��p;���	�H&ǁr:�/c�����ٮP���p�4Q�:\he�-[���#a�Y?4���,K ��ߌ����bb1~>�5�(w�/o�Q��j�Ɵi�Z?�蝻='��}$��<Vgk�v�e�J��x�<3ɧ�>��J2Љ�M�RNY F�T��)eGm��sA �7��՛&)L��-�yfJ'k�UW�5�e|�=�O-숀�.F�Ce� ���/��;+�g�E�$П�0�H{Z�]kD�����@���i�,�Ӭ���YM�>������?=!�������F���9�S��?�(�	�j����V{ɘh�*,-��C��B���?�dt"�Gm����sn_bif��gtfԲ}��w�#�]~^�'wIxJ@;>/N$��=��y�#\�:�6�krJM��5���L�z��A<g��i���Ͻm52��Z�s�V
B�@���HЦ��2��WF�̍���@���n!V�~Q������l{"���o���P:ߘ�[�X�5LL�3YW+&����P7��;BF�퀾���3}��j~�� � ��
����%w6��X��2�7�'�ms8kw�%���oy�����8�z�Ol����g�d�SdX���N��"��g�MЌ~H����D�NQ'���� �%�r����|RXe�Y?�)��Q�t����2Vj[Iy�ϰp@Ϗ"fM\!�V��ӔT� $���\���1���mh�R�>s���Z �Px���j�q! E�\�]��!���;�K/#��e]<6Jx�]�Bk�2��,���� Jّ0�����5:���.���.��y[����pގq*w���>�K���a��b�/���Kk� 	v���^�[�}U�N�f�){��i��!��IO�q�M�t:N�vq�:^�0g@"�È��Lug^� �E��3�1�??|����O�s�K&Z�IF3��:�!�-z�S
Br�	��`��8pu_���S��P�<;���0�D�h�HJD�� !<��V
�(e�\���(B���:Nt8?\�K1)UޫD?�[�m�y��B�B��i�w���!:��V�T5�:�J�3F�D�_��a�P��-�^g�.ɥ��L���T{��D\z�[���6��c�)1���		  �gU�$��A��(0�ɬ0��� �g�i7�L�<��ǽ����]����c���*�#v(�U-\���Z:Y�C m��,�^lo3�.�/+�ӯ:9�T�S� T&�|9�A����3g��KE%2��m�>��H�)7	��A�.���)�)ڞ�}y	��hm)A1�n���|��߈������ ��"��m���Y�p����h�	r5����
;x���p|(���*]dW	bY2
 󐿪>疸�S��"��<�i���V7T��"�e����l����Ǽ���8�ox�W����6��*�ߡ�Qr���Y�{�e�$b,���i�SI^�T��a�cO���ʣ�X�A��%���˴U��=V]C_{��A�,�[�G����^^	2����l�Ž�j�XH���[�p�T��<}��t�	$�~�0@����}z],ki��*��Rn���*σi���z�
���&�6H=�%���2�yEm�L�K���K:���� J"K�܊P���:��ۇo���)����"�}�o�c�/�qLzكW?�5�_4 ��>)!�2f��������&�E���C����}޼�ɡ���'�DA�Ǵ�C ��-"PR���)cr����K��V�Ed��@�$\uvt��M�g��>j:��*�cN�B��h3K�Ғ����`�V��{�9�41�㶉pm�L�]��M��N���a�O�?/�� ���]��92n��\pv��9Ș�j�D��?/Eg����9��պ	��S�֩���|x(Q>��po��×�k�A8*O��y(�׎��idJ��C�R�,:ή�o�د(�d=H��u�8{�M*�9m/ v�f��p(7y����"(����l徫2W��I��2ul@����[rB(�D�$|l��<��{8�l���.���EB��$��DwV�3l�9LLV�;e&A��'��ι�-B9�������I9Y��p!QP�����`�*b&t,=+(��H�=�9P�N�,��6�m�s��*�ѱ����g����{�n�%�m%�U�,+�H�)��K�s+穢wo_�J�h�Ahr��`��b�11
Y�rt������J��c㪡�='���\�o'�v��	�ȷ�:�x����R�W8;�1�ܐ+ڇ�Qc��9�ؖ��.�ڪ��ˉ5��Z�.i^�-C�=��c�2w��]Z�
�-�[_<`]�$M�F*��nkTz5�p�������К��^�+?]�Hv�� �5BR �A��꫄D�|�ҦE%�TT1��h�M`����;t�A��{|���u�3S'Nsŝd�Їt�K!&�M��<sM�J��Ϋ�@�x��$�,�]�=M�.7�JX����fk��r!9���F��L�P�f^:�H�^wtO�V'
V��AQO�nNI	H��OHJ_��[����(�Hn�Y��vT�A��z�����$vc%%a����+J?�9ΞOͲ~`"��4��k^ ���������G+�~͙}��:��禗����}s� �����E����)����6gF�� n���D{����^=8?����$��A�f�<l�R ��lxd�݊���7�P	v� ���:sI��;�Ju�E�>�^�n9��g�!�k�V�[�N�m��r�h��]`o�M��f�s0��k-�Zi6�����C�O;�<��g:���R���_eG�ފT⵰�����56��M?I�co��n�������#ļ�T�������-_�����?���`Բ�7��|���U���u�d�K��
�󒱻�t�>�.߲�	Qe�c�jTC�>��($�qX։r�
ri��#~m�͵\O\<����-���ٸ#DF��'BʸJi�Yz%l��C�
(+����'��2&{醛j��S�����3�85�VC��p!����Y/lF����đ�ҷs���虚�*�H_�~t���\0ǒM���>x�ρ$mx����ɓ�(㡕����]J��(�~�	�	�hp��˼�z�(�d�`��� u�
��7_�Tx&�PwF:s��e�~�r���vv臻Ĳ�ٶ��T;�\}����^2����|�m���Ґ�����\�瘂 Hz�@,�L����#�^�4>q������{���	�K�&�/��{�I �>���c���[A.):Y�	E�Ǜ'$��t�BzMBEP�S}̘(�e�]�Z�B�ū���z:$�C+*�Xmr1��(�ů�A(�8���<�sD���#k������ZRdi`��3���Joy �Y��*�ozI�F�9Jك��5�c����h�7E�ąHn��~D��B�5�n�diaZJ��~���'���kKj�%���,t$E9bw�؏@ʂ�!F�9`�P9:ֵ�(w�h/����^��:��t��?�/͕�I�B r(.TS�=ע��+w͆�$��e���V==��Mڂ¾����7N�hS�?�T?����q�<ꀌ  �{3M9H$L�cNÁk��qtO�V8��-�s��	$��\���V��u����(Pp|5��Hb	����.���1���t�-�xΝ�OEa��*S^��X�6�dA^����0g1'G�����:��)������B�=A�bZ6WK��4��J&��l�QI��j	�1׈i2	��ԣ������M�\��|9G	!�>�;}��H,!�'U��j� ?��e��+��9��:5����ׅ㻽�%8�k�x�s�7�D#�,d�Б1͏ N)j5 �g��[������eU�WR���?�����>b�|�#� n�~������	ԐZ��@胞u�钿KǸ�ض(���|�C���y�m�F��ˬ� #�eg�K?�_�ɳ8>W�m�������C�^��S��/'��7ǐ=+�
�ɿ��>�ꋔ4��%����Pa�b*���b~�Juh�,0���V/������+������� f�,M���aj���3Y+ԧT\�J�$��SE±�����R	���O8�0���Aʾ�bTT�3��r�F�vd){7�3Ym�������vϘ��B���$L%��u&B�Vu{�o-(�{-E��C�mp3��U%vU�w-���+4�&��-0u�&hon�j�=!�>��_A"�U�Od����>G�J�)���<~�����8����{�����4ف�%:������Fg.2��s`��1+�^��v�K+�ǗW+�l�f��6�G���] ���O/O�[�Ko|�w]��
������EYg�'4T>��:Ό8]�M�U�z�W��:������}��~_�����T2�H3 �z擕]�i�}��xW���yPn-�o��`ۅjƩ��C�go���m��|��ikC|�Z-��j��_}�a������d�l���͵N!�K������>`��lI{�t�i���r T$��LI��#{��:uv6�v����b9��&(OM�8�1�Hf�A�.j��p2�A�2d�Q��
�hfi!�t�в�h����]:��?�~���yX͓A�x:���0m|!�9�0���h���05�4��I�lzc[��`k�&���u��?�o��e�H�N2����z�i��7���i�s���?aRM[�)�G0���&�Bc���@�ʨZ�$�M��uK�ؙ�C���E[��ݨYC��}�LH�����UI5�P����Mz5k)����������/�Im�.n֫W��:��@��l���g�S&�(j=P� �l��}ГE�C_ڃ`*�8u�G��5u���Pt*@�wW D#�O�Z��8Z5,�pQBԤ���0�i��4�������l�'��LR�:k^)��ܱ~����ʝ�E�=͵O�~�!:�z,: �O���uKW���)�� �$>��o�����4l퍣����]	��
?��٧&ʃ�Q�&�4mxJ���s���U��`���A�k}��A+��kA��{Zycwc��8&E���u�0졬ڛ;�"��g��,j	b�[?R��$����V��5�H$b��S�����o�}�b��
��~�I1�@LѠ���z̒=#��49�
@��qq�q�L�zD3�����t^��GO�d�^������-Q��	~�#�z�Thg�Nu�����>֮�ȷ�k-���=�W�)~�N�~���g4l|PHi6k����W�..��[q9G�6��?���%�؅9T>Jb Ys�^��n�mh$�U2��QC�a`4C�`,�2p���P4su,KΧ��4����e0���7e��t��,ڭ�7`\K�ᤇ2�c0@�#�W�z��L�p�`P�GH��h[�S�KO$%$��o��^z��+PP��Xk@�����#ቃ���(��D�c��'q��2x7^�V�U�q(���b5åZ����?��0N0��AUv�(�u�o)���dF�3�h���]Uwhwr�}Q8sN�!n���M���>̞4+t1�����nt{O���vJ}=�;�RZ��<��z�b���k{C����y��������h�2(�;C>]9U��
y�u	��w@@t��J��8"}ASG�����\*���&�	\�X�G}�Y\ʺ��h��61˘l.�}�QE�{��a��o��N��an�v�PN���Y�\��ć�,m U�\٨��V�^}:���8�J�ݩr���0S�ԮN&��cK���#��ʋ��(������� �,Q:^��k�.K�k�ב#Η5�Si2�����ᩒ�H!�����Aw28��rfw��h��WY�q����\���n.vp�5�a���PL�i�nO��N��h�ŋa髬����tp+o	{#~�w�@�_�O�߫,Z��w�ѹ��)����j� Ĺ�qv��S/�#�uWF����.G\u�ً|!Sg"�_�����&!�.0LY>$��nT8{{�l ��x�����4D\��)WRe�O"_�,"�nw�%���|��I��E����s����	���֢1���cd����ӓ�X�j6�&�~������h�3�)�t�䩖I�d����i���>��%����k��Fܖw�ܟ�;V;2�7�5��@GY���&$
���� e��n9u�`�
F���-ר_����/��Yo$�a�m���@�����u��>�z���-��S+�~%<��j����*~��^�����a�w�Y LGe�Xv��^�$�"�x�����,s���Ayp�ٛ�מ�n'�h�5#�s����،))��qYO4�}��R��w�����֨a��U���w����I>��Q٫��	�X���DB�O0���&r#��5d������4�S�1���L�Kζ�'���/����;�̠�����S��ɤ�Ŝ���Z^ ��U󑾋�E���X�!�-�Z�7�뺛�fr4�h�o�g�W4�o�	,���9��-3�F��:	O�tw3�>^�T8h�Fl���5�sY�;���qv�Z��u�S8	aE4�V1�8�o�ak3�S�Ԯި���ٶ����E�����}����YiE�GE#�m�i�j ?g����d�d�yėLh��p��0\-}�<�"��Ӛ��W�W��z�᮲~�\��
�
���/��A��<��I�V#CU�2������P\DϼG�'$�5���V�G��4�ɣ���T�B8�c/��F;�xs I��E��̬@���NV��@���Y qw&qx�sB���r��=���m��<ʾ�7�צI����v+��+����Fo-+��@���_��	m(:1�^�y�a�"Qa�=�k����n�@ٮ�i�ּ1�)7�v��{��p[� ����
���w	*��^��
�{����S����OLésjh?�����o9�p-t'�=�ј��1j��3�󰑵T"7���)��W:��r���Y}䳽uv��<��A��႞���m)�O&���ȓڡA�dѲrȥ�P��>�����ޑ@�k�@��{�8���n�E��>WG%���'ʳN�>��)"|���)���$��9x1�pl�WE�>%/�����[�k���ZB�I�W3r�������A��c�'���b����1h�C�����
�.Z����m�b�@��j��օ*�XwT,���i���X}�a���N�z�>���-�R�Iq�Sy���҆��5��xǻ瘍b26�X�ȵxo0"2J_/}�z5��}�}�28_���1F�ņ���u.f�$�J����s9�;����rYv��^�msm�Y�H�*S��.9ep	�K��yFp����:oy�F��fG��;R`��<��D
q]�13A7��x
�5���%�_�q���v�@�����ySs{��Ә��އuq7�jT��2��0�<�푫�S���-@���x0�r÷M=�z}3��!3QU#(;%JcZe����7B瞽"I�m��ƭ�Zё8���ẵ��R򚐾�PE��9q�>%�ܯ�*����/i�:�X?�:��za|N׿��[.T>J
��~3����������>�j����l�Mi�D.%%|>�F�L�ʇ�9'�6��[��S
-~K��O���]x���[u<�^o8C��^� 8��q�,�L{�E�>���oK4�z܉�7�C��?��6M,�5��$5�o�>01V�^C!0�b��K'�J�/{"�z������:^�˓^l���&r��Ϲ�͇
�' ͛�I�s�f2�_��)SFF�gĿd	#�@�~l�F�<r`ߞϿ�������@ K8+�Bƀ�o询���_�>S4��u���"B�N�9���	@`�{�^IS�wb�/�4pcQWP�fɥ��6��y���e��� ��pL��D�nr�K��e�.�e�r�=� �O�LDn�~�M�	�I�����x���������1�p��&�r��wQDPDf�l�k4�ʙJ��>�!��t�Q��H�E�4�|Q�׻�v5�s��3�]���vJ��YӨ@�cG�e����r����f5�-8I��TYr�QN�#i���Y��>�ش�#c�w�X��S�%��(�1��N�:juR�REgt(��e<�Ō
1o��w ��މ���A�1���Оq�$-he��=��������-�n�x	�[-�4��-�i̍	�ҵ�
�@"=��в�t�g�gG�*j�/b�������n�$d(��>Iխ���@�A8���B��Pn���.nH���K)Q��9�f8ְv8"}����Iz����Y9�zw+v6���/�LHe>/|�k.4�S�G҂eUj~�X-�uV��s�ysG� g��x�6Q��$�[�xWf���K�	�͸�n�24���>�	��Q�P3�[!��)���s���ɧd��
r��\d��6�M��$���5m��w��;yF�>��p�x�3!}��x���F�L�'�[F=���t*�k�)�.�Ԗ$�g>Xq�J����*h�̥/h�혉��,E��H_7���c����-'��~i����rJA�1��[���˾p:C�L��R�=����0�1�B��8��Z~�����_�u5�Grᖄ��3�׫��;���ގ�ȧ�4���������,TyF-��î4�B��jx����l�Nl�]{���	* o���?��	�&3�$� e��OyU�Ɣ�Y<���b��8��;�K���ж�+S��Z��i{�p���
��=�d��|�:���������c�@�Y#����}z9��6��c(��m�4I�`�h���!�#FYg�YHϱ�a/���0��i��4]�(��� �pT��b�-LXujy�}F�%1W���v:�}w��/��5\a�~�C�oj�'��v$��A`��",�ks*�N<���\*c7�}
I��FF�ۥ�6SG�A%Y큘�^B��d_�;�������m��;r���I�m,�|_n����tߗX��qM��ԖqU�e}4�O���K�8{#MBvD�d�\��!
%*^�s�T����ȣDe�p����,�i���Vi)�:E8�Yb�k������@vR'�:�� �_����E�Ԅ�$uG��1��C��֚������*P�:���D{Y��8�T5��Ռ���4�Ҫ�V�kHA��c�IsY�@�fC1�1}{z��m�'��).`��'+���em�x;r}����.+�Z���R] �G��!�	sR��H����[,t3�����΋O�Ǳ�?���寅D�j�Z4kۿI>��0x\�$��4��ŵ��OE�h��#��t|)!� �}jq�hv�C�ꪺ�I9�hćT2ؐ!iI�$,��mb2�^\qE�f����'י����3J8���du���i��$��U`]+頂*m���0Ea	��-i��G��	4�0����%~������R�y����-K����s 9�U�'�	[�3�����%9�go��+��֍=�|�ftB�W�� 3�����4+���;�t�vM:)חw@������bȽ/ٸa��ld�V41�a��Vic��9�����vy��(:��<��S	�c��,������ͫT��-j�.1洊�a��(|���]c �����A��9Q���&�����ǔ���l)1D�?�Y��
�෧j��Ե>b&h�p���[)���#����H+���O�?��|���[�������7��ڐ���I�N�fw*�Q\�&�w�1�^���Yb�oؕJ9I�&C����H�!���M���
=n�\���3���P�]�$޲k;�������&c:��\*i����ZBa�rm����1��I�'����5,����{I��	P��QZ�6`�ب5�n�r�* ���;y�N�c�i&�x��I'�%F\�/PN�<T'F�*E�M �@(�u���GTv��&JW��Ӣm�-3��,�	�9rؓ�P�W/�1-}Vd"We�y�q��u�R��BG��w�s�{���!��FX5�A�ƱR?��s����{|OcqشdrP��cF_����ܺ�5�$o���!��$�\|��u�l+T����(���E[�z��G�&��!k�am0d`�����^��jXPc8_Q�]�6V�n5AO����J���8LA��o�5�sWx`��k�:es�o�X��1�2Hi��h'`�X�B�{69�-R�)	X�È�b��7,]��L-������$�G�Vw�)�"�@�5Q��yRm�L�1U�`e�R:Čr�`D�E8�k*l6 N q��q]홿����u
��Ձ�={� _ߠ�}6)SJ�6����~0F�W���N*�a���%Bjf�ta9�n�n��qfλN�W�D.�_i��ƭ�&Z$�G�h�F��k�Gi3���$���.�,��'��)��A\#RtJB�E�pd�U.]jt������pMd����F���/�ߛ��ǲRX�^H���f��2fy+��-]�IDܭXWi�}3��[�tV��e���!�m۔���7���`�"���T��#�^[z����,��>~n:�t�Ta/��G����=�����2T��v��G5/��~��BBV�@�Lԡ��%�Í܊�M�#v	U�7�:я<S,B��|��Ⱦ��\�/��7��x:�P�!���|���wK��RN��~���7��T�6\�n��p0�Z���r��Ag{�2�{*'�	g�C�|��݊��1W\m=�b�<��}a�:^M$�>�Ի��}Fi���}v���m�hN�P�@��*f@�O������CV��ח�I�j�!��ʫ&u#��w��T�@W�p�kqoL(�����5+�BHD.󲊎6J���~��c�9����vF.��{%���jZ��Ო�����<���E���G=��
����7+D���E�9jCB�h���'081�b�4q�!nGH럚�"`g�O����d��{��z����!�,��ӯ�
}>���y%�๚	~������~�q����� ���<��C�ɬ�ko�g���z��.K���Dj(B�M���G�:�y���tR�����ON=&�^MR<�6����nF�� ��Eֿ'���Z��ud�i�U<����K���c��w���a ���4>a��Rl"Tu��EL0n�-	�u׳IV���ۍ�]�{���U��ލ�/AW`���|~�@�����|C���s}G/�G���=�|��A���M�{,����E�)Ko���Vf�+m��\��{�T�o}�E����;n�<8�`l3s�	02�G*�0��SLp����
�����#/��U"���1�
ɏ�Ii8_&��}8Fy %�.�˫��,���o�:�NI�=�~*��ʮA�0�d�p�c����L�^�+���#q{s�J㣢�fͬ�Zm)���7R�I�\Y�D6	X�ӿc�1����ƿ�7��/����uY0a,H��d����d?!�yL�x���,Ey�890Qj�m�S��]�zwR�|b��}��y�@Cg\�Q-��ѵ�:�w�ef�zga�����n��_>Mq9n�CA΃�01�f0�U
�'���tT��(E��w��pj۵A�֪��f(I���;-σs�[s�Ln�/`��x9�oVOd��Y�� š��� _ƅ�<�j�U����(��-�xM��+����M+\Z:�
���L��
̎�wQ5E�i�nT(��4+L�<�+�U�|���ϖ�7b��2lgkov7�j� \%�Г�j�Q3V�O~��
^��j�D���$ek����?D���st�=�[+H)�i��g�a�!�;M�b��d�eyȈ�Zv�^]�"^���jP���1<uLZ����]��{|i�U���U��X.�r2�	������z�F��%���������|���~˱��@(O�iEQ��������-3�U����<'U]��Q�"@*Dme)��m�����@�2
�j؜��Hf�46��*ٯ���	��R�����]��-ˈhc�%�9ud�H���/���RH����ȳ{Wo�(;jS�5È$m/�"� ��fh�b# #Q����%B�.Z����& �ybh��E������ �o�����w��]�_�Z����N���59l͠���J1�R�~w��`9BP�Cp�i%7��p�F���4%e�T I^�*ؐ��1Z��uǯOPF���(v(x�7�J��)���	�5mP� Y�޽�2����óօ�C_x6e#x��/�Oz�r�z�e�ل|)�*/��������TǓ���>��9�_%-	�Κ�?/�%fEd���^����4i�b���,n�Prh��+���]є�M���*�<�,���{�����-p�E·���!8ޚ-�� !���Q�S��8˾��nTS��6�-��pS~�ݲ�ڗ�8b�6 «����l�4�;���^r\��R�i�(����,�/ݣA�z>��4t�P	2�)���mV�W�<�)��Sp��p�A5�{z6Dd�6޴��턟���HݪuM,�wy��������:��;�'�\" /<�Q��޹L;�oP�^���`�״�k	b�r����c�c;�,����e�cE�y�h��◴8z6�W
"�5�����h�����0��s�f�9���er��x��0p�c������l&o�8*�P��t=7�ڑs�$�H����=��sw~���	F۫��a����`K5��!���$�y�z���Ⱥ}�l�:i�����\����'���PA�ݚ�3�r���D������Q��ݤ���ݖ��P��8X	�0��\0DzV"u�/x�&�)����L�n�X'%|�ȁ�f�7G�x�>�׼Oј]���^��g*�����,En�:}}m�� NT��YG�a�V4AF����8��p�#Ė'��C����E�X'����/Y����9Em�bkr,�h�	
�y�J]'Z�y�sٗtk6���O`;w+q�}����ßoT��v���iZ�������O�㞕
@� �U7<�]�E-ՙ況���������E"d��Ny��x�nF�`���!�Z������y�o�`�?r+�K��,Nc��T<��_�M�mdX�30e���$i͐�u��݃*ź�����p�����{I�W�v�.*[�i�NV��rrs��w�R�g��X[�!f�U�@�+�\ ��^����Jߘ%�z��Ll7+�k������w��V<�P�P*K��,4�K������2�)9�7�S`bS6%i�c��ͥa/��WH�t�� /<.�c��G&�{5��Gs���9ʩ*�X�>)�Н0kU���Am�q+����=� ���*�yL�#�Q��*��)���9�ѫ.|��&�nfR�e�SzRpQ�X.m�?]�w��z\k��2�F
8�ϖ�1ŅR�z��^��b��dx�JĤ��8sҭY�������X]U=kS�v���q�.m`8l��,P���G�}}��&ֲ�V:�Iy���s���`	>��`~+�
�t�5avK��	���Yj��י�D{N��׾z�e�g�ܔ9 H�{�ȸ��j�����W�S���c-�9k��u���{j�h�>Ai�I�����JA��\���Ԝd́���]_���7�i��2��(���"Z2�6��e�K=�e{�&6� ���VlL>��UdBϖ��Ͷ������F�m�YE;#��Ը����K�Vˉ� �/�Ci�֩�#����G]�8jߟ�,�,����	�4y?�YA�;h�$1���Z�<yd��B�����l�e�3q&z��1i'M����Fi5m�R�t6s�S�i� ,A*�g�PuvF[�*<%��
��n5��t�A��e	�	���W�� �����p��dN͊�Ce;Y�u�S���[��,� �3:��� ��M7�R�<�I[�-, �- �5Of��o��!o��� 88z��ѺGwUo�^��f����X�NV�M�8���F�.�{�N��5\�Ǐ�IE�sĖµ�E�z����c��
[8�٫��	Z6��y�#\L裮'Wk҇�r�KuN��쮈B������hk4zt�qb@��^��+Ԑ�|�D�D}�����8S!i��W�*����&myl��-�����ia,���D��;� ��Gt��A��K�M��hD��_dL��o�����oPߤ�OQ�j�b[{�X��p�mm:�p�:n���r<-����D�n�����
=���Z�o����7ǘ�Z]&��:99�0
�jr�`��J� �a��qI �8$;���*D�Y�7$�.�A2�>x��ʹ�@dq��f%]5��$}};��بB`��鎁��O?hc`�W�Kސ+�$a���tsY�t���o�z�9�=�%}
B�531#�`ْn�)%���v2a�ś����u�V�\ȕ�&�+v��a��i��.�j�O�cy����mك�3���W��m�6���=�j\Nػ�K.<X�t��<�9ǆ�1<�{��4}�sc�pK��=JEȂ��P�rp�#���Á&ԅ��{�,A����_��L k������0�U��[�Z�(�*z� 5��Qu!��+dЮ�8ͭAabƽ$�2Rw��E����H^4��08�p�)l3�'Y@{�J�6k�&2���F�0#��`t����Wc�c>:�_&�����bQ v�M)�[x��ժ��L��Zl9������6�N���7E�s�x-��l��ޝ˙d��e��Ɯ)/Rs6*�E�2��{�.�	^Τ#�S�f���;�XDa?�W�®^��x��wN���/���z����b�F38���j������Jp�b��.�'��C&���-q]F���scT�ҝ-� �G�7�jͩGY5� �##ˡ\)��1y�R�q���:ǣ�=7�Y�YP��͌9G`��d������Ȋe�x9����}o������C��}���Z��ΫA�����I�]v���l�^w�]�'A��`��Xr�O�%��N_��	P};�T'�j��V��f� �|��R�9�L=Lߚ����m/՞�h��po4fSWZ�<�=�͓ns���f��3�e���Yjmٯ�X��t�c�~�aL'A�S��>(m?w4X⸺��qvA%���H�ڣ�����V��{�&t�nIN���*[�(P(����sHYy���:,z���� ��T���Rx���
�a�J�6+����L�����>F�W��,�=�����ϚR�53���~N���O�1J�VeO'�AD���F\\����8���`�=���D�k�xBn-�&
��v55�J�yZ/;�J �]�ǐC��xݖ��^�v�ꍽ���"V��$p_����U�8����U�#�W"��	�71�ϼ�R˯Eеx	�mH�Jӥ�|B.\9����|̳ehX�BwUzn_&�Sz�0�H�����!*��IW�X��(s����~.��Z����	�O�"@��aI���\��wJ ]�|����M�&l��!kJā.���*1�)�]��z֐��;kL6^�Eb�A�vX��O,}/l-��c$Ң�tv���.�} ,ՃZ�.�o0{t��=�/��F�X'�RK�'g����Y+2�G�-�{�.q���]��S�P�^����Ny�MU��6�.z�J1�%	
���ɿL�`<���/l�l����uX���t�Qj'���/O�F��(��I~ VAwz�?*ם�W���ĕ�tV����Gt����sԄ�R��/�+c�����_a���K�d�[��rA	���m�M�59��d�办��:���]�:6o��;	Y	�u������<��zBl���B)n�No��Ӭ�U�<��NmE�r�X�r�+�<�N�)B|;|/��1��$��r|iʤ��g�Z�C��5�ќ�����.�)�?[꯻���㱮�e�v����W�_�2+�g �t��"��/قN�a����jO���X>X�B#��|��5��PE��5����x��C�؃�x3zc��?�����q�Z��@fg"�4��z}r[��V�X��Í�w�@Z�K�%�$��Zߖ��O�r�����d81~��eC"l9�D�cOA��%��%)"��ըP��)�&���)�ਟ�{e������4֛�$��h��2���[�@X�������a˼e\�������[�Sm��5�I0���NZ��ag��
c�F˶�UK� +"/19�>%�%j��b������]i˄Q�zeᗫ�-��e@f��@n6֮C�f�� X��ĬۿА!i;sz &��B�>k����OS�m�����^@�_��Κ nbܱ�|�*&�L�#�k�W��n��Jfj��"d���f��^m�,T��g�yZs��b��c���%�Ŗ|Q�e�㵳B߷��'J�JS�Ҹ�F��%Y󽰶�`'�_��o���9�{��q֜����Ln҉�����5��]&=�Κ�\y	ғ9DDv)�b$�Ef#nA�[�*8k�����}� *eV"�E=@�}�a���|��o��}��
�K�H>�r]³"���|܎啻�`�o�`:1����M�6T��c�%}	��n99�0� �N�M,|L9uڹ�K�78�'��2iĘ���Ahx8歗d�Us�8�c�.Q��Q��Y�d-:ffF���R��!Ϟ�4F��n\�B�9"dX�,!���f�t<�iE��7m���,����7g2;K��*@+P��o ��Sw��^藖�Yʷ�U�q{�uY�#��uwL� �_�< �U^5�P���(��dz@jmSi<^��>;L�z䛆��hl�i-��f� g�l�[�J��BO'���f �	3���7+��8�.�����$�(��w����J�����cR��]rW��8�kv�pt�@���r$���s���hן��0��/�c�)]dSQ���Z҈y����d��#u��9=�P��4�M�h!Kz��9>�IO�YpC^h^'� �}�Q]�Fvՠ��ɴ�n�z:vk
���@tp%����(%���T���;f������\ R�+�;f�e]nLgXNT�!����e%#˘d�7���U�D��C����^���ϓ]s(\^$��V>�Ohj<�b�\k���G����L��p��ֻ��:�ו"H-�s#eư mћ���da�3���"��gE�ct��m
\\%(*��Ώ��t��p9WA�P�h5\1�򲤙��x���s E����6� qivs��� s����+QW���g����َ���p�Vs*�{7�c�����ڇ�*w~Y�/s0���`_�=�:48P"4j�f�\Z-EE��9����F�y�2����r�^��vI�e�?������ÆB�5`�oG�(��`I�l:G���D�nz
�=l��#G�2 A~ߵή�e�.=��A�#�5` ��m��:��`c�
�Yk�o��	W�ע��׮�8�K%W��Վ��M)ʎ�j5�1��`�~`�3�+Է�_,�>5d>����BH���̮�H��lj�r�5���p���G�U�&2�ÚPy��z�>8.�KG֝��8���76 �Crӟ!�iҴ>�9+�r���#PO�7'
Aoݖ}*�;�0�i�ItE�s)\�Z�������ԓ�1&+.C�C�m�y�>)� ��2�Df��g5o�'K�y��_ ��Q85mi15�0�^/1\I�91v5��j�Ti5�nV�,ff���`N�U�"�Ƣi�_.;���^�\^�1-�-�$d7��W��h��h\)r�$ڛL�d��S����+d�W��u���&<k�<Ct�N'mN�T �ώt�Ǝ=�G����
�&ǼaJDjv(w�<>z<����1m�wG�Xc?soUW�R�__�䳫2M�L����
Iu<� ��������X*��;<~���U�TZL� P-�5�	܃ԣ,im�3kV�`������VPM��������/Q^�S�`�!Mf�L}0�O��������N�?�J4y7���()�LX~5M�O2��"���	�If��&s[�ڬ[�&r�*!������XǕ��D[j4�Z��c^�I5�B�{�D]Ґ����c���������������VR�in=�Aa(2�3�ȫ7�)�QJO�K|�\-���'��z�>
�>�]�)��4��L�jPb��̆ch�un������-�U|̔	N���������2'�/N��!`��7��x�gP������_q3¾ �x�IV�,J�6'�gb�7j� Bs��i �a�������1D�a�HJ��HU)��&!�A�y�-V~����~��k��d�^��/9��U3�]S�=h|>=��5�i�@�b�U�rU4�X�Zٴ(��u�k�	d��砩�-`�1������QD��N�=�IK�+�,�)*=�U��-a_~u }��b�_ͱ�(T�� ��ї)�}[q�`�|ќ���ksظ�_u&{b֭ �jYy�cw]8�B��*�('�`u}�~��k��x���H����a���)�����SRS�P��)�Fo��fG�ٴ��CЩ3<��\����59>v"׀(�o�d7ǉ��K�\!��QH�YK1��~�%��-P���4%����K��/D���wF��s��1��'t])����:(D��є�)��d6VrG(�ts|��D�zu��˻���Q4c���+�Af8|��[z�������?Ż���_�]�Fd��+��f�������a�0 w�����l�t����F���6D�N��d��߮,���~a)ہ��CDr��Lg%���:��C�F�8*�{��<6�2o�d�g��O� ��g�i��)���23�J�e�HJ���v�z7²,�^ܰ��������I*'�3�`DqV���)��Wl(�W,�w �:BO��+<߱�tG�L�wt����kQhC-��9-H�)�������;k��ٚ��|]�e��zT뼕�gWs�(V�w��
�4l�����5gj�5�&q�ϵ�r����l��5��4(F�Y �t���"-�F<y)�u�W��2}����.8�a��aXj�r��F�Eq5T�H/�e�`\B�Q��P�����e̘�8�+GJO�%[)S=�.�7oIw�lt������J�����硸a�T^/�v�nrRl���;ec�;����ғZqb��7j��EPXL�'�p��hN����񖧚U� Q�(�=��Xa��y.77�4k`�_U��]^��K�Ńt�&��sX\�pt���9����v��A�����H�H4��ki4�(����޲0õtW���[�M���w�w��<X�4�� �U��
_�L��o�G>MO'�Ć��2dv@�׾��Y��+pֳԧdaN+O�\��tO	E�� ��X�`VnATI3���x.��5�,o�(�R�4R�C��e��X�_������O<gb	A$)Z?��5���=���â.&��R�C	(��>0�1/+�Z䨮�u$_���2�=scf[�aɝ�[�O�0nI��.�]����۞3���!W}��i&�7�ߙ��.�CnUL�n�1"�X�e4�I���3U�L�{����Us ETc�a��TO3Nc:a{���U�2&��B��22h��LE*���@�1Qp��I�T�9�Ȝ�d־�˲G)�m�{	��K���N�����T\-8�m��si&�a6�ۥφDaYE�<��'�b�n�QC��b�	�d}���{�v-Z���Ǥ6���7��.2?�������p�#��{��X:k	�'�~���v�ٺ����ʆ���Pn�w�;_9|�t7_�q��1�5��DñǬ��^"D��\l׿��E�{ߗIC��Le3��3�)�$��(`�H_W4F��� ��l��Z��#Y���ӎ����Q~��b��z�\4SH�g_��p�Rn����pS.���+t�{�O0�t4Ο?��8�IjDD[�5�ZvY/?1�-���H��<������$[�
@O��]�;��4t,�0�����w!U!+yÔ�;����>�+�Ek��QY��6�qn�S��\⟬y�
f�����x�C>ͅ�Kϱ�X�>��K
|9�&�������w
�(dL���A37��l ���v�0`�9��$�i(�昼n�(U��E��r�\�;P�h�k	x�ٱ�teD���jG�zM�fu��P6�Z�r,�貆��[j���8�Z>�U[��\!Cֱ���N2�V��-�V���wu�5z�pj��s���4'�Pל
Y��z�~v�����S�t��C�ޗ�!�LWX����V[V�]0�g$f�+���t��<]��hut��n�㿫���(3q=�I�"	���:/lg�Ce{� o�{ZwdW��s)�۾�r_�j�c�7�)'jT�߫ �^_?�A��׷���`��QD$3����_yTiޯ�w}���'��sF�h?��An�G#�����������~�ͪ������33'�U��?��^p�BӁ�s����尬R�a�&�;2�21�Y���q�+�Bq���:��c�]��`'��P�Y��p0g������ ����+?uO"�Bj,�Jw��<)I��D㋭Ҫ��b`�P"!ku����
u�"�:뵴bY��&a�|�K�l������:�l�M�V�bt�y4σ�� eM�v%aBt����5�(�!�JeQy	�j���ӯ]3s8(�B�;^>�P8``g�6��O顀�O���WĻW~�t>\�M�N������<R�� ���HV`+/:I�@��w	*��"P�:���I8���$Ǐ��\������>4�W[p;˕�pW��	����*�Wsp�k��x� ���~�]A��x:OR������:��a�&=Ql)"�r9�u"�{�b��1ݾ�O���7h^�5z�^���p/���!�i���p�%��ԙ�{�����O�����^/��6�4;�6�9io��$��Z�N�'�@h��Hx;��^�/�m@-R�21��X����+o=��w�4�E�����4r���)���U�ή�m���	���E�	�F�ډ�x +��ȅ���J�*G�U��l��9����b��l)X����K�����~\�D�Uc��g���P^ 9* �S:�I����m��}��ě34O�pUqΒ��x�*��܄��L�FA�)]�~q��ɢ�^��k-�p��:��(�Pᝀq��M�D���] @�h���(MJ�@|�<�	h!YU��w���� +VPnBn���=��op8��q����_��Ɲ���Zo���l4|Ldt��F�_�s^K�N��.�@'efa��9��-� !)��0��3t`a����:u���L�4f_�~���e��c��z����y%��)BY��nda���V�s0���h]�4�F�ރ_�Ipsqz�ٔ�AE~!�uݣ|ӂ�����������dR� �1L*^-�T�+�B�[\�F�ƑG�����ڛ��X3A�mfar��r;�^ �BMN췱oGe����wc�BbITʇ�k�y6�E�n�Y�ō4�^��� �>?��3���{�]�$)�}��2����ݞ}|�5AX��>@���$��ߒ��_��ﷄ�X���aϽzBA.��_x��fyl�1[��f�@�*�|Y^X>���t� ��!9TfUta9lU_W~���IZ��F�)��߿c�%y㒂�)����3���:�G��I�Y���9�M��Ρ7�ؐ��� �cDTS+�;a��9p�~W��(�]Ef�?=����r<v��v�)Aɩ*�t�!L:Y؊m*C�4_�PҰc�� g���TQM՛��e�ZV�IM$�v�Gt����}��9����m$�!1�wa�=�|�
��9ՙ�'O&1�!B�M��f����-6Y�K����n7�/��"D	��y"���9�������RL������|�m��p���Ĭ�F�J>g&��؀�C�����M)	�m�W���"�Z=\��,��v��"b��V���Þ���C��޷*F+�[���i<|���r�D����\k턓j�)��#�������)[�y��97�j���+��Dz���%M���ﲁ#�ѓߎF͝wy"��v@�8Zd����bS�=y�N����8͇̂<H�b���S&���"�"�C���̿˛@��k�FE>��L�G8_�G#4��J 4S)�YnF�)�<�h\��+��W�:�^9�{4$��_�_�Xټ�nŸ�Y�>�X���س魦i�D��|Z��J�ƅ{�u���+w�2h�����a��� �k#���GCո����]��sly�d1�������ER�X�Cg�#�2ɨ�k���ҷ��(a��9PP��9�FCf�� m^$�ĂrJ���b�)��9�|<&ܣ��o�����e{�;W]J��ع[F6l������l�8
UX�k�_�L�]��M�@	E�q���(<*\�_YB9)|Y`-p?�yJ�ˇ=��_|Ul�yÇ��Y}=z������ @�:���* �k���fQ(���������s�&�r��B��Bt=��0B�8���Me7D��y��VP1�5�K�>ɋ��R��� ��;�$뛘����B(��[��H�Kȝ�-b�8��XX���#q��!����^Q-�vًnH�36$I5U_Kw�J��1�0����_��L;lG��C���|j�?��R�V���勩b�M=����{�<�x,����m��1��~ l-r;�A�^c��|zO�gV`��(.���S���V�����Ύ�/�2b��`��ӓ�V��sy��ҽW:�9n�/�N��e���	�;JU�ܲ��szd���hD� ���s:��(�_����A]՛J@;��m6�Ј�2c%�\��#*6���3��u>xr�7M�УL1�1G���M܄�Q�"�:dA��l�(pF��	�:�B��9Iypc������h	�6�\�)T�So�K6ö�g5�*���L��	 J�JfL&�� YW�#�jg2I��y�o����� ���U8��2N^�u��%���v��X4r:sS/�=@��V��1Y�#�O�YŸ��r�|���h�OհpuB�&`Tk������9N|�t�O�>�A�"�5��j�(C��[;e��o�}�a����o��ۧG�R�94п�0\��C�<*����
���k�S�K?��^iڒ�����F�S��{�퇩��hg6Q([oȗ8Hw���7��;r&�0<����[�g8���9�g���sT�I+sW��#�B
��	�в�+����\��"������Y֙[����hR���;��:�qdf�ٴ����|ۜj��z���"XE��}��9}C�lR�]DR�� �� ��f4d���1�N����I��k�����|#=��$s^C?h�-5�֢�>6Y+@O�\������q������[�s0�	���}�B+��$��	'��gv��#
�"���z���՚�m�H�������𑼋�,�0���QU%v殆1Wܭ{��@M�Zv��� ˝��v��#���̱�+5�1z+��1/l�f�q����,^���+���U��)�lX�M��Fs��g��}���l<"&��8ѫډh�倦��-����L���;��ZO#��v�ѿf���1�P�7юŘk��S�oEڳ�r�-����7��	?�|By�	|���{
m�����.����h	��,u�J(3$�Rn�&f�|��/M]^�KB��
�#t�T���&4"U��ufNr�� ��m�ő�� ����>&y�RM����_�w-��`}��y�)"W�-ض>mx��<��j��HYb�ntO��G]�9�Z�6����x'R����Q9c>�l^�8�SkQ;�X�?��Mu`X?piA)) �D	»"�s�M_dgFr9MraR2J��+�`؄���~	�,��?��.N[��j��r�ƛ^+�Ɖ��ʱ^�en�O�M���da�`��X�4�"f���
4�*��Ir��Y.Ɣ���L��D�i���S��?=�Q�\���Z	`T��c�l�,����6��@
�hu��,��w�t^�g���ߒ}H�f�e<�u�G-��Q6 �u�c�I�~%�T�-W��}�V�b����]�q�}��\�hi��N� 3� @6E�3�o��)�� 8�%��Ů���\^3�n��I��%%T3�>E�>�W���8yha��v���Q�L�F��M+0rEz�giOu��V��W�U�����ʺ���6
�� E
ʂ]��	�Sn��zco5�T����G��U�A`},Q�f��ٖr}�V"S(�o�~�k����ҁR�,���D|����E��2��p�qd ��m�]:�D=���5��Ū+~��y�E���9~��a(�����o%]�U��Y��$�/q�BK~��=>+}�L�Y��/�Y�����~-��r��X���:��i�$Ǌ7T%!�E�s��C�̌�z(��[pL�+/8��>hJN?b�?�A��Y�F���i���? h��"�|#�Uz�� �F����0�7&L��qV��09)���W_����P��[��e�j����Z�)x�nuB*�I�u��T@۲N6�ވn��:>C ��*C�����H?���G2��c4{-&�p��d-�j�8�^�!jN���m��~�K�X�ȕ�à�I4�^.�d�x̄b��6�R;��s�uu��0jۄ_�b����Fu��1�8شQ�={�~�Gm��X�Se�da�g�B�&�}���^�
|������z#�F/tN�x���u8wQ�mTJ�>|N͊%6��è��?j�B	���	�!"�u�~��Ix÷9��|ŅӚq1o:ɼ�?�u�^��YZ�*b' �Ը6��_�NTl�O�"��M���,hW�M�}�@�:��T0�R���w���g%s�9H~��_z�Q3��9�q#���i�����5l�֖�@�nh�K�Hy�f����~�."���wr���\G�w՟_	Ґ�1��xv�j��QK�js��-�?\��̌1��X>�����!��s>��p�%�ђ�1ԃ^拓�j��Uk���۬�=�U�7*���\�K{�;��HזPm���2�mWܟ˾^���5)�MZ���K~��;�a*қ<�٥6^�e�w؞�ϓ~�?�iN���rî�����{Y�O�P�[ă)�A�ZbDW���.KK�:��x!��F��N�a��E�9��i�+�_P���)#�0����b�Ikp���+���zp�=�_a�OR�cpIW�<@/o��4{e���[-�!tK{>�ϐra�:1�&Y�T��u��z�,�z%����N3��7�_�M|;�;<*uԼ��[˘�2�\�%��bp�
��y�]�&��i���٥1�)���.�C���)�FX���|ZWs+�&^��]X�89�}G3O�C�cZ�b����c���]����-<�F�����zU�E�}���ܭ]*�m�ʹ��t
��b�P�H���6��"�J��f`��85�iLf��ψG������@}�?CB�q4ֳk*\"��k��H4���tZ�pU��w��6�O���c��ч$T��KW�9�̸��fdB��������&���z�pͺy�S�O�XZ�Ռ�9��!VP��e���%;tj����2���"G��E��a�}�KsY���)�����.}�~�����騣eͲ���v��e�X�����9/��FY�)1&u�Ϙ盏-r%��,�����N~�Y�5od�&���4Q&/Q�t� ����%)~�CZL�b�k�&��ܩZ&��ysF�̫��/p���#��Ι��Vݸ��B�LU/:l �{�B�,�(˒���� 0]I�đ�4�y 3������9���GW9*uU���l��-�kb����Ť.u�#[_��B��M� ��8���)T��pJ�M._v��jgr\#it�DJ�C;c�ke�G���8΢b�2�	�hLW����FY·��0�
�#��5��]BNmpն��eɜh�,P<��0	���M�Ku[��U�Xe	�.SSS&t�$Ⱥ��&+/������쳗��A�MuupL=����X�Yt�u��A�r�E��>�qmD�&^����]� D�nأF6g�&�緾;gP��=e�A��1B��B�aQ3�kg.���25��W�����z��Ù|\UJ���2W&s=���qD!�3�?���.'���%%���N��]������y�<
��.X����#�0	v
�d����`���W�V���z�W����F��t�~2��q�톅G���eB�ʝf�q��g��ӷBW�,���s��xl��P�Y�>6M�F���~c��4���t�ѥ���՜׽f�M���ի�蠞@��{q"���1<�p�C�eh���7<nD�ȥ�#��"vS ����Y�������O�+7g�6�̦O�¦u�
��o�d���4��3f5��et��3^7E��{������6ǃV��$f>`��|sT~G7�YG�o�T�#)rZ��w|����[;si�h���`��E�L�l��7��5����uRa�n�h�������W�ؿ�a�9�'A�(��G�hb��u�P�D�C�I��ǏL[�J���
o����Avh�TV�|7�����j����Z����T8��<����~���g��_�,�k!���B����2��Y4K0D<P,@eԯr�f��c��a����i��= A�:N��9���yң�j��+�p�/<v1���MT��ӎ��p:em�O^-�����/� ���[ov�S\��f
S� pאk�~-�]�y�3�o�	�a���JS�3�a�Ҽ�B�>���*��5{�J=�	/��-�<�Ni�� �F^�{Nm�� ��?o`-���Z�I[��5Gtg˕��6�u����G���{�����w�"9e�.�$������zԃh�8A.e�^&N����3��'1Ϛ�澎y��w�O�pK%���FbU���c�x*<�Y�UA�b�h�zZH9�݄�@ةy���X����u8q��h'I��sQ�5���p��@�]H!&%�B�P�s���9x?�xe��s�_@�4��6���G����ɠ,��n�),�w�&��E�9�=�s�'�T�[���ǳ����.�.x.)P͓��8�}t�g�̀;��21���8�m�9F�uZܥgc� �'��8�myi:����M���G�������=��j��knĸ?��0MQ,R&=�����Ҝ�̝T��|����:`�S#L��%�S/H����~��W6�r˧�U2��O�N�z�a�p�R�D�U݄p3�J>��sШ���
�w�-��A�XH��G�Ƃ�C�][���f��<���o�|�c�tB��A} )��D�M+c ����Ȏ}���G��}}��&̐
]�����ūn��OGb|X2I��{�.��%a<<���ڪ���%xcz��H�x_����k�O�V �����G��7%\�v.�c�"��tk�C4��<5�`.+���Yl`��0����./�<�!�ݙ)�i�P�I�i;�
�2#Po���Q�P,E2g�ˤ�ܾK���^� 	�2���z��[q�W���ڂ��%lCo*��jv�,i�I�`J��W�4��4��[x⑏�߼���1+�Ks&*�ٖ��ysF�u� D��TVt�Vݳ�<���8�rO��\o�����_��Vs�=ށ��������5�H��YQ�`~�WWv�_�_�q"�ӷ)��sd%g"��"���z�5�p�X:�ZT������؁$�ȕ�W�]�uWT�dIB��n�ƳۊkL
��W�S�8��v������~�E,LG{!��L��4f��ø�{���?����f޼���|�f<M��Ež)4��WO�PX�:]RI���-�v���k���#^�$��ʖ�ST���zF�K�ta��܋-��v)Q^��l�o��o�]��3�Ǜ6���F32s+n~谬�T�NG�C���5V���=nG���d���)��hU	�|؁kr}El����K���IH���E����-zz�
�
���c�ţ8����Cj6Oo�~�2R���
�&* ���hW+��<����u0��2�+��DO�=�/��{pv��p6��Q� ��F0�53�\xm�yZ�f��a�<�ǐsF�5x�N���@p^�J��Jũ�Yf�ɂ�Ҩ� �Ԁ9{��Yy��GX�\����h�#W"�ى���`0d�Z?-�����!L�n{�جTmv�8:��B#���Y���?�ۏ���44i�&�k ��t`��(���| qlm�"�!T����C+���3#j�g)Z*�N�VDI䄾�c4��V�V۹-�07Ho�~Rr���4LZ���P'���{�K�!~�|�d8N4�0U'ꇲ�b�r�79���@B,.�%�]�]A"��<�~�jB�9���?�z�!�,�Mn��}Pb�C�G����|���0�ᇓ	ew+��e�ˍ>HE�Nt[����D�Z�^�ck�<��f/��q�� �j[4�Kӎ={�ɐZk�|v�u�%���zC�Ni:�]�ͭj�,N��"[�G_*+%�=r�E�]��]R �~�Ͷm�ʛ���9G����Yvg֕���a��w��������TB-�̏����Q���!|3Tr�}@
�Ý�]��6rg+�'�V���qo~F�b��#���0���:�~KyQ��wH����������Rv������b���R\�|��E� ����`SYq ��y����a�n�.�=!�o�ຌ�B�s��\=��|��5��������J� �Ӭ��yY�/>,��B@����ĕ��@e{;q-A�mWܩ]�9>���]� ��?�Rc�^�*��)���dw�.3��1�������˹�)��B�N����䗉e��s�|���"���<t�
	}k8$�HZ�A9�H�'_W7�mj���$��]<�T��Y�S���- Q�#
T]K����ɸl��y���H�A�b冿�&���N��S�\��ڙY9i�V�,}�L�4�g<=8�J��X��@��
�����5hJ�U>�Ew�l��D �xR���-�9��ti���ǆ��4��z-ৰcHˣR��)*��#2�|�ܿ�)�_�������܆jڹr4����������PD�z'�p��[�mĤ��.A-��2�)�ef�o��T���TVꈊ|M���'�M�e	_Mz�̶�!�(v�*^�kn�6���o�^'9�~G�x�!L=�����h	�c;�?���`J?}E�+�cH�ڬ��+oV�h�[c���h�	�	�&cU�^k����9�G_.�!�\����Ն	F�Ԩ�������a�DXZ��m�m�e/�O	���E���:��{Q�D0v� ??��j�8��5ͦdr	��Պȧǂ>���ZH=�/
b���ձá�uq��%�w����v��+��3����t��H	�FTA6mƨ�-Q6�4�ۥ��#��4>fp�����r�S�%��2YS7� � �M!���)�������j9%f�}����gy\ >����S�P�'5ԈX�sv�������G��5�S���8~�⑖���E��#��O��雫��
d}�t��5Qm=�`?��~n�F���]�k%�ђ���a�]Tɐ�0��r�N7T{\rl��p��T�������}G���M��T\ˀ�bo�-�Y��hw��ߊ��nǟ�,�z@0�W���Wo�>�	K7{'佁����Rs���3�n�)ārƇ6;�&�1���E��������~W����R�#�������M���>��A�<7�VHV4n���O��k�l�^&�o�|��_,]�� ){\�g��;v�嘶I^mP��񙝔�?c�[�r��m)쯯'�,r�F|P�Κ$���!i`�A4Ih��tF�{�00<q~.��.�#�!��ѵ3ls�%(�iP��j�����	�Gx_�a���7��,��n_���GlRj��Jݎ�.�G1��X<�yB4m$�SƮ�����B@!��������[�&��	k�Po^�89I���4�4��%>���Ǘ������G7Y����~��ZǢ�K�h*��9�d�
���p��&����aձ�`4�&�1��p!ZCÀr>59��ĥ��f���m��r���2�JKp���
��Hs�p�:a�� 2� j[���H�b�Wu�^ظ���d.� U)��2�:�u��vqd6#H=����'L��$��F���І�y�e�����ɔڝ���v���ngU~wn��҈��_V���������,���Ɂ��P:��%<[�|H��ݘ/)Y��Q�r}�����*e���k��`]�8�]0�ȕ�n�N7���5~�k�I6�X��~���FZ��M��d�z�*w���*_(��RBE}�id�5��5�1���xη���U�}�T��φ@c�3<Ss4|�|DRJ��0s]!������������k�QT(��s�`�x�a�U�7v���r�u)Tᑹ����pV0r�^�ep��,c$6��ң��d��|��PrMׇ�{�I[i�ޮ͑��@拉���+�}>��k�	AU�5�r)eT	ޖ�&�QJ��ƖAif����� {C%�T7D�h�qA�Pq�|lޑ�d)��2bc����?y�R'5P�>w�6��o�"ʟ1���^q��<�v}�R����jj*��h���ߒ�I�'�a%nU��'*4��&�*=�������H4j���S��.�\��;�SD�6��t�c*vT�AH��U�z^���Y�W�MH|-�Y(-�	&�x̱�����U �`)?�α��˵������R.Ż�4ѥ�h���<��f���{�@C�?s!���:T@̀��zק,l?�5�a��MУ�B�S��6C��z\Z��w.P<���hu��b-��x�Bb�]��^H�Q19]ɘ4e�c�(]�`(�߅aeߙ?f�q#��uj0�{�����%6 Z%��#��/�/�KP4C�Lo�䗲��Q3�>�K����H�]�iL�C�R�i�og�⛭���5���>5�h1Oۚ��@���*oh�x�Y��d9w���c0�'-��x~?$�}����&C"�#��#��t+A!@Q臡�S�� ���*�[�v��Wt�f3��{䥵? (��JHٔ�K6�b=(ח���՝d���s�e�&8)�rZNK��IW?���Gt�uL�]������+e�`��2msm���$>Is�O��;y�w����Rt��c���x�< �bWGk(\,��:[��K	�+��FP�b.sdm��Y0^�=r ���&�c���ֿ�}�g��]&��pt#F�&�b㈗e���Nn�u`������8�5d�ĒĂb%.חӾ�w�L�n��y��Q,��:/Oz:��;,��8�Υ���jP7U��*��+l�*B���A����X&cS��Oc9��,�}�@�|���~����7��
����I \=�>S{##"�Ѽ�!�#��E�x�����	�ꛮ�u��3f%
"U!���D#��X��I��m�
������{��p�a�[��#���χ�)�+�y�}�'�Z�`{G�kk�v�Nf)Y�ܨyb���n���`������je��\O��l%�6�v=����E�������s>Ǹv�g�E���D�iL��xǜ���LI���0ф����Q>_�>��_�6��b�����\\�<�8������]�6Bbo���4"�ǾN ���w��I6'ws�U������g�:Z#%o�旰o������,�[���?ĉ���l�X��3p�_�ZL�GA���=j��[~RH3�#�9V���_:�Kh�D[��߳�����j&N����/TMIc�ڸ���=#MP�$��-��AOU�S��_�^D�](���Wh(*Iq��I�gYwU����l�^�R��ޢ�D��[����'�ZP�Wf�͔	�Wı�|&;�V}R���^��-N�Zx�y��f��M�xW��2ۙ����e�P��s�����1�Sr��F\^X�S���?+Z\#�ps�R7$Ҏk�(�<����vJN��:RϬ�c/�b��K������ڨ(�*Б|�� ?d�qyv=?�]q�+����rGƢ����*k�����j�+��I��*��и�Ҩ�K���(�KeVa��dv�KD�&#[�aP�[ďZj��'��,b6�j��F�?rQ�!�#�`��.��uziCH�vb���?���u2��	���3Is;�u��-����8�G>�xm�J���&�&Ʈ��dT1���;ܬ(��������<�ԁLD��Wܡ��HPb��E2%
��Gלe7�]���~b���Of@�+ ��άO��<H؟mpܐ��u>��Rxi�g�h��΁�TTb�;h5�����?��>�
2�+H#�J��
�u�+:��U�
�k��aOz�*��S�w�P"���="��kި�ݘ[���H��S!-��ϒ<�\Fҹw�σ�I���.hA�E��s������B�וY/�+�W7m�V������D@Tb.ׇR����!� �z��4���O�4�a�(����6�1�9��-�I{����uA�n΄�r�;�db:=�5Ѩ.I�+a�-��e"fs�F�:U���/��Ue�2�MV�������[�|������lA�2��%w���������*\��%rt��L�h|��g�v�׀�#���-D�����Qg�y-#V�w�>)L��YX�C�Т�.I�&k;���I7�a~��{�=�:g���'�ʔ^��:��	gBz�Ft�{vB2�]�Ur�Bkݴ���)a��F�'��#�|���_�N	v)�yD����Rט��ؿe�S�FFŸ����-�5R����}J�"֢h�NQ��/�l'�׀)� ��d]k����@?K��f�.Ճ�Зn�����r���u�S�W�B�hqe�% �N4�r>�-Y{ϳ&��K��h(�S��{ݷ�a/Gl�L��}��#��$(A��u{f�E� ��[V׋��&��n�.O�X	�:/� ��o���]�U��ϛ�����Q8cz����3�i��ܚ�{T���K�S�:���빗���|\a�b��J�sZ�4��a>:��'0�0�@�%Y��b'�� �Ա�H���/���3"�~�٨н�-a�v���Y?X��H g�]��xk�?���:903:�#�_!�#�fO_A�f. Ȭ�U�;����y�����|���J=;R�������#�|V�PKwKP?ď����ÿn�'9M�Ig��QH�V�W]���a�������'�Z����E5�VN�����?��Y�N-O�>����u�4���:�'j�B��;�O/��t���b�t7 b�ر����M<��dQi��T!���q�������陼{��;rTFR�U	鈅Є.�6$a^OJ�`ߒ�.�lI�ZE�[�y�R���wa'�C�zv��6���B�IHR:n-Т�D�%/i`��6�EG)/c��3ش
tn����^}b% �
���O\Kx�x���r^�zjY	�"8�
��7��)�äއ �A���i���W�w�[͟"hP%�'Qo�u���
�	92����7�f�Q�+g�	�4��:|Q�
I����k\�m���9���Pm�d�FL�М��G�]�h��M��c�4[���<v�p:,v�S��H��+>�4��Ѡ_VEn�#����~�l����=Qe�I�� $��r����&5P�=���^�Q��{l�W��q�zO�ǂe]*(��r a[�-,a&� {��˳�˼�02�@K���3|�U)���A܀Y��Ԍ�'�d�7(��H2�;h���'Ζ�����`��-�݄}����p�RES�KW��vn\<�׬���f�a���;��vf )�1�o�m*Nj�˵C�k��r�wЃy
x�Pj��|I����:�s�V-�~<�V����mQ���h@|��J�ǘ,CU��0��֪�D����j�t�<�]ĺ�T��z��5,=��żo�9L�)�ص��llܣCDP�䟖�=�Nܸ�`ĕuu،� ~��ԭ0�ɪB�3���Jbt�e׽N~�I�*�o
X�#99#���������sH�_�{<��+�v��m=��I��9�}W�'%h�2��Ҷ�;S����
��C�� ;��!�7�B.�ǂ���q5�F���?Dj[b�RREf���d��x���8!�[İְ`R��:?��_23p����w����̊\=@�5E�q37dAH۽��ˣ5*@nup$�����L������Yfūu~<�`����:q��p�v�f�y�͈ȶ��=������K�%(0i͂==��Z��^���Ѥ����-�*�h����*����y�E�vtY`�@�\���NGH�2�y��G�7�Y
&( �V��ҽ%��?A,�����d�p����v��W>��L�Żbr�P!���8�B��kR�>sۡ[U��>�'N#����U@�9c��r�Q��i�;�C���^L�oB ��G��b�y�+�h������e�`��_�WSb�vr}[�T����H~��;�`� Ǟ}��˸�[#՚^�))䢑����1e���GH� "�'������e���v�;7mR3�1e�R�h�͈��ϧ���6*��U/�y뗌�5�0��Z���ٜGjK�Ju���d�1_��WV8&R��Xl��VAT����?ۏ�t�E�h�b�<U��^��k����� �����X\4��5pX@�x�DcW�f�$�Y�Aԥ�7��{R.e���.OaF�Di#�1:������xd�C8B�P�Z�k`��~�]�ɮ�r�jCR���)ص��/�
�<0'c,{U`�X�>�%��I�m���xN��I��<:v6��E��T� �lG�YiE'��������y+��6�Ƹ�_eȾܭ��rx2̨�\̰�n;92�6UB�8�p�F��,\��ؑYcB��U.r�XM���=f6)s�n�׫��������w�~u6#+����(/�Xޔr��x�a|�\�n�BTn��EP1���WR�rje���A	�S�r��\��8������覩���F���N<�c�����^��,�9�۹FV�5�Y+�$���}����9RlsD�|��>��:Q��[ub�@����q��e]N4��w�$j��^'�� n��:@��x���bҒr
BmQ񀚠��윱8BLi������X���e@��|
s�9S�Hwv�'��g��u�*i?*"܄����E���O��c�h�����
+RY�n���V`dR��O����ɵ787W��o�
%F^RN�$�O�3�+G9&�l�XU4,��\Oi��RRU����̓@���A"8�>m��L2'L�9/����u
��V$'�!�Y�߯xk"�C�0,�+ڀ�ɻ���;m�EIE9ɔ�"�Fu���Pw��(��/�ɴ��>p2�A
���P��7�;)�UMB�����$�ˈ����ɒ܉��16��B��	;~���u��R���.ԧa��%��i�0C] �	�+�i�%Q��:� x�'�nD/�m�Ǧ�D/��w1ȗ9���6İZ����OH��T�t�f��u�Qb��`�re*�q����Q����V�pw�E�_�t�.�>�$���������Wjʭ�r�dl	�
��#*k/d&APJIR������?����8�{�3]� �װ�Pe��-Ӑ��ڥ�꒷W�/ �� �'�)������%�C����0l�2�j��t9���4u��F�kBT���D!ﹺaԂj�Em�Š�?%�~��`��@���;������ޙ�L�c"����	E�*mrvۀ�X��(�+s��kt�U�bx�Җ�Ʀ�g����U~SSm�<��;g�B�����e�i�ğ�=|6z����b�(�-����-6$kg� �}�0`�,>�_o�nHyf�M�t�^�����{��X��9ev,�7� ���dK$_�� ���[{��e�����}��c�4L���j�´[�T���8�H�r=$ $���;�	�G�0[�M��cP�n�XClKoϾ���BE� �%vF-u���%�9FX��P9��v��1PO�i[/,����B�(��Q���x�������enV8�}�U�	boڄ�7bv�3�/�|0���A��o��mO�O3HG����˗�E�vD"�UH�u@]w�>=R��!�>�2�a*���MB�VH�R����3nCԙ3��1r��~h�4U��"�[���������4��	\��� w	���,p��`zw�@VdL��T�yI|���X��B�ۡd�z�s�%O��p/^�k����c�	�tKgkt��s@E9�"�7!}�%$$;-=Ks[TW_W8k*�-Ѣ�%���0e�n�C�·��C��^w��Ch��U�v�&&-�ϮRd�U�Q	�hf�rv����+M_��hQF��gib��^M�;Y*d@OZ�� ���Q(���V*�`��o�p����?�n��u����2!M���T�&�n.�;~�7*�wu�/���\�H�r�kDx;��;]�_!J�iD�]�)H�*��R�3�[(������~~��/h����4��8�
���}�3���č(��}-AM���*��e���z���\#�n�C/Ѽ��M&mK~^�6��-�ô��dkeQrԗ:�s�aM���9����$�'&�M)Ie�ʛx9s��(����f���?K����_Fqh��#�Ȣ��Wƀj��^��0>�u���
�:��b&��Zb��s���W�8�Z�����`U|��_P�_��%i�#\�H����dL$v�m�^_�RE_H/�>`&T���Zά��\s�g�Rv0m�ܢ�ҫ�~v��q�� ŗ.d����c��/g�T7��r���z�j�B+��r�5��� :G�2��I�t�q(W\wV>�91���G��n�Y*P)흗\��<+��BXW�+#F	�J�#�����ug¯�S[�/�:�!R�{*��>7f�ɗ�o�R���8�d6�l3��1v�K�E��#w�c�Q�I��~�}�/	N�%�i )�r�;���{�vm
.GF��)ۮҫCz��-whj�EA�;��t��U�ZS����J)��U�@I�D���.�+��y�r����	;V��C���- P� ��?lR9���Wu�tL~xCf;K2D���RXB��w���r��VuKd
�D��0/L���"d�#�a��2PKv
壇��m�Qs�qX$���
u2m��g��
R*::����;뗮����mk����:+lz��;��4W.T�_�w5o��7ï�n�+�|*<IUȗM^��B��-�*9�Z#��^�dEu]_?�v��Ӗ���|����I��Ժ�֧�.=Pn�>�Q �-�m�
�W�#*Jj-}ho6�9e��&���6ꔶE���2*t\��B�Z�M�J�
4��֍Τ���~7�}�c����'"ɕe�#���~&��l���%�_��r��Lqk����G�E��52Mka�/�6�L^3�-f��su��sJ���1���\��N3�������(�z+��g'��_ݹ|�.L����='�`���qx�)�l]o1���ò !��f�JAZ&�'��Z���0Ԇz0���[ �}I/�h��[�癋�?;�%�^����(��i�����^�Nn�[H�"2t������r��1q��w7,��o�h0��m-$U�_��[����� +Z�#u� ��[�q?��8.4�
$��v0����'�Ò�YZ_��x$)@ܧF�'��:9�
�T��uh|T�	��>��@�oEKtM@Dd�Hz�I�|���h0H�3�c�a��<Z���+��1ǽ6�tW���Jv`�)�7��?:K�j�vQJ�dC��w�]x�3�}X+J5�c~U��%���ېG'x�ڱif=}c�J$��?���H��>�\��)��Nhc͛���Ҫ�C�-���H�S���`9���	䳋�:42Ȕ�X�Pxݠ6=K˘oC���`�"����#����r�����@e��.S�w���wn��{e��@�?78���3�[#�9Y5�e���߂;Ň�K�g��)�Q�� aE����AXj��9/��o��r���L��c���$�!���P�H�@4�/WU���A�r�I˰I���Z#b�؄��{X�ÖT�~�J��⢃�O!xr:^���k��Nþ���K��KH�&	dq�b5��t�� �~)3I�t��6�/�w����)�i�<$�1՟Wɏ����4'�]��Vz��5����ă��T �lK>���-�[ 2��������Q�o��`m�w��n��F��1]�,�r�JgatjBOQa��so¨��k�6�-�kT�,�0̬Bb�E��W���M����7WR�U��t�b�*���mݾ���P�y�)�B�P��bl%},S�A�fu�G� 뾮n�����F�\�_�0H�'�q�v�F���%�ơC+�Ά��;�6�g`V�m�����dp�n���������AKV:�d�=C��Ĩ���R���O_ذ�g�}��x[cL���+ҥm<���E:�*QN띵Uu%�w�����s�ۚ�Ah1-��0��Y5u�I�Ё0��OF����PgG�ş 8V��_�t>D��uU4P���@h��B!������m��a������	�s�nO��O����z�Qt��1��x"�����wG�E%[���B?V����{����cAnN���$�FaI=��[y���5�<��t �B�羆c1��:Q��I#�����#��Ҳ��X!;�ϩ����<��/�y��������}9`��z����i�J����4�ѻo��O���=O�:�ӈ��2
�Q;E�U�n\5�K'�e�LN\�a���"�FP�(C��lw�[�[���h�bu�Y�$5C�.¢n�������Q���U�v���ʝp�C6�WH֨������,%42橌i#��q�uso�n�	��	�R��D�vR�	C�h �ݖ}���v/`��կm� �1B���O��~��]����?�OF���e�E�,ҝy�<����t���8�i�Z��	���v�}��e��{��1a��?2��Y���5�rI�Aȼ����rv��@N��l�$�0 �v?2Zv�^��7��U�z��X�
~����>3_�@�gQ��
��i�����L�狳�K	֚�Hm������3k�iR��4�����г��f:8�e�����3����n+�ǖ�֪0��~ 
"bϢ[���<��>�B�q�8��E�z I�b�n0֗�O���ѨӶ� �"��#����w|X%q��%Ss8�(}b.I���.��YOd����8�=#O9�Z�4�d�����ܾ�:Ǻu1]KUaH�-h��,2B�G��%�����f�Iĕ��ur���/��0<��N��֝�E����(�'��P�ּ����zAb�K���T3�7�h3�k7Z�b�@�S2�����P��i�DG���CW�3�&-v�tpCNq�Z�����>��2b�]d�Ӕ��E�(�1	�`�d1Z�T��^�G�
@�f_p�.�!w�6G+�(�T�o��\Y�eM.��Mi�M�[A���������'�c]��3�{��K�'l����)n�����F���yzF1���q(���`b�P�r���b\�����̛(˩����tuc�Z�v�Fat��<I�q���$)��h-��`�V~k������芤� ��!67!Z{�k���Ԅ"�k4�;�L5�ŢD~[�J�f|t��3^��=ҥN<i��v�V�N�ͯP_Xƹ�H�1m�?߯
��-��4���Ru���S�Ɲe������EOQK�=0���z}���M&������T�ö^a�Ck�'��8������Ԍd�X��P]��@3���w���6��mX�EJ�'�8���b?կ�T"W����w�Pp�*����7%~=V�^aF�9Uro������z�f���Q���U-%���i��2]W�h���v�J7����5����<	OU���Jݖ���k�lk^�:��LZ/��j|�E}74N��"�(�'�\$��s�Q��{�@���^��	U�1�jN%��@�&rj�s�?Zr!Ɋ�|+��|Y�A[�N�E9�7\�}����Y�"0�8��<��BS���F^$����w��.IN��F���ki�O-�7Kw�`�E�0����x��z���G���r���c���4D��c�0=��e�2;���f5��?�p���+��ZC]���4��)X�f��leP�A5mE�=��F6�QN��JG�oA���#��NM�p�N�K��j}����W��� �#�+C;/��%#�(Lj8�:'�Ӥ��{ұ�0Sm�]���{Ӊ]6��B~�mVUl��L���k�_�����!'=bf~��b���Ʉ�D���a���`�H\�:�5l1�(`F+a��	�b�[i� i��N�t��1��W�,~K�D�`ty	6���P��8�ۋ���xS(:�����{��4q���j_j��^���jbipAO;���.$��P3�/vUX���ºaE����^���1��O��U���I��/�XN�b��I���-L�W/N�D��q2-�����Xf��n�7=o[К���ʴ�����a�f��䌉9���������-ܯ�.ո�|!�臺�?�L�=�| ����ᅹ�m��SI�2b�?�b�k" �����dY������sƳ�\f��J(�gB�;�d�Ͼ���I�_V0�����-��Y��m��eB��f����Y���[\�aj	۱fHTϼm�r�E�Yc�u3qAg�>�/����k�{�c���#�o����T;a����˕��;Q^��oD�6T}'��fb�79��p�:R���vD��R5���c�d��bGxʗ�*K�]�ٳ�@J9 ��=�u���2W�������BIaX3�M��m�#k��RXG�V����և�����}nv���	oxg�3B��X�.#�B85Ͼd:���]ի�2�@&^�I#.s�րJ�.�eb%�S�����{[���@�o[�wy�x~-A#�{��e`�s?m�I��G��ql�P⒍Guͤ���>�!e�����#��Un��)tw��D�YP��#�p���D�ʅ��gN�� R�D�e��y�F��n�d#�/A�K��EAq�
�� J<�Y���1��LB�=-MG
��A)nw}]+_����2?Q�q�K����}�'�f�T��oH
����}��;��9��3������H%�&�qYE�7�f���/��9��F`?�U����N��_l!�D�.~�Wt��h8�a�:7S�gB�uO�P`�b��~�c�UI'q�z8U�3N��ץ�u�t���m��\�<J��|�)���Il�Ԉ���U�.7����XG4L�r�X��X`9K �*cT+�d������&aav�^�$WfBH~N��}�E���Q�xκ�8�Z��K��U�@lX**�gr�T��"I�ȑd��ث�C:Q����J��fl9:.�'�Ҁ��1��ʚω#<ŭ7��LC���0������\r����:�L�y���R �����w����W}M���p.�r������(ȣ�QV��n���*թ��k�4�ZA�Kh�\�|>p"��bG�) ���gT�*�����2 Z=�?�S��s��Ŀ����
MuՖp���w�?�&a򽀅�7��^[j��,$�{���w��T��C%�u�T����S"��G���,!)H�m�����7W��dWLҢ�5�� \{p 'ՉP��h�țvHI|��|�X���Cu���� 4
����rX�Nq�K�IE	J7i�5�ʫ��"��7�՗���$�
�%���˭D�2�:n|�����o�9P	�{�<q���hSnєg=+J�뒤�n��ɐo]�� ���/bR-����t�
��h�Yݸ1��gV��f� �<!�nfʝ�EFغ#��uFw�o|ۑ(��e2f��N˯�i��XD@��v�.$=�﫳�Ąk��?�1�Ҁ��d0�5�z�G�2*��,��^�2�O9c4���(\7��J|IQ�5��ٍ��C����͊r��ͥg�5����86Q=�r�&BăP��L �d�DQ��j�bHAҢ�7
5?V Eگ�k {��h���$/"�Z��s��%B������T���%N��Ʃ��lI��)��u�1�g ,�˥*l%`
�]�%5Djdw�g�7�ځ��3�/~�b���~i��2�=]zB5vd�����62ǭ��gk���aji�9���a��G��Ώ�C�9�aWkG ��&����4>�K9Z�xH�5\��A�n�R+w���F�P�(j�,�Ant9io��P�t�|�~i�̹�Ф��� �24�G�66�ߴ�/�K����tQ���.� 15ml'6� �_�lj�y)L�
)
;�������T����0��gyk�/�M�w��EZ���@8�X�sG讁T�V�DņP��sg�~!��v��T�(�!jZ�:Lׁc��х��Z�Lg�����1/��>|�����eu{���g�����"��uV��������J:�dв(�@Y��v�Y�R{�U5*�v)�dL'�QJt@ܣCpa�+5�r/˨��X��;�[��>ٱ�}��HJVGXL��G�� X�l��;l���o�el�cd��awK*#��Ɉ7 ��Z�sĸEs������������ Y�D|��yD0�FR��[ISϺj�1v����K�AXBY+�*�S��vzt$���"��U)����!�k�פL'!�t���!�|}��eO��Q��&aju�/���Ә�`�SO��h�I��UU,��rji�Ԝ�k���b����n�Q
̝���I�!͓�8H��� Ƌ�]z���*6; ���M��4��Q<�oS�r�__��l��Y+��nU/�K�o�E�q�� �](�y�8��t)�Lg�q�$Z�#�ޝ�YG��
a?� �\]���C�ݺ:J�d�f�M@AN%�	�o��*����>���h8.s����-���[��r��!�%���n�k�Pp���a� �in�?�S@���+�Ӽ�?����}0 H�����
�[<Is��u���<%��:�d0B(�xq{��>���A �b+�>�C�ȇr����۞����G8�M��	O�kYK�-�z?+�i}F+��T��KWG�?1S�*���YD��=��\��z�Q�ץ��z���r�x�Em+�xT��[/c��n�}πh��Ꞧ���q�Z��8ns��eޣ����gP�1�� �t�L�g��=���_��� à,z&��3;����^�/��}�W�8̪.�(O�~�[�m6/,�Q��r4�ğ�����
qf�w.(M:p��C�0F�LF~"��8��Q?"6Ǟ灴�
H1B��8G(�)M]��N�ݧ��ioi��bCa�����`7�BvB/���ܑ4����9r��wh�f�����&���twf~J�$H��V�v�Lkj�C���<H�F�|��=��1����?�=�4���@���ގ��c�J�җ�����:���10t<�y��Ŵ ]���iL�������p��J���]�?�&1����w�:�*箎��	�k��ՙK��ݎGɵ&�{r��mof�v	?B3RO��+�����4�/�Y�����-