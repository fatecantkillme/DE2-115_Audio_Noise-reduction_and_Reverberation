��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�8k�)9�k���J�f ۘEN�R��>�Ug:�&�1��L�9��b��]D�޻��%9�r��vv��}j�v��dR��ï.�4�ld��6���?�n���r-'��:�Z�a��U;�۟-{D<����F�b�gI\W�]6�R`�q��𙒏�,�<��*��ج0�Y�`�c��#�X��M�� �g�l���(����,���A�,n9�W��q�ҵ����[���47qU��l8.��ZpZ�ا[86t��E���l	��*��*Y�57�:�V*p��1��'�Ha��Z�@��.D�䑦��F�	b�ӧ���_e��r.��z[�������S�du�.Rֱz�OK��~bO�	�[G� ���b�h���L��A6���{y,�N��ׂ�?(3�ݟ��������#�t "&��5)};\a	{9���E��q9�ŵmJЩs-��ڹYHCj�ZK��lP��� � >]�R9��|7�Z���YD������u�x���fl�ȃX1�wW �{��߽��QE��X�Ch2��ӛ?�3ZJ-rс� O�;��kk~<�ku��&��f����~'���MJ,�O���!?�Ɓ/!8��Ӓ�A�4�[�b�?�r1I	��MW���8qCô������[�TL?���Ŗ����Z�#=/��c�X��S��$�c���m���їj �,�Sy���F���]��^�m�޺(B��:i�T��T�@]�v9h����q%��9��y{B]z	��iaMD#jw��Rū<*�k9cNoCr*I���2-aO~�S�t=?� �J��b���Ds�O������X�����َ�ݽ�3��2��QQ����r]<��N:Q��O^��<}d"�I�3��	:��Vp~���KƐ��p��;|o*jxɛ��������)�]赽/�:�;�?�F�o`�#�oɂ|��G�R��U O�R��`��1A!�e!�~��Tۃ�e�7����M��N���i�h�~��0?���3���	s੸}}Tz6���C�)��{k:~X�������=�eji���@�O/�����,,��9�"'ѣ�,R���C�Ӄٷi��VcTY��NP�3����5_�\����]���wFv>B���cPX�uZ3D�3�n;����71�0���5@�w����3b�	e�TR��6TF$a��s��t�o?�XC��q*�\ׅz���n|�Ҽdi�}�?s�X3a��aXp6�.|�^�������5/��{�ܞg�)�z.�<����Q���'�M�-�"��HѬ��>�2ㄶ2���9��o><��l�<cfx{�'5�B����O�BhmaƹȥH���u���<�c\q^��-(bm.�`���e�.��u�C����{Q��|�-/ ��M���D�Mz�|p[5]�+�HU���� gF�~a�2	�$�~rEF�W�`RLoO=ӧ�����S��(�����`+����}���_�������e��xޙm��{q�#�z욣�|�������;?-D�yxZ��:0L&����i_�[%�Ccd�R�������>����	3V+h[�&Z�)AJq"�R���V��`�@�=���ǰ=�����To�����x�淇���.�땚�S�h��b�y��D� �w�������h���b��i�@����b�x�.�V�7��F������a�V��kH>��#ˏ������T���� �CB�䚆�x1��U��0�d�7P]�+K��.*�A�bpG��餳F|��sC�ic��@�[��I���%��~��nk��#���3a�K���$:�{
��lhO��Tበ����ə��tɨ��r<]�9��V��cU ����Ҫ$��<��dx�ix77P8W�;ĥ$�r�@
E#ڞxi5�3���hfj�2[%'GU�ӺvO-T�J%�y���M�|>��6)<�|̪Q﫴F����r��^�	������fP�R��2d���t;��j�L�H��얰Jga)�{����a��5��K}��^�����7�n��s�R������B�mmT�۽՜E5j���v}k��GP�JN�0&LZ�`�3�e���"�ݝ�U�;�8���?}=P\��P
=�ʴL4�}`9~���q:�Ue���m,�b7nLN@T�E����������W�����p�ݟV����sJj�eH�g������]V��nAz���1�K��"�f՝YI'��4��	��엌�`6s��^#�` ��AHչo�j��Õ�Fý�����-��L�G�PM�����мY,��Ȏ�)%��6r�u$�T�؈{?�0l�%��Gk���:�"��Ғ��`�ޟɭ��]r�yҖ��?�ć��$�}���~9�ص��2��CI����>Jp��k�y ��5'?i�N��by��R�y��*�F�٨��h��b���ݧr�p�Ǜe4��'彴c� ���p���{� �)Ĝ�k��no�5��
�(�׈N��⠜��T1�0I�Td�n�TE��F���0At)G\U-yy��K�3�� xo��L�c�;��IT�����f�C��=�د�xNȟ#��Er(_Ы~���	����ʽ۶�Y�ck�k�ׯ.|�H�ͭ�[��BtR=6�G]�CL�n5����������dU[Y� g��Y��gڈ��B��lLÛsu ��֠�����h���J���d�#��$f{2o۱g�HW���Tʏ�'^=�#�-QK����X��$;��DT����SC���-�`��}�ߓJ���<�%��ONF��IL���N[����G��GV�>�eA_��B,�]ф��4~��m�͗��3�����z��n���U8L~�Ug���a`�0�������_��u�S�"�Bh��4��x�E0�S��O�p�oLh�=R2^�9$S���������:=_U��u[}=]$��3�dl�8$?�\���\}5Wd����Z������Ғ:�i��r��{a����<ft5&�ȬI�Dr�`.������_⢁XR��(��G���9䜂Eޥ������n��Qõ�Ҷe�I�I�SA�k,5V��3D_��N�|?R�m��ڵʻ�1�c:�]챹��4����N��9nO�؎��G�^ꏺ��/5V>�t�j.hW>�����33� '/=��2�r�G��փ�E:�j�==���sZ�nj:<��3��_�b��뇴i��J���IJs�w.� �=aum�R�y$Ȥ��Bu�g@pgV�j��kz���_v'܁�(ȤI�h W�����
 Q} p�x�A.9P�=��fû����03%�I����1�{�y04;[����P!���W��ZJ$\I���7tۏLM��,F��X����z�9�|�Z����LU����X�j��dFͭ�C}��N%�q �ͪm�7H���:��av����i��#̓Nzto �V!�{@��	�Gk���e��
���[���@��TjF`��ū]!rn��V�u�qI5U���r�ܥ�7(�+��Qzl�yZ[rm�=�
	�K3^���Zu��C6\ﶥ�9��H$�!.��ɝo~%7'���Y��#?T�j�
Z���4���{��^�����H:�f���#A��a���yQ�����L״��ͯ��p2t���t��4���{�QF�n�<�H�눌�S�T3-p��gmr^�����|0�,�+��TK�t��r7:�:�ﷶ�!���N8���Nk� ��h��N��356�8�Q�6ტ�ɦ"}\*���L�02��7�8X��%O��!Vh"WP/���8b[����c#z1���s��9R����Z��(�*�/�G��$��h�$�Wݜ�\�L��o�sh���&M�>3?�<�4��6;[�����X�D��t�]�����ʵK}����0@%xj���([kSp� �`�(ٱ		��-�م���E^]{L���v�lWn��z �mco&�ק"��S�[8J���Gjs��Jk��Qi�Q��vǢv�J˺v�Wy:��:�Ecq���D������qǲ��
��,���bS�{��u��E~��Ν�U��@ӯ�Y�C:��x]�Eg������� -�.����"_����p��GU��g�el�Z,��������9c����l�bS��=�p�C�cs�R��R���!��e�����_�k�Lg}�2y�X9�>������]��Mロp��(�o�YBt>�$��e��!�ޣ�)���>�`�������Y� ���+l���"�"�\�׭d��ϔz.�]�JSb��~���ħ�Y��G�9�m����	9:�߳�?���l���]ظS!���ӅJ=���8��#���'#_�1�x������0�ȩhrc$�6���ـ�f�N��G�)-��W�2�hx�I\O1?_����� �0�wfϋN	�<�⬑e8Tf�y�"(���&<���Ntge��ɇ_	L��d@v���jqIzNJ*��,~��
�.9t������ea�Y���(PSϕHcVTV(n��w6B�^��4�TNd�>�C_R`�ך�%�ǖS�JC�.�ܘL�O�u�$���0xW�Hs,�d8�+e4�rDX�d�ZU����UP�dA�,A�ո�7��~�����Q�$}=�v�?%��g2ړ�[�<M'c6��5uD�Ae^E���p�7
��F�q�����\	;�c!jf8�փ��%rx�fb�*(� ��@�wr��P��ڼ�,"Iꔡ�d-zB$��xK�
&2e^�����h�`_���6�7������_̥9y�l�~n��!�{9�5��bap��#�W�_�~��{gN�Z�����C�Mv��ZT�����=X\廩2�ҙ���MkB��h����M�@LM����1A����Jn+U(]�X/�5k��I@9D��
=�?� 7
�W
�:�|���:��:���S��k�b*��3�_����±� 7����(,��[�cx�s�J1��W��f���-�f]H4�I���~#+b�ʷ�7����-ۈ�$���@�>i
��5Ĩ�w��0*��n�����U�Ouy8���0�SƁ���	�ץ,ù�8�E��<��'�GD���[WL�+.\���e+�dbؐO+��D�λU��u�7�0}���1�֥A6ުV!�/�����9;� ���Q3Ӟ����<���ஞ�휧J`_�J-`@���ւ�/�䙫���݀	W�]�cŻ���Q�is����0-}�]GRw��$R��Ƹ��)��d��͑�����Z���
�g�<��C6�V��ƙ�j0��j
�*�n =i'oMB;z���h�c�g���6<�@�Qz��K�Wl�;4I�: =���~3>⵽���]"f]͠�1l/��иN+�2|��H�����n�cwsj�ʵ�3��o<`�{ �Bf��L�]��^{n���+�<�Ά"3Z��B-�k����H�a#�?sC�3R��kn�*��W�ޞ��juA �vabbt6ڨS�~�t����:�*���;BHU�A�a��3)˞(��^%k��VFd�u�
!&���v�"���_{2��Y2+�՝�ݟȍ�ɥ�ܽk�H@_��)ln	�d���zev��bzy�)�'/�i�ᷛ��.;��ܰ�6��ţ1>	��l�UW�i��R�}�}cTlf!�Trr����~k2`�&f`��\�spcBܥ}��ۯ;G��%��{���š���X�=�2k2\9͈ƪuц���d�߸�����ͲM���C_�e?<* \@p��5��j�#	�Qyx�z�l:���+8��r���"V�OQ��&�E"���K?�'���:E���A��֩ʧ���࿵�
����Ò|�WA5�*Z �%�W;{�g��k^��-�k{�9?um��2 �<�+��85a�a?�Vv�T��HܾI����I_|V��o/�;��7{���zB�rn����Ε�`����4�x̣Ev@=�;KMw3�; �hh��}0(�?��ь�|33؇�gs����4�cy��Oƕ��|S�p!)YQ�4�l�Ō�j�[�)_���eE�a��RcH�S���ς4\�X�P�+ ��6�ʵ��"��So_��$'B�)Ї^�S	�DɅl���Q��1��ҳ�H����ۙk@b��M�*Yy}�2Y�5�fWӏ������꜆ݢ@�a�Kѡ�՝Ƭi�ܭx�eG,��r�K�)����s���Ⱦ����#o�~����{LD�o��+��\���ĢB���<��C�R��j��)кCׯ&b@n1��֨@ڊF+S)n��ڛj~m7�6KBz_|�`b2�Z�M�y8� Rn�U��
�߆�fH�c��Ҩ��N�����M�p[�啌xa���f��W�y"+5'@�S����̃�����W�[o�D�u)[H���`��j��0T�K1~e��||�y�Y��φjx�zp�B���~F�>o�j���!�r�&����Ms��)ݥ�Ņ��x���-��,�o�8���Zr���g�T��h��}����u?��M�=�X��7�*
���%3/�ܣ}PO��䨫3o{*�]�tqi�D��b������P����p���]4HNq��<��m9j��r[�H�o�R<)5Z�wQj_GC���?~�(t�:f��B��U1�별��o�s^@m��C��Vg������h�� �l�_�*�u����'	6�����9��%��H#��āmɴdW٩�bKI�~Uee;Q����EB	�$�\�z	��g9()��>۰85~�"s7^�y�⯧t�ó�-����-B�}N�!ek��j�񞊦����W+�x ��?',X�Gl��e�c ����l
���6��q���RE:��ʘP� �yٝn|��IUP���c:Wt�o����h��9����A�Q�M�׊ؿ�w�Y;����b����qq5�z���<�i�(7�ח�ң��"w�AU#�K=Pz�?k�N�Q���B�;@��z��p>���P���I5L8�U����2co�`�:+Œ~$��G�e�~bSu���q�0�P�����(db�i0�.\���^Xɔ�KA_�t/[����ꉙLj�����ˤm!K��lEI *�}�x�?A�s#92蠱�� b�@��*�� �ʚ��k>P=��+�W�,�
�5i���� `U��U}n|+ײa�ߪ@���2�h/J��Y^�h�1�pܦ�&հ�ɤ��� �����;���������f���L-i�
(����'��1�t�B���֒�nOa���#6�M��׶��?����K"}f,��ֈL��7�0��&i�|u>�hDYݦ����OnN"�IY�f��c즭ˣ�E��d��V�RVH��*��`΋�oЫ�D9�h��B8D��z֎ LJ�]��
�!�Nٽ�`��F̠\\��o�����6�-C�Ղc���Ahvc�ûC�bNI�d0լL�{u���q-�-^0o��e`�����Rٹ��PL,N���R����_ֳ����3vJ�(aa�F�ܺ�s�Mx�
;����OSv��?U��o� `
j$��Q)��gu(�Z�}Ӥ̻��7�-�/�*�!<�ĩg���'y�3V�ƀy�t�8���m�-�;�]=1������g�h�P�G��@�|�GO�?OG��y�#�=���F>�ߙ�h�ն�g\����"{6�iNd�h֡�{��.�
Y�{�+i�oOG�}Ñ��j�I��˫NT��H96��Y�L�^Y'[a�0@�����%n
�h�i�=��w"����)Z��0�w�ޒ�֒E��W���H�8�\�a텯Oc3���A�B3D��Ԩ{��#Λ�ܣp �����
F3c&�4d�d�zy���F��G��X3`	�]K\�X����g�g���w؊�S��u��f��.?��x�e`�&�-f�~[�(5ۺ�fYR*�㊄]���վt�!r�^�Ga�W=�f��C5��܀�'"�~����]N�45}����y{�V6�;R.bU���7�O�r+�>�ky�����Q#�Y(�*�{Õm0�z7�}����x��1�j-�T�{{4�0=C��͐��x=�5�R����!���h�ؚ���b`���A���<�*I�7�/Z�p.�v�r�R9��KΤO]��ɣpc��*���
*4sj�@{��1T.�Ǆ�Ls���)�WDet��� ��*�G�o3]>�Fr�k��r
��Y���>F	�Q����<�(C��=J��,4�����ǯK	`Ӂm5��Z=�;�E3���E��R�Э�DIQ9����ORB��T�c��ߍ�(�.:�z>�3�Pl�{R���%UG_T��Cg5W�r!5��n����fYOU��T�۰����m 6Ma�Ls�g]�@w�R�BQ��ͩ�w�� �nr���y*�l��7H�i�9�m��X��L��C̕�Z:�W�[�^���P����F54K�U�q�Z5���$뚍��Ɂ�a.�� Q�v�w��v�����L�'��g��x}�/������
�u5V[,�\^�����ª�
����?8���K ��3Y �D©%��I�t� �����	�IR^ ��T����������
���S�s�C尡���n�땚�h|x͍}��k�kF3�h�ܶ�t�}����@�|��]D�k,;��&r�\r�}�0#���z��8�?J�~�٥�#�c��E=������d�#�0���0�E��T%o���a��=�b,��V<T���NdO~Z�	����K��]��X7�ް��6!!�̮�f�ٵ �Z��%n@ll/������<�,��'�y�H��:�������(11��䒈��P�d�Jl�P̧b:���_&��"E(0t�BM�p��J^�I�b�8�j��`Zԝv$�do��x�-��GҼQ�C�5}9Kw�ʌ�����BC�=�����wIg_��q��Pi��2p�#2�lR�z$F� ��59�ĺ����'F���}�o� ��1O�w=���X���r���K���0]��6"���W>P]�{A������qI�p�W�j�ƅ���P
�GJ x�)l���/�?��sT�@g�3���b̸]��K���T=���� ���Zf ;]�,<{ֿ�K�cvP��w���~�t� �Z��g��=慉��9;���8G�yLy)z�2~d���0�D���iɻ�@M��������h۔��[i}aX�l�`��ɋӺ��v?ڈ�ϻrFg:��X/sĆ�#�P�p��Y$@+U�d���ѥ��o�Z����G��X��{��N�=g����+�[�Vx0����- ���}���5�!�Lym��|����Y��%�d����(�.m^������ 	m
�`�r�ľ�{����_�x1�EjF�'����V{�O�"G�A�U@��5�)��l����y��fG�����㳤�~{�)Ry�t&�JWUCe?��ܐ�0�N n���(��mt���V������ŷv�
j���Y4,�4bEN�aޯG���Ba�]l8�O;EZE��9���4q�}޹h��F>��a��x"�H�w���عbP6P��F�}BI$�$��c�o7#K�A�I�̐��/i.t;Ǩ��x���H�+g�8��R��1R�
Ά�u�oh$�1��LW��c	t
�2�h��~���庒\ڝ���-��]L����+s��hU���:]��F,%���:ݎٳ[�mSW^(Tz�e<�Cky*��u�@�nǄ���b�L��.(�w4�r9�6���4�i����!b��$��MG��,1�M���w45��V<�>Fi��(�Uk���J����V�G��B+
Z�9�2R7������t�����F%U�č�2[jC��r�UOK�v�1������r�Zy��B��H�Y#"�#�!�b�\�PTF�A��G/�L��������?-Y�U>3P�[L5�;}�6x8��3���EߌV�����w3��<�z9
���s�"��8�F�4DB�S�e�򍑺t9�H �d���#�,�������5e�O�C>����}C�=�=)g�o��~�II���ގ5%�x����>�7C{��M1>/8�K�0Z]�]����4�t�|Q� ��҆d��>:�Z���H3egl�-d��������Ŏ�d9|Ȑj�C-���=t�婿���zZ?�i��XC5z?gY���c���� ��,m�r'�Z_%��+ WR߹�\b��$�\��#}��dQ�:]Nz�v!�le����,��)3��J��\��+/zY'
��x3ݕu� {��aW����Bs*v��tQG���մ5%���j���� G%a���	��N���O/�|:2��?Q?;��� ��6�$�D�l��\[�	;N�Wb�J\��'�d:X��!vV^�u�c��Txa�ȼ���ݰ7��ٞ��$\���8���'��i�������~x}�_���I���>J7�X����C���U�$��Y���]�N�$�̼ozVo�,|�c�����|Wq�V���ݥ��ṓz���TbA�dT Λ�a|������B�I��}*�-��J��àh��ЋS��V����~7��6~�:)���&>�i����ÉѸSP����C�n�(�qÄ|��D���=`�}K���t��\�z�,����U�D�����B�L�S�y��%�ZMn�}��8-	L�� 
��)��������&_�-B�t<)h6��9|�2�7WY0�خ��O���M��5��	Rڌ4�MU5��y�b�������F*�@�c�n���ι�N�F�j�3�����4�uB�Èf�s38��L�����$i����\A��f>�c!�"4V��EE:O�$��ғ�ׂ���?{��`U���8rw=�.��H:�Ӑ].�"�e}�Z)�!��ʟe�03�糗���IօEX7'9���RU*��7��-��.YZ��ov�m2+��Jd��~�A���l8Ja��{g�qiV��Pt�W������W�^ES��"�rop��&���x��� � ~c���j-@/��ON���rŃr��P1�+׃�U�S4�̓�w��Hxo�1=�]�w,�JɼU��Y��k��aw����yh�D�k{샐↌~����)w����`4�p��Ո�K8�7!��L�Ն<n?Rx�@�Mؼ(�-�$`�9��ZB��8�1B��
��1���K|ɸo�7�0���<�T�����M�v��^1���n;�p	�LN�l@�k�F�+���Z�<����R�6~�m;������L�h�Q�dCYw���v�t��j��\�~2�
���'�����!,���H�C��O����y�\�ȇ���UM����'F���Ja��;ҁ��\f=i�A�L��5�g�����VE���A�;�әj&�T+3�p�:S��+�8�a_��W%�45�?f����u�5�?�R���:C�F.�I��̶�h�:G�y���%�5JE��3t���
p�'���R(�nbrZCj�_�����Sk`_ �_X�hzxE�Pb'� a���͊+���E/8Q63������!=��6�)I��R�����I�ë\�I=��ЖV �����1AJ���?-|d��S�^'x(#)�ċ�Gcc����L,/U�PK�So��*v���d���\��������-|�š�Vp}Zk���w��kIЋk�:��`��D�����P#O*��0��ܔ� }�~�v���p�w�A���<{-ԧ*�"��6�� ^Ʊ�Wk�a\[�u�zOh����pFb5��!�L)���;7+z� �-�ߚ��Y+K�:���<�G�ܮ���ys�p������FW���6�6�0�^� ?>�2�_د��x�/�˝���:�Q{�oR�v�H׾W�i����'�i| �O�d�`���!�"ɱ+�Dw3���t{� �1���0.MH3"�>�
�3s��c{-�"h|^��<|�빎b;⃇h�s9�т,-�;�N4�k0�oS�5�i���'xaU����2v�jW�N��]�d_;"��@�
�>�q��i �oF�*f���+)<r4X}��~��-J����KC��8���0����8*����xÔk��>�7����ā��jxu���çZEN�57v��k���~�-�;����3"RIA���͵r���$>�4/�;	.�g�g�c�N2F�߾zA-�9��\z��RR�!΍~:�f�+�������S���or���y��Zf�m�$ʿ��X�=��b���,�j˲~?�R=/a�h��ae�"�ʏ�#0�a2�0l�2y m`�l�t�07�$c���dMD���d�����i�r�nrw ]�rz V����\��<H���A8��ب�J��~��k�<Bԭ��&����NPYF�ˑ�mݝۇNk�aK�d��+�ԝ����_6�;��ǁ��C���z]�H�U�}�o���?t�����2I7��v�o"��C1xG�d� I��ҧ��e��a���3?~�>R��m�Rd�u�X$#���Ȉ�@��1�n�2�w@.�� 5���a4I�w�;P5m�x�r�ƚ�/pC8�F+}1����15��.��(�j���
*4�\���l
�|�Ԛb;e��I����i(�[>ب�A�Q�F";�`�ـN��ר.��Nם(Ö�ݶU8��"�sm�zu
L�C�%�w�|�߾�:�a%�{-�x��p���~ۼ\��s����P�Y��{���u3}�O���=CVڗzk�w�
�+�� �wG�{�������lwx�����{�z�Uy*���0���S5p?�c�B�}'�XP�U�Wʖ�ey�\�~P#�1[	#^�	�[�ߑ��^K�7�L�^	�p��=�*<1�����Fe��{R�V��K^z�1jW2/s�N,���������5_��\Y��d
��l�R��+�g�aU�WR�0p�ݍ!��l�D�R]E�&5��z��8Ob��40�	�bQi�R�]p��_5�8�k�g�i]��<MA��G�O��G�ǽ�H��I�#��:hs?�Q��vL���'��El2P&�Q�p���)|益BZ\����v$�Hc�p���M�LyL0�m�K?��|tF����H9�m��$k>�±����Ћ����� �a�끔���I�rm
����6�p��Y�|�@��]16�%罂O���;�x��M5ש(��ݑFE�K
[}��^�WjH`׌yg�v�ހGl䧘SKC���Ud��r��.�E%�9Y�M�8���m��Ǫ��u� ���ϩ�#*)�����tD�N��V̞~�k�3�Qr|£�jY�eD&[KXIP�q�$Kd��-��SL�ӫ��<µ��F����JmA��2��o��E-C��~�y H͗;�k��4K?��tw�c��礠�~�1(^G��vn�R?H�Z�!�gI�<��8S+lC��D�uZ����$=�H�����&�}=�ũ,�b��@Xxs�Yhzƀ���v��=,Ã.�*�k[�
#��%�K/,f旔�GK��\�K�y���Ź������N�@�g=]OD���?�I� ��!o(U�9� V�p�-eLϟ�sb�#�m%�k�hT?���gk�j䠳t�`��9x)[�#�k2(����ρpM�6�j��E!��;�T�'[������o���\��.*I��%q��Z��*��M n#`C��Y���!_�"&9�D�	�v/��<�=199��a=Z�	�Z�t4�:�٤7%��6��L���8W0hH$ؼu6�o�O���WϵZ��@�(�����q��V.����k0��v__i��pxQ|w#��Ya�:�L�\�j^���&�C��ƃ�i�[�������>�2ǋ+��d���r-�Q}R�%���Pٙ�L�a�i�ο7Q��ę���֊z���"׶B>ӕ��R�r�tR��ׇsh��׋�ng�9r���h�]`Od�
FE�.@��)�ç&�xe��_Aפ�!"N�..�T(����z�O$���Q&���,&"-����!y=�~��`�nT5�7��3����}R{����q�Γf���"��*��y��_Z�
�Vl�x��j/���7�Q.��L�5�ȇ �ɦf2{.�߇Ax��C��p������\� Q� ���'�f�+WX�j`�£���?b���h�͕����eq�!а~��s�/���sI�Bk���u��w���q7���ɇC�<��\�曕�u���kxts����vl��e�U�T@�7hI�ɴÐ��Ṅ��T��p9M/g��o{����֗�kѫ}�ږ�#�EϨ$�w�Z��V��钪�T���ģ��HW��m�g��\J�4�/���VU��D���ˢ�HSu�n��N+�AjIY؂L;{!5c�T��S��]��i�%���u�;���u9�H$��8ر̋jǞ��P3�O�`�L�����x~X^�Y��X��T[
Sd���0�o�} :�g��({��y�עԙ}EI��"�]�.z2���w}�]1V]�y�oD_�m "�} �]��v'\��|�Y��o�p]��<�G�yfȿ�Hjv��+sk�ގ��I��������\{c�ρ~���2�2�{��u��,Ӕc�U��ј�����z&a},U��]F=~}��S�K4�`�=����tP�x���S�_ν��g>H5��O0��f����I�\�$�rz ������
Ό d��7�:��)ق��OlA��睈 +��|��=Y:� �_dE�j<$��RM�A17^��K�� 
��a���20��`�O��u�lS�1�Rt)�������1��|Y'��И��@��Emp�: ��uJR��Y=.�!�pXZ�ȕ���B\��4ͭ7<���ِ��6�+Ug����PǤ��:n�ϫз��&ĸ�ʭ_ьӺ��R4�i7�?0�����4g�YA�V��RU��?�������B�+@j��8@b��?ٺ�>��W�sr�I��e��|��%�{�����
�65�b�^P©� eV��P�,+b/i����_��h��P�%HjI�n e�/������_:�x>�u�y�VQJom� ��;��
��(�=�mA��"D>��2�>倣�r5�:���e�.��C�N/̓���J��ɇ�7��q1�w��(8 �`_�Q��>��J�R1>�xQ/ҴZ��;�aF�"[�����R %y�T)�#���v��,-�t�Rl�K�]�S#m~��͓JR��G��(p[x�R��+� ��3"(lٿ��hn�t�-·��$!��.Qu����`���ۓ�N~V�DIo��X����yIo���ubݬc���JcPm"�ܥL����TQXs�- ����Qs]um��p&��x�x�I��-jvE�]���(>���� M��2�<�"J*��T���I�����l���z^���z���'z�x�|.�G�:$�u,qz��[�f3�3���-p��0<�A����ʔd3f.�H�S�L.\1��B��Xu��O>��(y7銩���H��ؤ�8���yS�B���s=����^ց�Z�7�
���L��w]}�fT��y�m�)��V�M|��2RmK&-!��^� ��0�j'�Ǳ�;QF�4������6b�L��[�F�"�	c_<W�{2Icx�����P�IWzO��t�)ÿSM���>��t�TE��e~��w'�Z�Z�Y1RB�}e�ֲ�H���0�n�o���J���S�9-}$*�,��s����(T�6B H٫sX�&��Ґ+'"b��}b��K���h����c��ۿ<����"���? K��R�PHJ$��*�g4,�jU;�Y�蟈{'�a��g	m�m����hv�H�����to+3'�Xj͞O�O��gw�O���f&e&����Y@[
 ��K�H��u��p�"jH��i�-�[�SƜ��%&��VX$��{�����\�dR�Ŵ�F��B|�� U{+?�R�m�8Gap���X�]�A����G����}EU96��M�y%fQߙ>�r=��D$�o<k�A`a�ܳ���P��ID�Y���n1��"����ߔI���N�������3kR������H� .�Ea-�ƝF��%�\lg�-�Ȩ���M�ֶ㌬��(��e,��Ha�\�(�iCM�g��'�J��ܜ����//��]x�Fk���Ύ)VY͍�w�*bK�k�y��e��u@M�;��!��D�}Q�����#��D��a�jL9�����{ҏ���m�
���r�ͽ�,4�T	�DEX���g�x� ��!a�.˓=s�&�}�0�3���
��'�[�����.�d�u�c
-�ѹ���� �g'M\)Z�/��v�������Z� ��y+�����Q�����F�n$~� G�lЌ��G��[W;N�-BN�?��כ���Dt(��F8L�W�n�j��-�S����pf�� ��2�bu[�ˎ�t9i{T��CN�� ���hlr|�t�z}C�!�io6`�����$�T��!*c�	�)�y͊�i�;��1E��dM�}�ʀ���fC`�Q�p7k��$�Տگ�mH�x���ٴ�h^c V��5o�r-�"���+���C�����v��*�c�g�447r�O$@^>>ϱ�§�&tc�[ȹ�p��^�?���R���6ν�~>~C6�
�S����N��42n����7ԪZ[��z��ø��?/*c�{��|(�����r
o��+�v����?Ꚑxr|�u>$H���ĺRE���HG�^%e}�j���� Gl��y4<�{ �TYr\\A�A\_s{W�6�iH�����Դ��4#R�E����[>�%�"_�LT�A��{R�F�,�t\���0yS6�3����:q2����ȲC��%t_L�wA�AP��B:��;G����x����Ug���S$)���M��Y �ۙ�6V�QH�����)���˛��1./іZ���]l�ɻ�fE��7[�$,�=���^���ѿ_~S{"}b���^�86`]8;��*�����ߦ��G�����߇UΕz�s�x�H�`٫dx^�I��?}�:�����5��V��{�T���=��ϫ���l*�!z���|Ql�S��}��(����iW�g�����J%.Wq?2�,K�Fϱ�Mߨ�`��o)sK�8�h����'�YV<��M�J��?�?����]�������Y��&�����%�!���f/{���#�3kyp�9T�}d0�;��Z�I*�D�=��}��#q�{X�Ğdfk�\���Qrñ��)���֢�0!� �i�� �a��/ITl$P�oW��{�� �P������3��-�9|���M�H���o�L*^/J辵W���J��	
�vz����i���n,dp��A��%H��E��SqƂZ�ܽdm�pxb%z5dz�^�o��h7qy%�g��P���#m$Aa�Њ旔d
o������}+����/9��@�H�*|����g��	�t��?�!������nY��2j�b����8����_��B �5��F�h�M�`���EeF�d��<7��U����������%A�v���5%s�(�vbE̤��De���.-��Iw�C�v���ж5`�d�<�����-��e(M�5��Q+����(�",�k�"e�%�<$�fD���<�	%�s��
f�@�9��g�
NI.��` �Cāi��^v���㎌�@���M��?�9V�2�N=�A�j%���8��K����{�L���2���@,��hK7�a�������������u�/]�}���+��:�>ON  Ǧ_�'�q���T�(J��f[�"<6���{���y+3_^�j<�I���o?X+��؅�����	�t,2^/�?�̚�8��g����n�"����1��\&��zީ���\sb��%�n�!�y|XKF�r�7�����h,�����'�O`}�D"t�����b�|��ن<���W����R�J�Y�zU��x�?�1 Ό�/H�L�h�òS$,���\���=7�{1	��]�I�!���f�'��)��:�M�����A!�a�G� ^���<��-Ь�c�{�Y��G���R7�G�k��B�"��"U���T�9�?�z��>i1z�@Z�3ٚ�<�pqu@O��Z���iz�s�K���&�b�:ޠ�I|1�ș�t�l��8Hͱ�X��$yZ��p�(�T��z�|�H��6���D�*V��ᐠ_�X�h����ו&l� �����g^}l)0�R�Č�<#��q��,����z�]�%&IN�u�ս�㩂%MBE�:�۸Ŵ���l7p;��Fb�բ^&�*LL�{��=��)[�������2:��(�(&;��
�|��x .K����6Jjs�O���Eeĭ��:�p�4#~��"�������u�4u�p,��x0�a�	U69Z��vb�r�\橩�2��p�L�a�0�ed-�_y�p�rP7���*Z�p�B&���بkT�S.yų(Fo¢pֶi�ú�MG�:8�	�*E��ɝ�Y�ݮ�����ai���p׿��ri+EK�HO�Ǝ~y�	cɉ�+7Ðy6�؅ds��� ?���+NӖ8�V*`*Mtf�8��9Ml�� �X�am�Q�1ׯ�j<Ʊ��@ulQ�h��ڎ��~���=Oc�gS�0q�H�|���ߑ1?�@�䐻��0`B�-K��nc��o-xص�d0�X>��⽂��mPwW0R`�:(��,���$��3XzI�8�D�:Ϭ��W�Ǫ�3i�c����:�;�{卤����iF���7�Mt�lՙ�*�)m�3���D%[�kjvܾ�ëN�`2��Q����u��CQ
U�؉X�ߩȓFr%C���bi���`{ɖ�a������!V5u���9�"�milB�"7�{����6�r<���NܖT�
���D(qp�g~�����muZ}~�����X�JgD>��a������Y?��λ^���E|t�q�pv�O�ѱZO��$�?Y �8�na�ne,���x��J��>KΦt���M���uK'y�TA��+@B�����������+����J_��h�Ɛ/d�Xu��v��;!�1g�%�3��C����7��޸���{i�If���qS:�2��Lb�o"R�o�]�Q�}����K>,�f�SŦh��p���J��������_ބ�MH���=���n=���Z���z�]����B*�7\XYF���w���u\�:��][~sW�Q:A_SZ�B?��~�:>�x�J;�x���hcoШ�r&e@����p��L��L�`�zܲ䁋 ��Q{�B���]��e�2 ��΢�qzޗ�5OT0���w )�-�0�Y;ب�'g��6�`5�S��]��;N��a��
	v>Z#E/OmW�"��# wS�"�M7��m!HA>)m �*�M��M��6c9�bD��97����u�mz��%������vs.ճ�o�H�S<�)�=YK�"yx|��#i=�8�o�=�4���K�%etF��+*�y+Kx�*�`$�ҵ	��)
)�K%�?�m��@���0���]�"&�Mq8=��~�AD>���1�\6�3y��Ŀ�d�^�c��:����$�k�<�,��j�>���bS_uu��I��F�
�ϸ��5��q��6��gg �k��V?��!MG��`�<����>gx��2%��7�WU�&�[u��%GM��'>�DS�иe�ϼ\S�Y�����G���>� ��W�V��Uyy���O����`m�e����(Q�M��v�+=P���Tø���aG�^</͖_�CF��O�cT��X�6���ǔ#��2|�F��h��b��!��a���M��S�]X�B#���O�
@?:6y��q
�˖ce�I�?���w�Y2���EU��hs�um6Ku��.~�?���b�w}	rE��VP:���fjWәq����P�z�aw��$�l{M��q�������-�:ο`L);9�eد�7�2Q�0��cS��tk��g#��������12!Z�_'Aϱjk4�ƥ���7�Տe���5��9[��*ؑ��������~Đb��� ]�בf����*�F=��0�}o�izJ*a�#�
�G:Ʉ�y�2ِ7���:z��n�b��u�ej�45ZV�L�_٩�^=�aZ�^�kr�2�3�N�r�V�zs�����$I�����*��U�ɏ�hs��d����b\r㈈�b�V
���)�ua 8Q �Б!?�J5I,�B�	O:5�Qq���wh��>t�8j^ʞu	��aA�������(q˙�j�n���QR� �ٔx��UwT�fS��W���h=����[���s-+i�"MT&\�^.��mA������ϑ"F��o��ۥ%�r�v�x�j�-�"7c"��P�^/�no$=��Ą=�T��p���6��HFpߔ~\����;�����]	HY�T �\=���o:���j^�~���{о�Ͽ��
TF4�����U���h"> �0r�y��to��&J�� `� #Z$c�i���0�n��0���{ypl���'��Do�����6�VE�S҉��O ��9����o���P�`s���
aR�DO��q��%������&�Q�١QK���K�)7� �۷��j~�!lo���!y�2^/��Na�}:P3`F�l��s�v�dk�5C��6��]��e����6���"Ӱ�M�+��B����;4`�[�5��������}�~r�i�$҄d{@�[7Y�"AÝ,�R���n"&�7
(t�GJ�_�٫��]<� ���&r�;������g�P���h�G,j��E�%Y��X,X6N;�C`{��>��2� ��Ţו藆k��X3���?9Ӻ�ɛ��B��Y���m;��"!�jSq,6��i;ƠCb�oo��~��(�V�o)����*�Cܧ�����E��>1�iE�?M)B	w-��%�)��r���~ 15��P����7�H�4ϱ���eƪ�+���Z`\�v���t}��-�F�dE� �Ιю�<���9�����[�t6D� �V6Ζ������H��S?�n�G�)d���F嬛��?ƾ�̽�#X-m�E���i?*�����7�f�l��!���u�g{�J�aZj���/zZ�2Ĵ
fO/�G���ߴ e6��8Pq���D?	�$Fk��IA��_0���-���
g�6j[G�+B7w)��I{. }�~ݑ�	�8SXt��_Q%X@�;�P����f�>��3��U4~T8�k� ׎~�1r��Ǝ��W�Z�5q���N�h���鬭��'��E���&�N		�},��,%�R�4����8�X�K��C�i2]�5!��Q\�4=��&'���֊�;ke�٧n��ּQ:�fMc�{v�mL��F�\O�&���y��v�#1H��������+���a�?zH�H)��D�Ú; E�nIHY���y����Ր�s��G�!��הY׼���c[f�y)uw�j#�:��O����3�G�1�D�j\�	���|�k!�n�Z��`��s��s�t� �� }�&�Pbu�D�-�[���ȩ���,�a���5z:�{��R������tWn�d*���b�!���1cz3��ڜ5�uƃ�����Nl��.	� d_������v3�V�i��`7���:u�\ �f�]�>:V�?��<Ѷ{4�&|EN�;���ߒ�>*�L�ڽ2L��Ԓ�Z�7#[�%c|Zq��8�`�i2?�PkE�^XT	�|��{1&�j��;R�k6�^V�����1��BP��D{ɞ����3�@�o��T9p\f���eh�l��מ�&d��u��|�~%l½oA�+t�>�4���,ޱ_�������RB����M2�d*Kb���6,و
�Ac��n��|���a�&��F-��`���83�%o*����f	#�I�`���<�2����rż0��`����~�1�1Q�s;�p��Lk�P������:}���N�UB�N�4�+��Ep���^IB��L{NS��*4%��"t��K�G��4��zo��rZ9E�:�6�ch@?� �m�E�o�L>���2H�+R����A�^U��´�MO�?/��`����Ŵ!��j1�~u�0�^.�A_�1��N���aϴ��$���k�7�(S��K�cӻݽuO%F�B6��F��#ݺ��ʇZ؄1G�ylL�C�\�Bڥ<�X�%�u��z�؆��|�U=+�cV�|��|���U�`4���҃:�8}�Dz�u��1A�[��v��GC�8nI`5^24�Ҵ;g!�7B<�&�e���&����[܍�u��_R?S��-�-�)�$3�g�A:���	����䠘t���=��E�:@�i�`x�WK�׳�w�t�d�M��w���"U�[J9�Q�q��,��B�Y����)zZ�6W~�TI�"hkg�P�$i`�x�\��?mܧN�w��D�o�;9����`d���ʹ̭�%L���Ou:���c%);z����m����]����˫�8��8�v�'�X�>�I���������.~2�t�"���Y9��O�7�����J�s�N�ÚUK�$m\�H׎��'o���W���֑d4�F�Pc{����N(�5�J�̥�3c�H�/7�Rsyi�e,T���jy��֢��0X-��$��J�8�O�ﱙ(������B��p�C�U&�j{;u�WY�8�olO��$�o1O]b�5�{����'����G�2<��9��*Zo�b.�p�ƈ4��TQ2�̎���� kM�"㜏�N��C��Ң����Mh�T����nJ��5�۾4�Q�;��M>ÍP���iƶK�v�3su�kSOR7���a�b����e�]�冤]�_W��� �;�!	�������E�kdzнd�#��ŻY��n6��������e[�T����9y5P���e��ӁR	OQ��`Q,L����_�eEȕx�6N�k%{4��*�t�~[=�r�l;��E:������{�/���ӱQ��0�5�=�\�;������*;O��e�ꆆ�ީ���*ql��Q�<���ʁ���@O�At��l�����~�[�?c X],�ؑށ��C?l,s��'��[RrW�>nD#-go_��Tu��}6Сu_�G�Qk}��i'1�%��b]z�2 �3:8�DDP�]���`%c� ��9nq�JU�_���z-4L�0�2]�&D b�4_��%�\�?�r�j��F��	�nYp���k�����H�h;��		 ��/�����*?�v�V:{M���|�9*d�>|Pm�@۾C�&��{{w��Md`��pEQ)�Ƣ��O�)`������`ӽ��t���/X{�^��|�63�Δw��c����Iqx��B#c)uh��'m�l�lK=ı���"�Or��C._.f����ԏ��{d��]E־����a����1u.�M�A�������n��DX���阮��x���y����r��C��uT
ߖ��3�w�n����f�QH����x0+�x���R,HpT �W#D��KI�ޔu3�+AT?#����Z�G]'n| ѷ�\w�-��h��<�U�wm'�m+���ju�v�Id��1g_ˁ��z��u�}���j�i�@���ך*�����$^�^��x��.m|/$�!xp�rٝL?� �dʆ�Q��D�טcEih�R�F����� c��#�/O�����[mN76����֓M�������y�Tm^����~d�u<���
a5�U���:)�6rE��(��ݩ��D_특6���4�|�g����9�;�B3�~�ʸJM�Uk���Ź�KLtX�U"�����m��
��K^<��.�����������y2�VoE%{̛�|��\��	��* �J<�jS�2f�V����z7��D��0�+	б�\�$��ۑ��&&�lO��&<�CVգD�Z��y�)�1`�LK��y���W}�a[Bf?S�n��0���w�*B4}���.�~���u)�g�X*	������=�Xs%���+�������-�a�:B
����If�`]�tJ>� A�C�Q�*����PA�0�w;��V�k�N*�@֐L����u�t�>��M�'�K��)��P8�t�
ۭ�NMm<q��"e�ފv��O8����n��!qp��p5��M�J�nȣƀ�d*�T�Q}*A~`V����3�=Iwh�X4�#�/�ѯM�ȇ9���
P�zْ'�`�� z�QY���&��] {V��Oh7��i��;���b��r(��R(+Ϣ��Ϡ����Z}��%~�}�,�#�+�u�M�Z!�Rzx��B`�=IP�v��}j���7��h��f78��I�`��ƀF��a��H�1ԗ|/���qz�w�E~�+�b(I�/S�(�I��6j���-�h�'b°/��4��M�2�ka�ŉP�Я�)��˦�uP�.\A*b�81����HrTFȦ�2:�
��D�� OF�k{��F��4�`hJ3���2����Ψ�nPL�}��]oȶ����@UJe��eG�l�g^����)}��x����\菉���-h�d�WP�85��
�l6�Vd�^���Q�9�>�W������,���,�h�z׺e�o�2��jq���z�4كhD��A6�N�ӌ�4.^�pJ�� �_{��T�P��g��A1��b�����i�����_yq�uG���E;]*��XUQ֑rұP>��O<S|���7֨�rnG���T�S���/ûg�=���j�b������9"�%�ir��0t.ox�9G�!�?���Jq���m�7@�O�3ݱLc^����.F�f����L�q#PK/����V�p,>`�sUVm�����2'2w{[/��B�% =���qP����X��΁#O��?K���(����VI8|�'��@!&FU[/�f�v�γA��LT�j�Gm.^���Đ�-��Bq�I��}Jr|���������������>p���n��*<����������<��_��	��էa�5��BEg�E*��7��(�E�i̧.�RȲx�҇�!� @�����~c��=���]�еK��'GQo�@�D�?�	˺>���[�wg�Z��&�#)�p����İL�{����/'��x㪊�F�q�8RD&��㩖D��\N��n����2\��A�}n�3P����6�����*v���ˠ�Zß��X�LF����i��9J�M��%,�B*+xN#.������Y�j�Z2��f-L}��;�]�N� �},BW�lr-�)"3er^���ȃs{X�=؍bB����':�����
wG�c�2��
v����9�ˣ�5��O�|01�k�@m�p���,�oƗ�)yrH��y�͑��v2C7�3L7��&�����,j5mg1��{R�\�����8;[��׹�:�`:L�-�?��[���ݤ^:{a�K��r&s<�o���59?`�F �U0tخ�	gyw
O��Q_O���gн�{��O&�e�+��3z���@fN�e��e�ֲ�c��8x�KϜ+]�x	����cj�j����K}o
.���Pb���Z�k��*�{�Ŏ`:�fҺl��Ȟ�ì�LTX���O������M!e��
ߡ��2�����h(%̳)�ڰ���L��7Ɵ8��Km"�C�w���}�'��B���.��٢}�"��\�5Yl�L�t���nA�_����H���;1�UGsg�嗭����n'��fL��
��̂����$Q^-+ɰ��?h��ĸ��T����i������tUr�Q���T�Ľ��DL��b#����@$����6��Lc��g �؇fFU�_����B�tĒ���̕��ׄDĲ�T����<)XXT�&�{�	j�ŏeA`�|����I+K�9�ܨ�g{�E!�9���,�b��MFJ"> ��)�����R�R^2�mR�Ѭ��$p�%�{5��3����RMp�������Pa���N[�&m?܊�Y+�6@!���ǡ�ų-k��]���[gn�~��Iӹ1���VbJ=u�d�U(��r��$��)L�%�#$?y�eEZ�փ�\����':� <<�f� կ�2>@d���I�$�{�����X�A�U�L�.�E��S�߶�h��]ar�T:�A�]�k_2�A���8\��ׯ����A_J;HB���h����F9���(2�͓��o�ѷ���Ru1�Ͳ�-���c;A�M:.����������ϩ6H1E���I
wbLxZ!xI ���b�U�Vn�{FЩ��AR^�{�u�y|��rQ�wr_���a�!�6��|��שv���
�+���S���+�Kv����g��F�0��9B��sV�	ҩ��8�F�c�w^�A������҄�޿-�d��x�\)8��5������a�.�����:�99�͔+�FT�>�BѬ5@zuf�k��Yn����~Ua�і�dv�P�?��"��(�Y�*�������[>v�HN�>Fƭ>W�S�6���oK�͘��_�8[N"��U�~�͡�v���9>a�QJ��(��r��,���*fD7�]��fL�S6�ݝq�T�{����ӭ�kܷw(t���[v&%�]�� 8��/q�7k@�{wJ�������IX�{n\����"��F��R�~��Y ��eXH�lC��;��}��մ��.G�b���_g���(vst�t8]
�3��<�&(n/�
sy�%��T����g-_ی��\���J��}rڡ�����u>�#��՘x��v�K�R��0�Z��rd!����W,�/*�/�qb3�T�WC���쌅T�8�D��Æ
�6�**.uЊ=�#��L�����Z!2J
[^&Ѿ�[{������U��p�WHF����K(����۪�u��G�>u��k�蛵�ե�s���vI@"��r��m�7��̢U�|�Ur,�vǓ�T��zpg(���4;(J�����*�������'�&�}�)�;xP��k���"�R�s��'{$WO+4�|���k���]��s��lWb�5���h�[E�V"�!ȑ�HLF��Q"�����v�"�& Y*�W�y��V��N���7��aF��f�%�<C�S�SC��\��u�
��4��V$�;a�cGՌ\
+Q��`�-��f�&lr1f���/3��?�>̟(�<�)����utL���$��1*g��S~�R#
���8��a(���yR���v��	���v�N&��n��4�3���R`�����]�¥QX�W��4N�0� U�J�q	N� �N��Gy ����I6r��?��X�+P�Q�B�=�pQՓn[W��"�o����i��(jB����Ĝ*{��B]�s��p�\��Q;��s�V`��1�ECbf%+3�����a�����F�p(��o��Z���w��󪆠�j�s��J��U���>.�8��hPt��kZ��(g:=�>��"�A��z3�ݗI8��M���6�T1�<��Ѳ��3l��
~F4"a�r
f+��{,�_�aB�t
l�1W�F��6$��_,�D9D��3_˴��[��o�:�
~- ���W!���������^x����E�o��K��cG���}�=
=�Sot���;������ױ��Lm�(�S�����ip�P[�U7���q����N+�Gc�D
�[�$c<LD���P�<^h	�L��L�<����C�+�Q���cd��U���&I��7�J��#H���?���]Ɇ�g�m	��ٯV��a��=�����k"�R�����NA$���M@��о�|��� 5�É�Ac(�
~oR �;ArR�2Q��-�u%�(��������E{s����E��m��-�.� 	f<]Q��b�gAd�Z?�&B��;���cF��~��T �{)O�eJu�8��W#q�t���;��}n*��,4ѵ�%����X�y�R��q!]�=6�cԨ/���@)�_��<Mh-�L���6��U�n�c���mIRS@�m�P5����?����ޑv%�3;K��.��"$�4[��ǳ�/Pn����fxCl�Y:^�%�C��h���UBf�B�A��0�hj�ɗ�·���zB��gz���ٙ��8[b��.�A��d�Y�g|���U��7<��{�
���1��X�.����qf�z~���{�o�\8�l�/�f�._�e���P��z�E��U�����pŕNn�'��o��N⿟����
�u�B�.���>΂%�7j}@=�;!7~���ܲ�
R��&k
�Q����0o<��Q>��^��jҌh����~M;C�jx�N�̆�PX.B�g�00;u��)̔&�a	�؃��J)'��
�D(��^P���f�ˀ���7F��@�%c��J.�6�VW~i��\��L�R��)���X)��5���� ��*Z�k�#�˧�(�!�Ӳ��»�v�m�a˩R��s�Q���u9���~V�h�D�(�$�~�{S �*掻������<dg��i\Ywp��f ?���0�w�G�����O�طM�W�d��պ�~OF::�>� �tY�!�G�1�`G��J�]ogv*�x��Θ|q]J��-Bt�z=6	�x�E����(�*
��(1��K�ܱM�a
�9N�l#����}@��t,1�G{qtK�J	�y�-7��Ta�7r
8�o�n�qJ�g��,!"�����r/sk^z(�j)��S0V�G���_Q�	a�Â]�
u����2�<F�w��'ᦔ���(�,x�	o��0����qm�Ox+)��J�o�{\,�},��r�7!E��OS+�0|J�M�D'^`s[����>}{̙ۤDF��G�Ѝ'R��!�����p�ЪP6-jVr��z���=����	�W='񰄋�)�"���=��l��@fz1(y�5���%�w!�}�W�<T�{s�Vy=EM��5!l��9C��tS�^������U�\JC,�T`AB��ڂ%zEӲ���'u��h��������* xsw�c��=@	�<lQ��a�M	Wk��"x D��
�7xR�h�F8��*��FRGË<��fK�w?�����#>B�R:ޫߍ�}�������ڍ$j�Hd\֩�ī���!����ؐ�}���{<�Q�9���R����O����j!�F�Z�V���l�����Zl��n�r�^�x�u���u8e�i�0~��@>u�Un�/5Ũe��ች�d�Ӿ�8�;��U��G���\Vm��Hj����������m<
��ϖ����� �E��<H*��A�� �G 2���pO��Q�p�����*����2�d>�b�E��&�Łt_"Ժ�M4�J��L���E+f�����h_����-}N2WG_��f���ē�z"����!�Ĺd��|�aC/��,P{�}����l�&.6Ӊ���I�'[�H�|���*�%b�c�!U2�5)��(1_`�C{��LD�+6�@��@����.�;r���Κ~>��*,����Ը�l~���*�����-�L�Ջ�_���M��Q�ÔԲ���5�*�7!b�`���h_<igV���#"@^�����������~�ְY�P����	b����µ/p]�z�W���
��t�R�d�ӿ�`T��#��ib�l	�{1�[��A�s��*�)��F˛8�@AǎC�l���������O��y�um����#�l�.4�?���`r����s���e����!$�uz*��n7��E2��1c�D�G����U���t/���2%�p��+��A�XU �NA���W)0x;��S
�<��tڜ����^$c?���
�`�<���H-e�M����j\�w.��s�u=B�>��K���,�v ���x�Q�3��i��R���VCZ��M�+}cu���[V�ԋp�D�W&�i�o�n����AO�K�l ����0��ۙ��+�ֆl��N��g73�`av ��2����%R�9yG�Ǥ0�>4L�Vن6�"���b���^�&6��q���q��bw���1ݍ<�F�T�x>��{�Wҫ�@yXbb��tU��3��Uw!.�����P���LX�?�����͠�F��Z
6P�!�,d���+Ȏj�nc��+���3t��a����.���Q��:�C��E>۱���D���k=�G�����6s	P&|Q�ϝ��C�(�I�#���O���g<y�����<K^ �r�9U�#v'�8�&M�#�0l��+��!����(��ذkh��OI������UF;�S���b�kM�{{�3���a7-��:5�y���V=�e�᪬�>��=~C[��s��yKAx(��Bf�9�5�=�����U���]���K�L^�F�j��Q{ ��_��#���B�pB%h�m:iMJ9+���P&jN%u�
�q}�C3�ek���5.ϯ�<�#���h��c'!R�}��Je'�K��}Xa)0��z���ڞ#Q�̠1t_h�J�o7�g6z�0��B�Z��h�D}��Yv�=qY18�Ih�d�����v�i����؂Iz1r$Z�v� ���k�y��WC��Ct��ޣ�(�Or������ՠ���ێ��p:	���Fe	��G�V���2Þ���Z�JGP�Gț�Q�!P쾦M�v��4tVWS5jQW�3��L�ߐ�p�AX�e�YIM��&/l(	�+Z׹8:I�N�lo|�\�Ŝ9�A�[_ԩ�`����˕".���ӟ"�3{r�aT�����38LT����5�劮��b�.�&�i;|��Sl��	�p�i�������G���j��t��������t�  �Ȍ�_�g��"��P��~q_r�7��i7��M:;��=m��n����le���s�$��I�����fH�Py�8�X���2Y��%�؍��	��6
�R��_zZ�Śh-�̵�A��d3��q���UVLYL!U.4�	�Ͳ�3���̊��$���v!��?��Js��B�"��E\G�c��L�τW��[����ۏW�p���H�G�3@|F�|jXܧq�2v��z������#~�P>;�v�H}�����i��O�;^n���՗?�a�e�E*�ۈz�q;	<T K�[��mB���p�lA *Xn���U9Y��¡�7F��Tyj�+2�l��Eְ�U�r�[Y���{A6jO�V���,l� �^�fE�,8�������^	�PO[�}�d:u���io�%��J��c�z��)�����W���yp�S
��O,Ŋlk/Ι�W!o��Q���/�o��=���]h�������P��f��"0CfF�9��-�W�a%��_��pJV��z�|����ü����g�Hq�|!o˺پ<�vo�_���t[,T�]P��1ʶSsb�%z�h��'zc��8����L��4b�	Ph)r��"����!�_oU�;��X
��hx��:�w��WֲH�R�C����6�3�nd�&ڇ���q8C�,�95�n�4z��^#�/��E%hjt��0����̲}��E����V���J<�?�*�ar\���7�/���/
e*��`����e�����"�+bBH7��0"�c�^Q_��ď¢Q���* �YQ�.�J���?�8},�`�DE�%����J�`+pz��\x-1�Ss�k�t��������]���)XQ����-ː��Fu���'���� <+��������#? Jw��	')��m�,4�CIqv�O9B�u!���-2����ǯ��T�\��%��,;� 紻c0y?���U����o���#_�l,+�ިz1�ꪟ�Pb�X������`��a�2����/JҶz5Y�ЋO�
����ޟ���S�/48���3�R��*�b���H����M!8�����1�"���o Ѻ?�<��/����ɸ�v��¶{����SI�a�ƙ�9��RV�x[�`%�n�x@?�z�(��U���ٞ�j�ȸ±3��t��F�f�#�� ���sY1{�g�~�	-0Χu��3�jV�~����F'��&,���m����9o��%��������E���9�~ �<ٌ��y�ؗ�kBY�v�����KDVy�Y�z)���4["�2ΪK�Pz�
J�tQBs��+K����'�]b"�rD^��n�96�!�H���7V(�*3���������;��N#qݠ_��&�ń���#�i����nN�S�����B���?�D�]�;m��@~L��:�0dS��� �~VH�)����m���8�(m2�^I����v��A�xc�َ�؊�!���(9�iR\�&~,�k/����F�I����P#@�L�(?g�?�I��-1<7��Zm���6�v$���s���ux�ra/��1�9�'�u��0��}��!�
�u�5��=�������S�!q�m8� ��W������!�i�..��pA8�2����،������I>��u��h��wL������Bu�!��c�n�ӧՅ� M��}3u�I�C)�����6��j�K�}׿#��k���7����?b�ڝ/,�<���N)�Z����֏�N����������`9oi+X�v�o?x�G�U3d/$��ܭ��yKe�|#w���@��H~k]�CySS|�Y��،*�	K;���7�Y7E�a|���-��P��1I��'�~�V����0|w�9��K4����6��,����#�
�Z+�˾rX��|#�����u��~������䵬ע�6�,��
V�*jd%�f�2Ѷ�Έ�k������
nܽL�;�@W:���D�s��h��K�>���O���� ���^�����V��,mp$-<�K�4��G^1��NeǇ7iM댕�m�|���kL�t],��zp��[S�����ݜ��������֘�P}��K��.�2d�"j��+�!�n���)s��%���:��	��<�l'��S͵�)���E�����-�.[~� �ԅl7N�������M
����<)F��Gf�#5��I��c�o��q%C�O޾T�AS"G-v�˖}��5�VO��ky�D&���>���Z(��-�L�mx�}�7�[�o��u�_�1/�w��-�i?���2�4b4���-�o�=��f�/ώ��G[���j�J�c�
����cw�8w�5���g�<��[�vn�:���0|� dh�$c� �/4�
�U�鑠VI�a�
y��	�K�\�w'k�q�
���K?�3�<�1��%�J�g�s�e�i��� s$[<䄆�E�������	��;B��֑A��I,���hؒ���̾��Q�+��[�{��f¡�1��dXg���
L�u���˅<���8�՗N}���U#��إR�C�w�TS�5�9�6Q�����ر���u"�5`�y
;��ǜw�Nɛ���g7����_j��96�w��aZRbY��ik�B1(�dl��tE6�1݆ĳ���b��f��cQ�xp�V��k�� W�y�>e���`z�ftb�{��z����\H�ߢ�d�-�0���F�Phо�;7Jz��E_�0=�t��,��\�E�U��ч��l�'��b��a�*&g�2�&T�o9���Q�N�EwO��~9AF�]�(=��6?7�JK�
<��0k�jh=N�G�^g��:`�e�t��܍��N��l����:�#��,�h�
��n�vk������YH���*��a�F���z��[c��$0C7��	i��`�kγ�F�b������:.���!��F�Fѝ�l�X|vhw��d�v���p�~ 0��Ӎ���y�������%� ����>j��3��Y���C5t�"�ډ�n��WD*1|=��"�1��8c�Q�R,�v�	:A-��oP�$�I�W�����lQ�����m<-��% -R��'XJ��>q�~F���uS�5:<���JFĊgD��w��g�ڏ�V�������#��?��Y�?j�F�P��a�8���8g<Ν�@����Q��y0�\����2/Z�щ�V6�hE�?X�Ǻ��;�%�t}�+գ���w=X	�D��&PE7U�)u��xw͇��-hfa�걒��:N�V<�)y27�Ke�qy0� σ��9՜G�)=�Z4ӗ��!�L�aq8�=�R�e�n"w��3�r��Xn�O��!�rF�!�3�T�8���c���Y����9��Ȼ �s�썖9��{GNb:��P�������j�����]s�b��lD�@F�q�]N�p �\.�N��z��V��x)�F�|��ţ?�w��%D�B~�6�^=�xjG�*�_��թ�yf��#��e��~�*@�˵c���{�FN?����;<�A'w�ĕ��2�o�\������+8�A��V�kt�������	�$�Q���5��vAL�^o�>�_7�r+�-�
	�1��� ���C�\Z��� 	�|?\ٝ�R���7��u���]h��3Y���qla��/^��\,���rX���n=�p9Yt�y܉�ޒ�b�j�B�MB
��_ޏ�E#�n)���5��:�#�d	��M��\��X�<�2gJe��'K��맘PL v��H�J<Ѯ���|��7cɦ�8���9�]"4��;��d���KwFό��kJ%�Q�y���+���b6�V.������O�=9��M��2���757[�1��I�#���~�u�����z����`�`|p�)�3�$�w
:��y��r��u|�'-�H�H��+�@�T���K�߬x�:��ZR�!�s�E�cܼ�Z�$����怐���PR����EE�^��17���1��w5<�-I>��uj�~��{g3�;�Ǆ,n�*����y��G��ۇW%�)��D����P�ٯ�[������㡬|"sKA�d�>lbw�� /�)\�ys��x�$u�L�?���'l��GH�L���}��� ��솺���v�K�+żu�z��)�F��3�����]��0ql�g��_+�[���Y��h�Nnԉ�$ʏ]�j��� �B\�}ɡ�.�Κ*S"�5�ЮNaq��{�+QC�Q}�C�yRN]c_ɚyu�?tt����.xF<	�>�2כ+�!P`���/����Nym�=����-�N��b���~�}�����o$A/́�ǃ}����C{�h�]�?�=.�G���L�2RgԚ�$
�΁Pֱ�X��L� }�I}�9d0!%"jv�.�R����T�!*�d/k���O� �������Kz5�D2��Ӣ&4Q����,$�)bc&o��U^����۴��x�eᩤe_���]���4�|A�K,p�� �J&�n����C�P�w���Je@�(_nE���G�!��/�Ai� �'���;6k�QDq�q����w.
F��1�_����E���KӋ�!*�;�-NEQȷVG��"-����S�~iE-
���þy�Z���xUͳc��pRs��]�YA�O������ju�֭���<� �hH�v��x,f�u��y�^9�<�-�n��!� ����p�)��.�x���ꌝkm6ﴌ���S7C)��Hq:��)�u��0!ݍ���jɋJ~g�Z�⟩���~B���7x^C�$7�� uv/���vG����Ն�sƔF�lC�ͷ�S���mMm�� ��daʹa�	L������w���b��
f�Nn��n�מ<[?k��O������_t-	LHs�JW�a��p;�1}��l��̙C�|�\�Ǹo�Jg��⃶⾛/����$�v��r�I;l`jML-�G �IKWv�jA[-���tIRY���'ӹ,�a޹�;7A/e��<�����{lGP.����%lUM9@�� a��G��m����i�V�wJ�����\({2��,�{.������hwN�+b;��KB������7�P�}���rR��di�ɧ/9~>�4�449NJ
JEG��� �q��j����l��=_���d�p��~��'���-�������	�N�j��3�,���g(a�^غ�'����HV�I���zW��d-��Î���p���8��W 7i�����n+��b��C�NH��"U��J遮	�@oS�����H�齆Ɵ��O=�(�ur'�(�ՠ�fE��-���z\��DA�����15��s%��M7Ħ��R�%������*�W�p	W�6a�lL�*�>��]d�Y)cn���L�"W/�܂8j���%���}�1���SHX39���֍���Q�X?w퇸 ����鏱�� �˥��_��[���r���r�7
���*���T��X�`���v��i��I��$�<��T�fg,�I��Y�q`�)��$K�yo<dt�Z�E���� 1�
��.���a�B��\!?�"�^���b)�=P �"����N.�g��(L��5M\�M�B0������_�OR_%�B2.W^c���0H��J�p�zaД��)y�#n('���C����XT�lF������]��8��݃DeH�ҥ�,cr��fv�qJ�]�D��N���{����q!�~}*�ba�.�O�f�e�1�1�ñRD�cn��}U�y�٨6�5����.�X���=�K5��M�ESt)��?�~��Ǝ���D��;Ku�sO��i��=5��֚hX��}�E�*;�ȠT��iy�*BTs,I��|�4'����g�k������'�^����]���[.�N���閠R�la��&�s�\����$��V�R�������e9������E(�H@���"-�
>�G"K�����I=�Q"�;bشH���ض���s������/���a�^%�Ժ�&	E��W�Ӎ�'�fr���b(ⰵ0��J�i	�Vݮ5>��p;xs�"n/h����\�fg
G��{��A���(��؛H>N�+�X�:�b�`T�ە��6���p�bT�ȉk���X��Q{=Z��s��V�!�pYEm����-)جd�����b��BI�(_Kg��$<��A�,!���PR���\5�|Y��̺�}�|R���x։F6>"��%	�߱��NeT��k� �Y�DG�~�����e0�'r���*�E&C�������1*����) ��x����x��je(�Is'!��d�c���ܶ�w=U�l'S�HH�$w�S�	�1�b���K��>���J�k�F-R�'��Z��m��-���o`�����5�Y5y�4�u�s�0���?G+?�
�j|�m@�OO)��[ɸ��stxX�k�Lx��b<� �yݏ�m��@��|����(�%  p����lc����K��Z����I�Ģ��U>�)Q��7���c�ͫ�tv�{:���N���-ӱ�'��.���fƇ�����l��
�<�\K�j��C8D��"!�9���dq����W�c�i��|��q~$��<+{r�V�6�|"ڌ�ܘ�7���Gx��o!�g�vA�^ �[IY1:�X�og��N���0���#~6�X~�q��"e��7�q���X&I�]� ����@X�ߋַrN:=ߴ����ޢ9��M6<I;1���#a��d�N����[�}$�Ï�(�I}����@?T���\�4,�fi��Zk�%�L���[��il
2��dָٍC�Z*�9���#+�u�?ؖz�����`�2�Wڃ�*2�B;,Q;L��$��������rh��k( �6����S�U���kȫ0��Fx�^tTQ>�
=�{�F�ߞ.I$�x��m"�^�9�'1JPk��s'P� ��Qr��p�̳l�ɴ:Q����/^>�S"Y��b*x���S��툔z�h�g��'��k��n���u�y��ۦ��\"<=(��4a&q�J��a8O�s4'�A��^f�*�����G��
�	�Hס�T)�z�f��I�e����(�^��4`Y�`�&jK���{����w�����U	5p��.�!�Y��%���	{�]	#%��]k���u���<)ڸ��Kҡ�h�e���J/%�3�*^Kv��+��un O�8Q�hL����:��a1���F�Y6㫐��Bƒ���-+ĔB�01���%ߟn���3�la���G�ljB=��ίќN旻�( �İ5[�W{j�y\�3�Ӊ̼x,�1����A4�V��]�Zó��?���ݻ�~�����i��Kj�cT`͌��\Ѭ肧��Gz�.��C נ��-A�D"�.ԕ3���-��dx�r���?�U����� D�J=0��[�'�O�O��䕊�!L�E�v���qP(yPKt��
i��!�k�g�B �#��_��ї����FHL��������U�a�Z��۶����ً��)�`����ޤ�4��I7|���Q3� �2�	 �Jӽ��ۖ0#Ӭ��cQ����N����5лq��%?E�!{
���K��
������US�7� �	��E����iq4��A�d=2\��H��`m)�r�2������|��uE.�OԘ���xgǝGu@�an,;�/���A2⤢�z��bO�gݤ"��T;���9��֭��*�,�S}�g�j2�֨�#��	�N��{����"��T�I�a����]Ǯ���W�	�)�R�'a3�q����=Ίs<�o��I��m�1U�9��Y�r�O�7�=��")���.�Nm�uO�����]�cȘ�&t� e��|>�q�����Q�ME��s��/i�K��Ȇ �d��������Wӂ�R�z4;n���"(o 2y��t���WN$�߫%�j��lM�إ�<Eŷ�k"�����d�3�e��l5)���.��E�LE���aH�(AYw�[3d�E^��CI'+Au�]���ٳ%��l�ȗ��zʋ-�������ӿ�6K�>#:a�<�K#��G�zIb����,�::/`X�LŠt
"zQ��7X�� �i���a�6Pݍ�52т��ʹ9�!���X���/���7�uB%w�ۃ���v��6ȗ?Bv��Fb�X,���Î���G�E�yhQъC^@�-E
�qzD��Ija�Ye/�!�r�hB�(2��͈�i	������J!Lk�d�%���]�{=爥��A ���/� ��3I	)���Ṫ�gsvŽ��LNZ�(HF>|��/:zpEhU����P����4��x��V^\&W�U�|���	%;� ^�u���X�B����<$^�dF���()Z�[�
��8}3���M%�IV�d ?��&iD��v-�ԩ��Z��7_����橈5y���H��ʩG:w�\Q�ϭeǱ��,� %��ㄢ8��ϳR�����<։�Yd����$��Y��ظn\m�5�-�r�wHGʯ��  d��Nbdv����2g�<�=f��-v�K�6W#:�� �]���hHcJ�J/�����	��1��TL���4���v����9����[�ZE8���3�%�%��4/Vb�Y6k�T�e9�8P��]�>���E�~7�]b��K�2��c\K�C8is�`���i/(�f�pot%�����߄��)l��K��,O
霊ٛ;.4Q�^:h�P6�nHuU�v�@�kS�4��ܬwα���RK�5F�
%�̅��uf`����E����y�(�aK�+�UJf#ر���Ѥ�#w��1�l���W�
ګ�x���W�S��MLU���	�X'l�CA�#�TL�\�Ax�k��Ժ�#��	_�!
�qUv����T��Ө|�˩�H5���#h�Ê�O��/n����5r�wX�p����ygb�������_�aF�w�N*�W��7/�Ԕ�L�N�M.�0r�"��-��܊��[_���������(q��¼h���y�UP���k:.���$��H�Y��̥JIG�Z�ɻ�6ԺL.;q7�
g�e�"��MCL�oSt���^�|-�氫�aO迟x ��0LAɻ<h
8m�W��.�8�r�Ir���]�50-v�ڣ.2e��Ͷ
E��|�ֵ���������g?�b'&,�7u�^1[��Ͻ?7Q�*~��Z����=V\�I{��R��\	%̙=�iQg�e8l���'�v��ɣ2Lύw�-r^�C���
���X��\�A��0ͻk<JY�1$��}� A�-bڙ�2���k6���� G9�����Q�		�]���ug��>��{ۢ��Z���Ӈd{�=M�au6��%Od��$!���y�H>��8�+��z!�<ǰ�������ڠM�pK��_<	��8zJvI-�۱&�R"߭~r������M2���|\̎�K�(_v$panDx7Z���M����Rȶ�e�@l8k������3ˋ��q0 v�d ����t�&�m��}#H����	�{)+uLy]�5���co��Kih`z�����q�T�ȁ®N��[)�EgU9�����7��[L���� ��#5I��b����@���l�)%��q�=��倹
�
�T;���#2'(�R���"*��=y��ܚ�QUP�� &��+�/��U[B�`��*��UE������Ae��E�ܼ��J��@�>z����=l٨����L� �<S<���vR0$��aƫ�Pg��Γ['��.���p_=���i�6�E��d��H;����6�e�
pkzNQ7U���5.>�iٿ;9��?ɏ'=.����ݦ0�we�r��i�J�&�����ro1uT�!�T"�6�~��?)ɪ g}�&���%Ռ���j��K����3�w�E�8l/�����?J� �hH
��탎Z��1�
D0�� �5Cb��Z����������>���c�8l|��+ݖ�l����G�<�fT��Ơ��6�hOBʼ��� T�+F�*�A�����H����a�S����K推G6ge�1xu��^�[�Ҳr��"�+��F�5E�Z5�6Ms4�� z}�~��ʟ���ka�⁍����tp!��b4v�I&��VO�ty��	�2���S����[��7��j�/>���<�H#���3��ge����Lkt����ၭ`��ԋ:�{l)�nv�-�@��8��A��O�%C�/�:���6����!T{}P��f�:�K����#`iRW��~��<�ܒ}�W�M��{��;��U؉:ܔL>7���k��`�9ZC��/M���؄��s���8�f�N�]�dZ�G����%�f�%ȃ�Q˶�+��DaP�qU ��k�!��=d+G�x���Uf��W��Fɸ���=�Zw��,��N�t�=���A��ywRㄖ�a?����5�D�ښ[��e"z�r���f�P"p�%�����5WcE�9E`()�9B{E,Zj�s�~n>��q[ $/��x�@=��2���8��c�u"!.J�(����T��r%�2hTc|a6�i�"��^�Wh�^l[�
2�^X>k��%��ӾOEO���Y�;���� ����k?����i�� �F[�$+q���ц�.^\�y�MS�qY
��%Ki��_�Tu���8��=˃5ߺ4���r��В7C�����`Z 
����ˬ8�G���%���<�K�G�Ix5�Ǘ�1bD�Lo*�)��� f$9dk۱�矹u��Ҫ�����K���p~�Z�փ"�K��x�;oD��MroZ�����6��U��ū���<~^��\;�?�G��;'ү̹��j�O������+!���˭��G���m{W��U�CyO��)Y�ad�<��`�p!���}:H3uaV �Q�dHj�Զ��jg�cj�>?t���P����(_yb��K��|
�=�#��P��v���h�,�q|@c��Zɔmfv���r|?~��q�g�͠�S5����l�ђ�����ƕ�w0?���R�f�"��8�O^�v;9��0���&�=H�l��#Nf��9�;s��Y���g�cKXR��aAk2���Ea�듕D���F��P|
�fΝ.<�L�u�]�3$�U����vij�^�� �հ�M���M��Ǟ*9�i@�C��������,b"&WJÞ���ݜ���Q.t	�\��3q�X��B�c>��XQ�8�gp�b�#|12��I�P$E����hw�n��ű��d~��]���jZֱ���1"�AJ":d��[�/R#�\G@�o3�K �~L���
����!�\�L��͗K��ϊ��Wo�m�-k�іfH���}P��"�4/B%Pc�F.$|���X(qQY*.�@�p�H��V"(�%y�vs`B����LVE3��u�
�f�"�}/�'���W�B@�����U����8�[�����d���1��# 6��SR\c��үQ�.��k-��_�QI4�fY�9��J�b)��#ʍ���o��.�{�bn+}�y6qB�V��k/���|�\��b�� �0��~�S�/wC j�o�έ`�)�E
�p�O ������������77�v�b��i���<^Z�MT� ����dq���}~����#K�js5cN�"�<�">������D�C��=��ft��wϤ�\�h �t���Ǆ�p�ñ~�}������%'����܈PΓd��g3@�6�,��v�^��r<��W�9�����<�����wm���;��o� �"�и�Մ����+��� ?>�/7����&��!�fI��ك{O� #n�%��-Oխ�T�`CF9x�QFe�D�r�^�-^-�����Cz�@��+~nB(�� �A�Ar􆇚+L,)w�UZ�:�L:�
��Zs8�a�5h0"���lG����1�.�hM����'y]��(�!\�;2�$i��E�)��vK��՝.��C�>^�w���\'��
���c%)��D�#b�xp�g'R�7$z+.ʻSE�<�f�K-<y	�#>S�s�/�f�<+î�b���_}�{�4i[��Ϟ$x������p��S����hiQO��g�.��g1�����r�s�7�U"��r�i9V,F����6�}v�SG-��!&����6%�7��8�{{��jT�B�:��Xэ�-��A�v�2�e��.�4�����[�Â�*b�[�1v�����e,�c��K2�m������83J���g��M�#<��a��f.��i3�J�쏦d��v5�S�p�8,�X/i��.C��y61��#D�`n�n�CA����ܼ��䥎����͹�$
�"8k<��2s ߴAWqJNYW�O���ۥ�{9�v ��ǽL�}?�	.v����s��ڼ 0��[����Yf)��`fO|'A{(g!AΆ�s��Y"�=���]�a�&��:i�yh�,:Jꢒ�J�� ��|p��Ё&lw���s�ٔ�5VY(
i&FV6���s�0�^�d�D���MY^8��r:e�>��?�(=[{���MU�NvL�M�N���)>�FHm��Z�h�&�;�J7���*P��<2reߤ�p(�D��6�I�����D���9��g��4\b��=�
�̓��N�,~�P
E*_e�pU�����>n���2LT���u�r�ٕ�4�~��g3R+�it�݇��,�(�AEj�ݭ.��s��i��Wn�~L�؛6�O9���M�o݄�<�*��q2V�F���^&�+"�z0�Z�x�JY��d���i҆�05�|`T���4�Pg�jRM����4�ה�/1iЉ�k	G�32&
N/N��a@��/����V1��M���й(���"��c�ۑ�q}0�奬1�3'���	b�j� ����(o�$��?G1L��T�Eb���tE��_oRs\P2ĩ�N_�z����H������k�S'�A�J��=$P�8�H_��V.&3����#뿖7�E�,����A�A B�2N-��7��F�)��Y{6NtS�@���b��K�Ĉ�����љ���F�o�}�� ��['CF�������Y�����:
�ض5���{l���L�Z�G������<�O��0�Ҏ�Է����AY[V����  �pi����p{'ų�W֏ �� ��;k�s; M�K���#Ĉ�O��K`�E@n���^��r��_i1Xi��Ջ�����R��}�?,A��z�L��q�(*c�F"��	>D���u|�	2���`���Ҷ���Rٚ�tC(*gdPH�"��Mع#n�R`1�o�����T�_�񤗫�3�t
>��S֘ˊ�!�d{��O�BۛE�Y9j9p#8�O����?c���r.�)H��_�_� �'�ᕓ"�G�Q�%�l���3c�p��!H(boܝ�&8]<��)bi=0�z�o������O��M�G�4��u?��1�Y����n��p�H)���ko�ʹ�պլM��wVk<U�WfV�w���,����"zu���f�!�r���H���߁-��u#l��nۘ^�т����u��ZA$�E�orIB(�L�%<�B��黒a��&y��L������o`�Jp����Hz���:�Y�iF!Y�����:�Gf\��G�竵`���s��g�P��j�+�o��=��'(80�H��/kkw/�$5�CAm��n��eS�`��t��ϭ�ZU�{3�t�o�d!>u._���e�%`���5�gi�T+��)!��G�F��� F3��kRĦ�[1�oe�R������H/Q�~�gyD�=w� (�~x�������&�ۄ��)�V˩��>�W;!#{]�R�d>�m|�n0*�����,�r;C��$R�����l��!�l���c+$/��+su:���������v��k~� 	��&��E��,h�=a&��mX�/ë:���2�Ƅ*@� p����kEw��䍪|���r�"��s�4D��~
�+4_���m��f�P�;���`���J>@�l��ZW���p�{�����j�&�E�c��~n��D[�NB鞷�\���G �T3��Q�����'���f�	�wq�DG�n���e[,(Q�Z	Y%V�)�4�|k��^���j8%ø�m�$$�����41�c+K�.��Ջ�0�����y��_* 1f����lYa$C߀�0��q6���d��iJF
���:p��=y�_�By"��_�a�8͎9������2蔻��F�B�����^�<�mW���6�C%�2?�'�*��S��~U�$Nr�Vm\�B�!�i��u���|����o�j����»T��k{�.�N"���wݯ�{���b�xI���¨�T�N���*./��݋��@\֦?���q�W�4����FR�Mk!�mL��=�D��J�4#���z�!����2�:A ��o%]�Cx��]��1v{X�!ȇ��6�3N��"Er%0����7j�I7֣�����U�Pb��/gY��݉�|F��y�eI&N��{b/m!yH l��ϞX}x_)w�����6������WM��׊r�5�,�C�o��,�S]���(�J�_ш9��#ZF��u���0�$3g:�i��O@��iЎC���h�5�Ӗ�\c!�%�N��e:Õ6��i�5We_���h��F$5Z����B#�;���K�1�-�Z7���/�/X~�4�7<�2��N�N����:5a�P�Kw��p�;�RN��	蒇o����8��=��R[I�4]y$rs�6�CN�V��è� H�:hg�������a�>;�b��H���
�3���5s8��6��FVld�tCZFn�'$e�)����\s�yz�n��0�	��y��y�o�N*�WkM�z�u�I��4��K��I�Щ���ڸ�"��Hf��҈,sM&��7�Eʅb�hG\Չ��.?˲W�Ӣ���gg�ʴ/l�`�|�C���օ�V<ڿ$3��ec�W}T:�{h(����	ҁ����ςT� �:�)j�pBe;;īU���n&1�l�n+<�O�m�{�pE�$��^��O����,��,���D�T1tQ�͎�9Ɵ@I��̉
^��$�83��`
c�G�B�J:��m<;��^sr�K'�'�U+�v-�:��\2[`D��\�R��<���n���(�uDlP����q��S�<Kա�E��IQr�x�3��D�n�9/��V��b�KO�I]��7��[��k��� cK(�f�w%l�R�fl��v�����"�ڻ���<���8�OD���-���x�"�\n��J������`��'�����O0i,�U1%���;�Y&e���F����ظT�&��q�"�R���l��~���P�<�Ĺߧ\�谊��m��<B�cV���㧢���F
�zTW�ZGz�s��9�}M��x����C��(��K������CF�jcHy���BI�ڽ�49OB�]�A��/'��T.?�ͤQ��:��� z�a��F�M�@r�RQ(��2���UB��Mu^��J+��W�y�!u����#ik��Ռ�tX����[�����Dl���._V���>uB���pA�\��}�Im�L�ݢ~n���!:
!d�|qf/�FC�Faι��� �~��Mg�`�|z^��*�w;���No��D"���#�W��?�y��w,q���� ��ɋ�7b|���t3�?���e����x��B�+|G��Ћ$��sP���5�1O@�J�s�qw.������g�����p����~`sQ��E���Z���	��^��.���j1���e!��qh7�Q_r�ףN�T��(��f�Đ/���ֱ̜��?��%K[�&L���Ի�"	<+� ���%s��<V��nOV3�o�0��>���-��w�����8��P{m�|\��1��;�p>JZ)Tޜ>�z��q��f��a��7�Y4Z��W���KH��S�Eb�8���?� ��$U�|�Ժ52p^��S&�{N�F���֜��ߞ����{�|5�su73����X�'�@�@q`��W�w7�������w/'�{�k�n9/i�eH�W�F�`��S�-~��&�ܕTtEm��#G�k�eC�i,��`AѯW�����4�8A�ZW3�������*$u�\��<��Z�b��N?XV���/;Fn3���x2N�.�>����=W�(̀���ja�%�^��(wi��a.��,H_pZ���uYQi)}ǣ� �?|��Eȵ��.l��xq�R#,�tMn|?	C7�
tX���d�d�����N�2�t�׬҆���Z�Ⱥ���,��w�.5���gw��:d�Uz��snFG����_&9�в�1$UK3�#o[+���x���#
[gą����%�'c&@����7?�]�7?	T�p]6���y�0�.3']j�����V�EM�8��G��u_���8����?�+�-�"Q����w*�8Y�V��1�Iv\2�[o+~���;�� �h���Z"ER籲�B�])p�aa�VtG�#�x�'��W�&�wm�������5�	��1�:sf�LR��T8C������!�B}��O���7B#תQf�Zdy�O���[#��n�ṦMSe��[�{Ηdwj�	���Ȏ��,!���#�/�x����_�h���4׹��L�/g���p��Py��f@p۫�W'z �%@�8�ؔ�9ѩ!0���_�^ILn���p��*Sv�e/�?P�⩨y�����o��ES�Z���[��c��<5�o�TCT���a��׵Cv�z1��o�|�3�|w��@�bq��Ի�Ģb�i6UldP1$�_k�y���x���Ty��Ϗ��i�[c����l_��wQ�۹)��Mv2�79Ԫ^3�z�"��K���3�:����vc=�p�B�AJouD�(IIy����	�<�7u{8Эk��{���U�aw3=����ؘ��~E� ��y�BCar/������El��%��x��q�-,��eF8,��S�v�����ӧo��M�K_	-g��*+~�X`fZ� �]g7	�/K�<˗�0 +�Xik�%p5M�ou��jYE	�^�v҇�[l7���N��)mPV� �'�V&J(�c�Pw�;0U�Ev�H�;|���:'¯�s-P�5�y>�ye����!HI���^�k��a/�`��[�s�T������*=Ǡ=h��,�hv:���!�*�w`qz#��i$�_&�d���,��nQD3��O2��U��F�.ݦ竏FŪS��q�"u@Do�x�n�ĭq,��'2p��Z�SdG�W[ѥ��̱>�Q��X-���5� �BşjwJ�\��綑ߚ��G�e�mp9��iq��Fn0�Zژ��Zi�8"f���o�Ӵ�K���� ���_����$�vA�o���o�${_U]����q>/���N�IγXV�*ը����tM�����(ko��*�_ѕ-?�揇c1=\��mg�a�&�m�33U�+5�Y���R�މH7�u�%����uN�ɣ&�z]��������j��Ha}ws$���El�-���)d�(�%��q11�!�U��M�7�"
���>�8���tv��y
:�aP���h�J�z]�U󋒜g��CA������6�@Po9}4�k�}ҹ^�K�v�����ٵx�CȾ���<E'��5�;��,�/��`b�/߶6�_G�?͔f�T�2��+\+c�R�M1�V���l�y�Σ�����僭`ۘBb�|tЊ�^���U�'<�fi4�{t\��^�x���t\&7C�"��7�pr�z+�����TS(��3v\3��w��S�&�	�0� "2u#ye�?��݃D����l���f��o3+J�,mKǏ9dy��5��2y\��6��h�<�K�	D�	U�ꛔg�␬�����iBu&m���e�E8z/���)KX��${�E�����2kq���t@^#(j���;<�1���K�4*�1tQ���虓�|<f��y���77�6ܶ^����I��E�ٽ��4�?�w�P��}�C�m3;���@���a���8se@��j�A
����:�� o�J�4��iY��^�2�u���v�f��� ��tˑ%����I1k�����c]���uؗ�������R�1K�gL�'�Q�#��YdрVE�κ����� c{l���������܃m�V0h�ƟD���(�p�Z��O�!?W+�U�\g;�Ƴ�$�0D�'H+|�,mPu�5��)H���t=R���T�K�����?�H�MLa����Em�m�@H"����_Rg,�/�#������_3f $��F���]��l-N�a*>����Z&�;m?�WPci1�7i�ҋ%ï��q�&�Y��AKm�th�ޔ��:9��r'_K�v���W�Ή j�kdZ�?bU�QO�5#>�YG�$�����	�FXɉ��tCŇef(�x	�fP$������I��V�o�'^~o�ѡ6�"�a�4���=��]2=ᆂ�jQ"����E{"�����	���,ʄw�/X.
]��O�QQ<��t����i�,\�����d>�}Y�b�8�;#�J0R�T�������FY��;����Խ��#c���rm�}�G�NOY��Y���z�k+G�|?%�Ϊ�ǭ
م�"<Z)�v���Ԭ�c������B�n_�=[T?���N$�1�7b��D��q���i�uu�z�8ُ�:U�g��0j"�{�w�� 3�n!d(-_�^��50;���7�Z��2)���#l�B񍡎ѵ]�	@��s=��5	]7���<��\#B����A-N�:���ʬEb�ud:js�N|Us:R~��)�&��4iF*l�?�[d`���d�<_:s���m�`�o��j��X�z�T�����9�N�!�εna���8�Kz*,�R��9��/�&�x_�x"O�y����{����0nV�/����*oFW��A��(����d]���'
9�Db7��-#p����d4�>0s ��?��:(��އ��i7��>	x����[ �	 � Y�)���t�'�F���X\������,��������{G�W�D����D�OS��ۥ�J��U��IY��}�@�|'_��,�|���?X �;�����-�ll_�M��$"�:��%�B���1M0J��=��,��°KP�>>�:�`:AH�����Khu]Po���dt��Q$o�hq��.8RH�|���a:6�7W��ڿcT��/�7)���� �7�^;�&��� �c�e�����R�c��c3q���{��k����+����;U����l�%��C�`�̫՟�#����5�4E�y������Ɔ�$�p��t224�t�~g��j*��[�N����J��⤿�Yc�`?���V����a�}��KH�gkx�$8�E�{b?����*��W�@ ���.�W��H�Ъ�.��^��� �F�|���T����}�ԭ0=0�/A�^�6:��W<d�c���K���i	�-��%�^��_�=q��AgVA�>��T�BP�����A��֬ōo79mh@�ߤϒb�*�����魹FΛ�s��H��%p�!f��*������[�JY��qE�Ec"��C	���Q�ɬ`M%������|�~$^��A���i��b8�J�}dd�
0��KI��v
�h��gJ�ep���ֳ���E3�����;�Ҥu���z@�\��py!��x��{F�D���J'vo,���4��#L۾s�e�M���y"�d��6��m!��.*@P�r�If8�gʴ���D|u�rvw��l3�B)A^��&4)h���&���?S�r^F�4G��B��-�T������7~�A�B�MAfa�����������>���g_�֯(�M�S3�B?7�6�-S��>�]� &Pg�M^�(�(&�r�hL4������ȗz5��M��l�w2!�Ҭ��j�!���ԅ����."6�џ�Ru���@K�՝Պ4(���5���86���}�lL�"�d+q)�4��c�����qU�7�g��t8	tO��:'\!�ڻˎ����Uu�a��,�1�۲)��F��yHc3���xsA�����Y�y�{�)�����W�ڌ���U+t�|�������(�%^:J��#*��y�>�u��ҿ���%��H��_7}`�=)�9�/w�j� �-3�mQ�}�s�{���;�cfGS��,��K>'6E�MpҜ��@r���;���(��ғB>r%Ɇ*��}޷�[M��Ő?��0=�
'���kT�*�
Ni�ppr��[v��b�$>�$��g.�z+'$�j�j$,��ֳ`� �f�C�������'�O�Fi���Z3�qsq���)�G�]ے��HO �w�VΠ?&;�@1o��'�2�G:���Y�Z��'9���XQ�:����2OƓ�&=�>�^��l���C&�Ԣ��w��� �����~�{��b4aTC�T��b��@]�����z;`6����k��¬ޱ1�50�"ܔ��C]�u��03�v�5*�jd�jβ�̻�};��t¸�ǾK�C�W���������9��t����d��1�����k�~�s`�ƙ�@v<h��k�M��yFP<��,G{�L�ب� �y��=�.�¾�]}�my
�k^߽�C��5eQ�za�b���k&Sȅ~n��s>ز�
�y�d]�=s8q=[r'���@�g��pUK7hsi�=]^����t���R[��bh��������Ǝ�i_�my`,��j&�|G��}�������\Y�Q�*�a��	I�q�l��'������fC��X<Ǘ�	�ο�d�U�/k/kr��-���X�M�	Oz�n��4x�$.��P���Y���2�*�L`&�sЀ~��=��mA:�Oi���L�0ˠ4W��ؗ�����@et�ֹY75r��+����v������I_/v������{��|1s?�OX�H>o[M�G���T�Rah����1�-gC>��h;�d�K��̥��f��LF�eu���#RU.߆ �E���y���
q�L�1����x���˳|f�¾%�B_3O�FR�	����S�:�'��E��q���MI���`�A���Y�,�57G�6O5m��;�sE�ո�4��e���DQ�3��LM5��a',W�-����ƈ.��>��ȹ����u��yĂ���o�c��(���Ga��f�z�"o��G����CF�|�w�[� JG?ol�����.D_�fZ|�鴓<?�2"�E9@����<fG)�l���2�!��25%�r}i�0��v�x�&f�~��� l��%��6�]��N�%s2�goYT����}�	1��kWz����I��������&E+��6�w'H@��b�F&�Ւ\�튥��ЍW���(DP`&��
�ۈZ��S3K�<�KLBgV��V"|V��냺
�[4��r,A�f���׌�3��]'*�1�Z훍ua�׫�Gt8��S�����\Of)~��ׁFӝ�Z��:Z#9j2 �@b�(c!��{�X��jx��Mv�(G���>vbWǜ��s#����ؠ���r��9[\�N���`��t��?:�+XQ(���cI�p[ƀ��;�<���HZHgO��`��4�o$�/�*��r+wfE�D�3�!��p�7h����u܍�IL/�<*M�\�k�	Oߵ��$Z�
�&+�Cf"#=L*$T�!n�,l�e4�8�d�L��͛sO��F5�>�0�|�|�� ]��v����~w���{���D���$�v#'��F_����l��3��t���Ȫ�5��9�i ��[^�=4�M��#v��  �<Og���4��Gs��
H�ˁQRK`Խy�������S��["���wT�m�^��>LaMH�Ev$5�> +���x�� �
:���/���a�UC� �`�UW[�O����>6�\���M�$T8���� ߄4'�h�iՐݸ�ރ�bJ��kp�L��#�~���4�P_K���xe�?84�����]�k�c����My1"��H=&5i��+�e��RR��H���CR*G���Ί�"��+����'�ȋ�������0k�_�:d��qb�$�y%⑥=Â�.��0O�ycl�?XV%3����>��||�^��8��0qC�����H"�t���r�Mۓ�jt��J���3���됼�A��!�uM�B�(+C��_���K2���\_ٽ(���X@��b��������!�kL%Pjq���E7*������Cd9j�{n|��߮��QuUY�5oF/�� F�<r�˶��i)�u��h�;0_]��y�e�L#�M�>�&�/�4��k�q� �z��$��ÉLh���2"�2�Ű����gQ7����� �����e0O�흕3k�>�?�ϱ�}�R�/���8Pxj����4y�C�3t�}%ʹE��Ջ;3��/�T1��,��]2�k:ˡd��f��Dr:����F� �%K�rZ{/]��`R�d�+ݣwQ�ʣ�G+���������VY��E�H[�]2"�a#S�W*7z��/�v��{�d�ˏK���xh�E��9�AQ������β(��3MM
��[{�(@����1)¾�	3f[����U�|M
&�w4æ�X{վ�M,|���n���A m;�,�轸��A$k�!E�`�#ě�@�o	c3\g�wL���fZ5��-�P��kjMOLY��|�WH�u\)���^�=�¡,�p*��ۀ�8w�O*�X�Z$`���mz�p�|+���ԗj`7	�lR#����ҏ}�W���j���i7ة��*<��J�M9\��S��?s�`��$��|�S�����rR1�����r6�w�jƝg�����!���O.h:����L���v5�{3�>��f��ƶQ��>��	 e��_����?f���n��Zm0�^⡯��#��mE!Ŕ���Z���ϊ	�`M��đ�Y�g���X�B)n��?��%�Jp����ͦk����Y[=����*x��Ǭ�g�l����+ܔ�m�Z5��1�^���`e�ѷ���?8���/?�x4N:����d�#�HM��i�D�����@80�VB������Ή�GYv�%1C���>��~8xL��_\Ei���,W���Ɉ�Zv���Q��u4�Rj�lW��Y�)�G�����J�B>��`?N;�^�e����wM����ֈ �F>l�Ђ�ɟ@�{UP�s�AL}*J���W���R������>�sՂ��U3E-����{R�����!̀����o㙌��������1�����H��-����諦uX�:p�8^��١>8�L��;&@WF�@2�l�u*��3NUX�b(�I���2���)��{���:>7��q�	B���ŷ�l݇qH�q��g�N)͙�0e��q �[�;M~Mx�}�	����'����|>��s]�C��	v��48��<�M��T)�/�Bս!5�~ċ�DJgSAp�\_k��+�J.�UX�A�`�H6��#)$��ӽE��IL�H�<������� ��H$��Rce�/;��pg��"�!���A]��y�y_�����h����h�����x$;�f3�F�q{k�Zw��}'�f��嗝`IqD�:K��M<d(�ǖ_P��6��L�K���sb����DG�8��<�{΀���)��.%s@R(�8�j�$��TT��0xj�����.d;7C`P.I�>fW�t,!7tG�g�����̕��%k��y�GM�`�R�dB��[������|�}��&nF���	Q�>�
���G� [���k[�]�a�v��l�~Sw�ۃ!��ֶ%7¤�UBo��Q1^��^���܇_���"���\��������ڮA��b���}@�g�����|�����W�@�=����q1u��u����'�u4�ң�o�$g���M�9�p��X���T�Iݛ�ӈ�L�$�JB>����!�n�����p���䵓nrV8�I)���{4s05�WC4FQ�1�]�H��Z�^㷮<I]+C��!_4� ��ǫ
�n�(�`I�}7��k����u5���rZ�(Cq'�:��gï�MZ��`��k���5 h��+�,��!���_@Җ��+I��!��H-1�xdӂ�7��3�K߽���c՝t6򆻘��^��D�]�]�z����'��"f�B>sl�󮫥��Bk���ב�i���U��Ԗ�<&)]��][����F��P�q�'fF�yX��(�ޒ�t�l[�"�k=WF��<K��U�V�E�,��L6E�x�n�ӒLI~����'؄�\�P�Ul���ڤ[ti��)mZ�1��=>0Yy�<�B;e٥E�95�� f>�ަ=|x�h�A�,o~ݒ���h��OA�� ������zE{��� J���*r�sg���&W��O�MU�+�'���	ڢ�ы����k_2�#rS�m��o��tC�z�(V>���uW�O�=��:���� �@L8��8���#`|��A-�f<���=$���5���	ĭ���f��~��JE�&@8���rd��jL�X��lW�É295��{<���:mk����:�V����%ɣ�u��r.iF�Rn�d& ���J�hi28��h���_�z���s��K�;IJ|]�N����Tb�8�k�9f��Ȕ��';B��i�X7�/l��r�oV��R���+�X��U�g8�-�H��F�%%�h:��O�Ǖ,`���)�<���Ps"(��h��؈�m���x����{���\�� ?��I;&����I��A�؍�b$�	��cp����5C/	[�\�&<�I1������DZ�3� j�?��]2B�'��u	���j���'i�zu��<�4
�y�x,Y���X��r�� ē���7�zb� � V=�����P9гH�hk��P�4��R��Z*9��=��0�v���D�.X^!�Qʹ��qj.m�8�m�]���	�V��V��'��h��-�\��aW�&
p�m
�֭D��ym�mu�~
M�n�aӭk1�־���V���z��c�SB���;�]�z��/j����;@�d�*���/d����h{8�\<� ����/�V��J?�#ow�oqO�������|� [�9��M��^�}d^��h�&T�Xi��;~𧅍p��Q������`(TT�8��A���v��i)@7΅�������vz����`��m������%��o�>㿾D?|l��u"�r����Al�L (iJ�g&�o���i��7�|��s�<������d���� ���9/9��ЁU-���(����w�j��U1���cz��@й6�Rn�ev.����֐�'�vؿ��1f��i��h�^L�=�Qs>�԰Q@�y7����	S�5���L���TG�/�7����gۥ�	���0�u��мE(���G�3�yn�7)'�����㊏x�����;��T\���t{İ|��O���'�U�t�ݒ��0��jo��cY�g���(cvGx)�<ǯtO��B�^�$���[�T�T��۶e�����8���)n��}��!��{ϥx[��1S����mN�S�{zA�y:�TWq�r;���&c�VE(�|�ZM�3+�c�����7E�8��=�C����@�ڼ����E�)�Tu�]�U�O}F9��Mr����g
Bv����Fq8щl�R6�oQ6���������yA��t<���D9�c
I#l���;��m6w!:�L�Q������
�>gwc;◆qF�9���NV�ݏ$*ld�Sq��ci�̔ {�U���������>����]�3�.O��v�����qTG�B��*�o�&�4��i^h� !=y���}�GJX�?2�7���%�Lq�m�wA�XI���/��TSs��>���"1z����4v����e MW����q'#��b�vjZ�$�3�&q4�p�un�uBD�re�V��.6�sl��%��ʑ���%cO�(���kJ�E
����|����L�0��7����x�\5�0���̿�����O�)[v�4�s&>%�*�Aˬ�󖺅J[w"K�?0va����{���|x�S�̖�O���K�+Eӊ;�^<�ʷ /"x��Y�f��[����/l����m$��i[����CK���.H��}/R� �O�;)�Eo����.`�Vم��4�͈_q��5��`������>�[�qQ��Lq�/���J��Z(�KL�#�<�m�w�87Z3��N�`Igx]nPtpaH�z}@�rn��:A,H�b1ڕ�\��8ϿܽP���x��Uoa4)��F������O�_@�Mȱ����D�T,���C7<ځtD_m�ݼ��$*t9_Byr�Y#
�������v۴&c���̣��Sc�z��K��� �*�G�j!��P�� T�����M�M5{����2���bX_�'9��������τ�xO�h͂P(���A����� ���r
(�s8<���F7�C�	���z�.�µ �(�SQ.٭��m��Sy��pOA���
���&^x��ڑ<u���[C\��q����@E���� �gN.,�=!��y+�TV�B�y.���c3��ǋ[͠x���;���,(�,y�*���VPf(���<$��[	��]��uՂ7��)�29��|J�u��Ԣ�i�s ��C��z��D!6��[NZc��qvကX�}4-�'��ͪԀ�z^ ������:2���Ȫ��w�k18��1`�[�:G�!T0p7%�a��Nu�t5������ߵO��tP\���1�Ϟ�Qk���׮�ɠQ+�5�R�#:0#��l�0��7�C����?�t�� aM:CسJ!R�E@�!u?$gk�������:��z����!����kE�pTꄋ����̇�ccG�BR��Ȣ�Tű�MA%Y�k����.^�����!��"�X���e�Kg�Y"��o�AY���dE!2�A5��	��!��p��_8@>l�#�-A nh���TTJ���3;)��^��&[��9����G��2��M�O�9J�Z�O����ن^.�;jy�����ÿ	Ep�%�'���R���0��ŔB��&9�x��i�H	ה��zTL�T���`�:^�]�I�s�sKc��*�����Vz^/z�O�	��{����ҧ�E$MÒ�H3��������<;/���~�j�'��+fE��U>D\�m����}��0Sq������̊Z�ϱ�%д؉o層��x���&��evLY,�N��ҥK>��O������2�xb����UN\��҈YMu�� �|&,Z�PY�f	��y�z�Q�v ϧ���6��}��<&��*M�{�o�`�K�<Ox3�����-܌$l3#�s���N��O>
'��.�1�y*Kr����ܫ�3��l�MCG\�/>2"-jB��|�!�k����I�\����OCϐ]H� H� Zܰ�o�Ǩ|\�scWw�P?��ќ��J"dQ�/5A���
�RBzd� ��ŷ����A�m@zZsyᱶk�e�4�s2 	OE}ʣ �2�0;��[/�[�Q�H�m^q�A�j0D_2�l,<�g$p�;����P�Or꥗����[FiH2�'
�;Y��޹�S��wȶ:���w��?Հ�!R�'�)V����,�����q��˲�.��(:�۷q�u�(�w@�.���3~i؝��Dy�7]˔��zm��^�4��E�BD�{�V/����3����ʆ�V��B�Ir��-W���$��Qړ�`m(%���{$~�I�3�+K��E�.
;�T�}d\ˮ�����H�(JɜV�c���d�Ck#l�|;��|2/tv��[H����y��� Y�9֫�\������P<�ߐb?�T��ʦ�z�#���c/lFO:ʝ�)xp��6�r��=8M�"��Y��B[wBI�d��!r��4�j�Ĺ6H���垣Ѝ�a�c�c.���T�d�jY(��%b�>�*��C��&�{���	�P�q&M�oJ�RzW����W��0Ęh L��8��j�:(P"<OL���n��4omٓ��l�o���U�
��+�򼦭���	���Й��b(����޵���~��W&)IS����od��Ҹ<~ � R�(ϊzCYQ��z�&�t]����"=�@6Ϯ!�#���Z�7�W�j�Yf?�Uz�Ś[GO��Z��o�(C���|g��E*�����]s�J4����ixĚ+�䎖!c��k�W����G�| L|3G�>��WC����:'���m�u���V&�zJ���gҳ�&���tY��r�5ߜ.�)f���<+�9��J<����p� $���5}��n��U���J�=�6��k��{�����h�0P��2�2����'u��-"bLT���4^t�\Ѓ�Ӷ,��f����Œx<���V�ɨ����3�4̿^s�i�!���\!�.���:Z�+Y���︲z�F�8�;Y���>�� }���Z�5nS[�Ƕ
�""{���6Gxt��q��on��Vn^������^��drRW�ݘjz:�G
��u�C�O.�$z�`����
ʪJ�\sY�Ov�́D���	 �{{(����O)�Q�e��遪6qف͝�hrUٺ���6�k.^Ai�k���u���I1~�1��%/_���܄������&�qKhWޅU�~m�{�V�jA�ʊM����X���'�ӈ�H�pS�-|��J� �
7��*�%��S�wq�uL .�0��n��t��6.�� �&c��m���U2s�'�MB]��)�Y�Wo]�N}Bj�X�)��_�̩�5�`�%Ǽ���U���:���:��f�Թ�NVQ[U��aQ7�8������N�ل���R>����[��X�w4���m^����Q��Ȓg�ح ��v=o���9.Oy��e�Bc��5mb�Hb+�+��K�]s�M,�}g�j�f�`x�&ќ`��U��|�ft�y,u8V��А�ʎ!k��8�?�(�)�I= Ө���^� Ly�����$0@^�+�0Kͧ�r�ʖLv[�����n�k��d��������O:�k��.E��-3��޺��X��w��5�@�,�o�պ02�����a0J��=B� �L�)�2l�
e낁�u���|H��#��2%7��4���Xlvz��b�i��L����S��1&�K���J{���Ψ�F$}*1k}"����e|��6�E��2(�R�l�6�7y8�s�w<~����0���AC�m�jQ{�1�����nx����$��^it��}����-�2-�q��s�'c�o	�A��v�6�4D��Y�Kȝ��	�"dŋc�-'d������K�(h7e+�!T�2�tU��\{�/����p�f���~~��51튩��^�hCy��и��cC�����oy�mr/�w��փ��!V^�2��߯)�f4�vf��4@�ţ�f�9�C8,`�G"��A 
�Kz.I�!Y����]��5(C��⹱���B}Æ_�&�<]0t�W���v�*�_�Qz����z�A6B�Hh���xǃ�F�Q2���7u1h�r�u�QxG�jb��I	/at�l2�h�wVE!���c��s��<9 ����/�p):���Ȼm��ʌ�@���N� ��M��yx����:�.|�K�|���>�eB���6��yn�Q�]E�\
v�c?����ܫ HP�Y� ����l0�HQNi!9�1�φX�\�&!�s���}�� ~�ԝ ��&��[���$�g�f5Q�S�l���Ϙ�h�x���,�}���ت󌳖e����e��~2���Ap!vKw��1 >y9'ӥ{&��c:��1�W��`�� 8��iV������F�ne���*��"@9�#(�n'��c��}�B�Nq��s�	A	!���̑oÐV�T]��3m���l~�̹c#d���.����2�b�.�� �=�k��n�m�I��w+oz� n��v�U�,��@����8B�CУV���H,N>K��g֍���:�e����`1-&��cD����U�����}���>9�� 6c"]Fe�L�.�'S�.�d��׫B�˫���X,	{c��mo§���'�%�BZ�~���|r 9ے0MLk����(=Nk�S) TV_����Nρ����S�}st��3�ڌ����Z{7|�mQW"u��zQN픕���y=�43�d�}i�@�cB�]��v 2 ���5��Y}�}U�6���FQ_�s�'K��4�rV9��p�7vp>��[���<!>�R�:�>��FBފ*ȶ�x���{V�6>9�՟�Z,W��<��IQ���R ]���7�zH�ˉm�F	��2���k�]7YY�@F��N˳1́�%���UQD�k��a��ϼ� �SgbD�C�nhnri��S��T������t\�a�����0���5
G��U�y��^5��Y'��9	���v˸Ȁ] P>���{�� �p���lwh1h�'f� �pH�e�
������H�m�FPL:1�e�ڳ���=o��@�,��栴��R�UC���证�}��&��,$��B�uED�������߂��B�*��b+����9U��+p�3T����0iCT�����,$퍂s���5�T�tː����Yd��=�IՏ���״���]9A=L��ʉE:u�t��UH^B6|DV�B����/�~i��$)7~ZEBTvi���ӹ!�
h�>)9�R0'�>���V�H�S�����
� �]>ь}��_ �X� X�>��Yi��3<gae�?�\�,-N��b�S!���̓��4g�ٴee�,]� P�"Ñ� ���1s-�QHj��v��<O�~YC@�l���UCr�(��^� ��k����0����Mq(��ls����sP)!��c���9�^K(�l����2FX	��S`2P�%���w��Z�1�9�F[��32�=Hlnb���x>�j0�0�yRWz%�����5�����:1/[w��~�e�}a�.�Td��Yn�T��s3)z4$k��YYq��ZZ�d3����{�w�Ǳ��Z/�r�IU��Hy\3�p]vQ�E���Dh�.k��[w��z��1l���:���=�.��G���qR���8ĕ�y
\���u)�8R�עq����r��#�r.�<\� {�4L���;���;mj�ާ�TZ�`�����d/� k�Cߑ��b�h~��o)��(����>���"�\�cc��_Q�~�щ|\�qʞ�ww�!���I@��X�hL�����u@k������������h�0
�W7���9}t�A�+n>��#�s���KY�FԖP�����(�dZ��a���X?Ec86s�����|k����y-F���w#��w5�r�4A�9\�CLn�#��
7|�3v�p�.@�%~��Lx�H�7��{������{g�W��u7�S�ܖ�7=��7>��*�7
/J��}�%���RĿ�Wo����N�ro�v\�q������uԗ@��=�b*�g���(hT��?����.A��_����%�`CQ��q�N�AK熌�����-�ʁ�%�F������gy�t��$���~&\��g���(�jʳ^-Æ��L����-��d��di;_i�v`:�&B�Ц)��>r�L�����������٣�r���aB_QS��f�}F6�v�s'�'���+h��Ӟs*�$İw�!�!�cP4���qD���ٍ�*�<F�����!���Q-5�2�?���IYڽ�.����?��lS���>��[�]Y�/�O��І}��>���5�l��D���%+ G+`l�+MFa�Y���U2A�t��#�^��p�`@����Z9 _�3Y*��n����%����T��&�ݴ��E[�i���G��Y��N~Q�t8�h���~2�;u���a�e�c�bM{����l(�S��Ro�a*���k|�O�o��(m�Z�#�Q��Rҵ����8�u,�ƣ�W��&�&�:�"՟��8�gքz�-z�I��XP�*��lj��������mq�<0~�LWS�f@愯R���U�Ay�"I9l���+�z�WU�$pS��N����f	GV#�?&�[B�*�����UpI�Η�p� ��$H���\EBhD��u K�|�,>DR��XeY���1���ݕG��]�Ұk��ahռ)Y�M���I,��~�ʯ���}{�-o6ڣ
Gb�
����i�t\4Sh@5�/��e@O��U��u����� Of4|�?w�S*���1�;�7�4n��¥LV~�r����z�����M�·'�Ey���������!Y�^��eM{�;T�QP��w�#���H��ԑiA) %w�'m��}�
k������նr�qA��1^6�W��Z�ˏf�����h�3�1� mN3(_�K{^�7+����3���*��|n�mi-*�<�t�n-c��x����`�4�O�)����R�1<0�0A�]���<�x�yC���K �{�M>��-5i�q>jK;����J�5�����J���l/3�ebo�'o�d)^
��,���{�ԲL���ըC��!�f=�B$_C���X���! �� �w\2�ݕeMPL>�>���;r�w��V��n|�<�P7�wBYL�3W� �����-LٳC�����l9,�wv2���!�x~ZgJ����q���p������VW�:�M�V8,3�>��Qe�10����N�w�ي�ߓݑ+�����nX	y�kۼÛA�$cZ�f�s��a��}C�1 ?f܊M��g�mV�K�y�B�2��Ć��F�~�~t9�JE�ЙF�m.�a���{�H�[z��l�[�=b=c��S�6�Rؕ�#�n�<O96�
W}��z�,Y����5��Žӳ^ih���,E�y���q>'�B/�lT���5/�孬K�d�R;.����O>�N�}e�5H�Si���f:�y�eї���5�S7Wo;(n��=�S�xj�n�(�P���n9_,�E�t>�m�ӹX�'�9�'��-�_�f=
�FI�@��L� A�Z�W�nt��[�x!]���̇o�4#^��4�����I��Ɔ�4{=v�<H����3��F��o^������w\��h���/�L���^��/Q=̆�M5N��D*+41�h[����
��&������k.Oa�՚/L0��b1	Q��HN�X5bm��?0���T�M^�k\;�h���`�1sN�n�¡�̌ynh6�Y N�72�;ٖ��ձN�>���c�3���%+�ի���zX�b����%�� ��&���t˭�4�J�d�8m��"s���!EHp�����k� jr�;��I�S��wù�$�ϭ�r_Jdl�De�po��vw��ϴ;0i��w�x�o�����kB+�y<]!���H�sS�PJ!��'_Ֆ?)/�(GGY�&��q@
�	�`��;ż��(h��'��"�5;�7�8�q�9<@��F�)��P(]%�h����&5�}1z���=z�zڵw���~�G��0ld����R�Uʛ��׆7�[W���ؒڏ�.�tH�lc"6-��0�Gx����.�:Nɵ�6���s�\�W%y�l�� �_�g_���c1J��~���1�=���j��;b�"�䑀Ă��D �ҁ��Y�N�����p�wB_�����R���\zl�Zx���,�͙�	4�%B��Xf�Ag�$�s�+�"�U��qU���7�64̑����y�p~�`���e��u�Yw����.8C�0b�+�:�9w�FzJ���.�.����N���r���uW?�X-�Z8c�������0� ]�B�cpw�?�h��"��Β4��~]�S϶~wU�ŀ�g�F��;�L�<�Ի��b�̨���`/"��h�S�妩��S]����*�H:?'�s�� /��ޅ�pfЈ�G܌�M��lG�������۲�\+���w~B E�ga/�_:�ZK��n�����<�s]�%�����H���mN �r����_�,�9f� �ia��QW1ԼQ��$u���cY��&�Y���)$y@��Rl@
�X�	�j�� �'j�8�#�<p Y?4�Px]�s�	��\��J�������R��pỴ���N�%�ݰ^���i���AHy�����l�V�����t �U]��S�V[4�����|��m�$���zF���8�0��+����u�����&CmFS��w�i�h �,���]��������E��*6����S2���N1�q���P�
S�����~z���䟨Փ�@	��ɳt��4WS�-(ìP�!��̟�C��!�(tںJAȲ!��ۯ�?�Xq3J�4�x+8��b^��	?r�"�9�ޛ�$y	6�W�@�����}�����6�?����|?d:���0M��H=N�Uu�ܟ�qϪ��G�	m?-��|F��+��
L��7�E��0��tB�TdDO�*ȷ����>�󲠅��c�O����)gD�;��_W�������: �1[B��# |X�];PhLR�&��uv�*l�3����C}qeY��}�=�2�-�;�X��[�vv���n��	��{&̜��λ�Nw�xq�y���z��";ДC��Ov^�e�2r��m�Ё�����D+2��,�&.���X�LcS��h��O� ��4��Ue����b�uCT1C�^-�ҳ�.՘K�S�'�S䵡j|Oԧ�A�`-��xt�����~���׳���?1�i�o�'w�3β��kSCe�+��î7 A&j�<"�#I��xJj�M��H`ڢ([ {��2	�S��J��Q,��@�¡Y���:x��0��M*�kH�n�1��c�A�q��v��j87"�p>�p&'}0����*�����ȃ��	��++-]/h�;���3J�%�@�����w�����TxDn�?и6N�ϗ��s����GD|/�����X1[����F���Vk�uTxt~7mQ�ք%����v�P�? *��2���KZR��:���<]N�^�0�&����.�N�9�&V�zE����7\�. �I3t�9�\�:4E
qͮ4&Ē���|���۶ry����Z%����̛M�)g�L�����J�Om%Q�)�6�ã��4!�|*��`��j$�<Y�ޖȣ�.�؛�J҄=FixU�T�Qؗ�P�FU��P�sP;�?�zL>�CW�}9t���}Ú���7\��>��Qz\���F�ؾco���H��L���+�%��#/A|�R�l=��]+x?Y5�1\�����L&���,#���y���I�g�;���|�:��F�*2��P�7w�.�eag �u��S`�U�ş�R'��$�0eo��U�Pq#�xi�DrE�����!�ܽ��Y�)�#8N(~��:��h�II���FI���q� TQ� s5c���I��
(Yحn��G��bF.�;
C�İ�ʰ��p�����;�m �2PP�e������)e��,8�� X#��z�h�J�$�:��R.�7>��k�kj�o����$ �ʓφ�J�J�d���y�m�UV��C�����>t�s��S��}<�Ϲ.��Jf�J{n��W�k�ׇ��;�:u����&|��;�,E8�M���$�!�R�~@���@����<�mf��axh��.&���{d3�N�=h�4�e׈2S��y�~z�
��R�ꍙ���T:b_�ȟ�1��P�=C��w&�mN@|BJvR�N�*��QQEDH}��m@|ϔ�髐 F��ChdC�:X������K������D��D[v��<NǗ8��X�H�QZF_���g��Z���ks�o��Jн�Q�����oJU0���G���ĉ��ө���"���n@슥��_��_�M�yn��
Sp�[�j-@�X�80�a�7�$Ƴh�����딗��=��~���W^��{�AV><m���c���䊒�qfݬ5��ʣ����6!�/�$�zq�J�tve�3��e�X��\��=2!آKR󏆉� 黑1D�{{1}Z�nw�Y�D9@��e�^K�@���� <�
� �7R=����64�I�)Әc�]�X9����A�" SC�ntBIP0����Pu�&L�ӿ^]l�7a5E��28U�HI�P�;A-֓��1oA���ᒤ5�R���Zb���"�u�f�߃��]��^����ܬ��ڢ玶������:C��zJ[�9��p�湵u33��:�����#��&������̊��5�����FQu?�Z�5W-!�iQ�ZL���]�c�˓%�>Â��|)rŇ${g,�o���>�@]�4��\7���J��T�
��SE��;�6����Rkd���:�ڝ�w6�Sp���7K8�:�,ͻͯ ̢3��f'�
��*
]�!dJcR�O>�!��
em�%=DHYV
c�x*���I��2�'���1�YN�@����z嵑7Y�d2�19�KΘ��ț�����|�@�R�6a!G]��Mb�h���(^�6���{�[ׁ�I��6c>�7с��	��uW�$m�ί�"mk�Xk�ǝ�=�H�~��1��#���:u��ʢ�d▄�B��Wrc2$&��rpd9�� �6�m�i#�4��t�#�K�C`=TE�^R����7 GvL��^{����MR�(�����&T!�kPz�H��f)S�!`������u��~�3Pqy|��"��`A��[���ڡ��+��kO�h	����ۢ�䎠�t�I���d����˹���KQeVu��O��):$�σpv�om�a����P��W�_w�`��0"��+�m�|����{l�(��>D(
i�T�Փr�Bf�PW�vk�p"��$�6�W�*��s�k_)R�3�%���μui*��S���K�u!���}
�\�L��:Kf��q�[��MQ����&�xtF'	4w[��R�N��j�c�l6o�LV���R����?�Y+��:�8�YW{�$3����G���5)�>[��'8��;�7A �·OUu�b	�G�g~]�K��V���}g]�Kz�y&#�eȚ��B�����Y�,�kBNJ����xT�����r+���Ee��B�y1W��)���Sχ݌�d��.����A)�-����V���{������ѯY]<��N�������!�׷��b"S5�q2��;�q��W<�X�Av�^N�e�#\N�n�nͰA�(]�Nnqx�t>�����rP��<��ߣ� H��;�ȼ eٸ}��vo%] A-�H���1��7�I�h0(�s��=���%=����*�w=��w�0��.��[�uJ��/2&�oI4�<��dn�)YM��7�Oe�T�T`+����2�b��H����X_���<��'$�$)a���e!W�Xj��3�Aj��_� ��5���\B�"﹒2�h{5�R���4��Z�B'BpC�5�'�����iT@�Ȝ%�j���6��lA�h�4	${
xl�H�Cj��Q�oȍ�|�ta��'��<���%�����#~)]�Ǉ��ʄP���!e y����'��E*fu��
����uYm�:	<d���Y�����y)9�b$�/Q$�s��o.܊,g�+���Sᐄ��A`+~/>�
!�`�h���>D�Չ�d��)��B}#��x��4�M�%��B�+͵ǽ�#W�؅T���a�P�������]`!5���|��H�5�._��jH�+]� �3US��
^>�xRz�A�㼝EN��('ә��k��N_�!������ ��q�%R�W��a�lT�����" _~�7�/�����~�`;G�2>m��1ܜg�c���Ǫޭ���V�4�U�a�N��Pe�=�+o`0h��W	�Ǚ�*�\�uE�q܄���^3\qqi�oI�Q���B�j|�EC�;:(bB�ɾ��R�� ? ���yA����^ݝ�IEto���U����&��k�*8)�A�/J�"\2y����p��v�~��ؑY�G�0�B�G��J�,�!���30HF�::\�T���Sζ�2JQ��Zi5��2I�Urc�t����B��eMl�2�$�79S�F�ו�^�vdsY6 uE��*ܜUօe:���Y}M��6\S�����,\$�nQ�Vw(�ݜ��b�?Q�'A���D	W<��R)��}��_�-�z췙AS��4��-^����=��V8��A��)��t�	8�d��S��@�)t��P�������qD�y�D��?
� 4��q�ZE�,�E�a�"H��r8i�(N����$�ĝ� �}�� �V!�2�D��:3��zp��EA�K�(��]��z�r���ΧjC��X�|o22:�Q&�� �ԟBT2��5-<�Z��ǟc}.�8̸��&'@����w�)0�v[���.o)mi;ȳ����Z�e��2��D��T�$�P��Ҁ��_���G_�C$^���7�;���v�RBp�lk��O$hn�~9I��$9f�ʽ�,�.�zq�b^-J���)���<"��ʑ�r(2~c�Aqg.p]��}RɌZ�N�58��"�l���L$�9�i���gkhLDZ�2e�A?�Xb���A�*찈_L��������dY4�s9R&��.�l��b��&v�"Xh8��d;�����A�6G�a~�h�s���-	7��)2'�[5�$HK�9�ț��I�|7�<�/���Q�(���̛p_$ǧw_��[�E�o�l:)��HC2qX���,�L��"ó_� gl-��,p�l�U\ޠ"=ڮ�7l]�v|d�*G+&a`��v�H�z��$h��X/߀y@���ٟ�u�b�Pr����=+�x�����y3gPI�1]G����6ƥ�b^cSܚ7�G�C�ӱ�'jA�;�Ëڙ]��XdΞ2�Fz
zN���z�Wd�V�t�äd=YZFӕ�Ō>)�/ېߜ����ǫ���^N��v�V\��{��8��O�׈sY���#�����R�|����1��VG6(#n:�5y;�ߘ	��13)͛��d��Tk��G�eu���f�a�i���v-��$vBƫ��:��)x�����5�n=$�3�ֽ0��l�(ō�8����.�:��̢x�魅��T��~`_6��1zy��������M�^�����6��l='�*�FL���*�y�n�� �11��J��4�-�F��:&��3�p3�1_�"�gp��|�!�����|L���fB�qFrL�#X�`h�t0^�D����dN?��@+�@��.�h�U���F\a�$7��ӆ��;k���0�Jc~Ie�az�S��a ����� �6G�T�Ձ�sk�ބ��"�٘$=�e�0�)ㆠ� S���1*I�� ��|w��/�X���8 U"U�i�uq�+Hc��9�_Jy!,�	�V]���a����lp����'b�!-8 󪪧��y��F��I��F!�����ݖUF�u�E�N0�c���Z�\�%���?�zؘ���s��kZ�n?��D"���=P1�.4�y�w�"@���������1T%B�����/
�[��B��?���eC^��?��z������W�NT2�J�����:�.��*U��F��RO��Fy��;A�U���K�uX�{��]��6F�ؘ���"*Ɉ��f��Ar[��?��ګ���^��*W���mD-4�7ĂY�-����f ��ۈ��;R 5y�+ ��	�Ӻ����I8��@��
oG��d��dgh��XF�4,SP�;�z��J��=�=o�W|GLcf��*���v�F�NY�vs7�XW"ɤ<3���8R]yMV�����k��v�t'%��wRI���5p�l��0-�ՙ��l^������}�q:�����$<e%��YX�!�G�J�:a��2fk}�'��n�F��y^3���֪KO+GD;�I����nq�D�Ez�a��
&ݸ���|`��_����r�r�f���һ`��#1�/�H�@��ف����������@ɻYg������Öi�2?&83�t��gn@-ڕa�u �!w����F�?��c��[��=G����L128\���%:��0*����T�;����ܓ����0!bS���A7�D�U�j	�o+ێ�����?�0�O%UV;<Dg��0\�'��%ѡ�/P'H^^����h+	�HC�t�D� g+��ϋ�	af4��ċE��!n��'nZ7�d�ox3��F�i��&��Tɻ�4�	���^8@�W�Wu�<\$�GM��:U�HkdYw:�ۻ���RT���uq�>��vy(�IH�qDB�������K�JE�й���MEբ���i�������<rlp�Io���Ũ����K�V�zέG4�s��t>l����̈́l��3�XP�Fv�(�р��pDQ�g���o�Cn�X�A~����pO]��f����w�mZ�I��@ \���Y����@�G��L���R�yR�;��6k�W��v�b[9Țƿ�k��������`湂��e4⪮ʉt����
)��ҏ	(�B׆�K��� 8\�ǻ�c2��a����~���3��X�7���A�+=���^cB������Y��ȍ���R�(9:�ƓH� �	����IX���@,?s��w��X��2}���f&���2���V���RŐb�Yh\J$��y�x��9�q8���`��FUi�]�t3��D������4���/�����g������T;�C/�\�8�������I^?d��cM�-�M[�&�rƃ�̹�;3�E��$J�Y�4��܋��N�,����;�^�D�B��G�����-�D��s�^�>�h��H��ߛ�	:Io"݋�p��K)tm׉p��P(j��~\��גcz��D2�M_��$�5p�@�@]�|=B]gLD@`���[����.F��ȝjr���ȹ���鄨x�$u���H�M; JͶx�w�@W�p]�T��;���\H8S�λv�Gg�3����>�h����VW��'*���ڧYM�y��k�:+{��(1"��l�-�9�Z�6������'>�{�7���h]ȸU
{�L�M����o���!�t[UZ�@�zmn�+n�Qd���EN��Tؒ
�=$���*0�I2(� c�(}j+�I[��߀�ǃ��X����$��YO;�(�#U �G}��U��{��4����k�z�K��y񌄲��j|UJ�P�Re��\��q��>)�<�2�WsC_����Ő7�I��>fDb�����ҠLe���N�ε;@8���j4��ٝ�H�������m��������'B��2�0,��W�� �}d0r��:���%73����E�[:����ߤ'���W�3��Ny��KH2��!��8�!�M�}>�c�ލy�h8��;���ei�$�o�yˉS;��cӄ�hb��_Պ�5+���;�h,��s�Z��:"�k��[.����Τl�עHx�f��"�:��7��h�# ���S@��2Z5N�=�u�7�C� �� "8^�D%~�����+K�G�A�O�a�n>{%��]&g��Ѵd蒴�ا�b������-�kU�T�I�uX�&�F��ZҼ��H\B�C��)0Dk���5Ay��$2cV�]��͚��Jd�i�j	*e�@�H������JC?���nMXL�W��*�M3�*�,zjɉ�Qw��6��Iw�8�ˌ=/����
�4��:�v}Ci�_�ӵD3��Mz���z��@|�����瘬	���	<p��C�+2��p��+���Z���Bvg���2�^�d_�>��=��` �5\˞e�F�ۨ$)��ۉ���=M���Z�%;s�_.:����G=f?s(6\ׄ��ЪT"�I�ٌn �dKEVA�Q?����t��R��z��ä���M�|��<h���+M�r��^�Iz�(�ܼe�-����l1��\nw؅)2��P�n�Jo!�	��&]Bf.֍�u����QZ��C�vJ��j���W���Q�/�0R�4؛R{_@B�1�?Z��'���Kۋf���8��{y�@�:�'�c
|�<����xDr��b���j~iଘY"��B&ݔ}��"�m�[�_����=H���n��8�O��Ҿ�VZ�̰d?�S[�/h,�-�J�C�B�m��l�F�}�@��>�� v
���`,t샖n�ȯGdG�Btu���;1�	c�����#F���O�P��qӕ���Nڲ��Ȉ��[����8�V�@yߴ�\�7	mRS��R�=���b���yl��A�S�������S�a<́����E+@灎oߴ���,!�V\�q��L�ҿc���-f�6M��9S��6�Ca�����N��Y,/�R#w2�O�c|�r��%9#��U&ޯJغ^�96�j�fp����1�D�6� LM�a���i�b�ia83'��U�}V�ՠ�Y�Ί�.��0&�n��^ˎ��C]�!�%m�/��J<)�l&�X�r���m��D�~o���p�T���U>�>Q ��4p���ܚg��v���J�	c���_]�i�f��]�19�# *砠��LZ*�����������Lf&\���x�ǉ�R�����BȑHaOn*g�5��L�Wg��<��3���$`&���"3zW��[�y���x���z^��xQcL�k�(��S��H�Q�M]��r�s!��z�^%������u�G
S(i�4 I%OZ�N�N�?Pګ�ڈ��9^��eF`��	l./k<���}s������<>'�T��[(�^�����Kx�.u	v\6KZ	��S8/m�~���@*F۴SGʱ�g�س�%���H7��1ej�0������Osji�[���g��ˀ7��$W��f7������s���s�Z��^�Z�Z�1���Nb�U�ﳪ;��\ԥ5Lzy��L���Π�7`�q	f`|������GC��0D2٣��M��{dPs�Wgہ��q�K��MDT�3¸%'SH�'�p!�@�؁s�n��J`y��_vк��=�zf ��{��$�)�C�p���7����f6���$�'>�_�X�M����m�
��.1����0��j�`!�G�GqSm;f����Fb>���x����>��1ϙ_{hG��jT���@��P&a�Dn�����X��cKTSc?7��u	�՞��(ڟK�"Q�_+��Z���S�E���Q頉�6�-����~�E���Ϸ4)�[�6�
MK'"�:�Kos�<XB�oA+�G#7󡑎�@�)�7>�z@��^'���R����r�ʵ�Gx��$�����I{��t�[jB��@\`��_��D�'ݞ�1A��6���eA5�΍�>q�u�̖�-N��
�Sg%�.��[�
��/�d�� ���my�gfr�9�>� ߥɎ���A� ���4]#�Lo݊���3��MU
w0��I�Q��S��1�Z�G}9���]Z�m"R"��d���D��j_s[��M55��;a8�HN>���t�KcCӮJ�~�������{[]wS�T5+~�Q�ì�~i��D2�F�`�VG��ɮǢ�H]hLK�Y��/��ɜ%xo����0��O��yrm����P������	�'��Q�#��auʐb���':>�Бz~]��T��K����qAy�~������<��R
Ӏ)̅8��l,囵�?�H�6���ɮ�,3;,�Z�)���Spe���e��=wW�_�4+J`���G?������f["�jbP5�ih�^�.�6����ؚ��6aj���~a_n��+o��᣼r���t� ̀qs�<�ud.�X���a��~�I��%٪R~��{x��;��4Fx7�}��ӑI��ҳ���:���t��w�^t���2p�NzKr4�U�:ߜ.�{��F���y�p�������+�Ѻ���39���E�i�[7VC{/h�����^#��'v@7�b_��?f*������{㻯4�j)1�W����HG�LEh��N��[�W���ҝp��<�|�^��K��{N�M%kh�HA
j�~<��E��IkM�HN�-����OA��y+}GT��u���b��I"�Ƌ���N[��#�o�i�2�N�1
7Jh�Ђ��堳ԧE �.�	G}U�� _���b��7���Q%|NbX�M�j�(p�bo'g(׹�*�B\c����1��9Wy�VO9;�U��SV>��mû�Lh�H\��� ��]F E��k������8@)����4��υp�/>1ʬ�υ����2�����r�8$���������ehL�d�>�BĤ���Ȱn�/Ck;��+`�:�L�"���f���q<O�5턷�8�,US�O���P�l/MCߝ�?�o��q���b�5Ja��Ȕ���ix�L�x_S�l�zT�QH�:��纬l�B�k�
k��7@s,�siV�!�r�/W�܄�/KX��u���k�;˶�r���,��3 �<r�?�?y4���V�����@���w�;��w��d6���۷�C���ۼsG+���(3g��s)p�M��d/���z�
�U ��G2��ķ_�L��JA˞.���+oOu�ק�"S��dѦ���]�AB;�/�dJK.�}e��/`x�e���箛Z9\J�D#-5x]uݪ��ݍ�����Ah26[
���-�}C��Z�����Z`z���1[�ma�s%�f�ʫ����vf ��<�̾���-_�e�a�� 6F5+5o���z��z���h[O~�:��p����<�D!��XY��b-�،� ����X0X#�;�&�>[�j$/(bL�"�F�h���ݿ:��}V�8���H@��֌sƯ)mj�9�}�6h�GkV���[�Z/Q��g>Տb��r�V�Ed�O�6Eb���Vp��F�
���8�$Kqt��
�#���pa�m��`�O�#
"�i�����;��f��lY��������[�]Wj����}ZA�O5��W���9sA����� �r]:5�"���*6�f�#>�1�`�xG]�/�wϲ���$�}����ɕʇNMP���^�8
&S�zZn<q���v� �	�}F���tĴ����s���S������6]s�ag�.�H#��<�%�j�'��[Iz+�Ar�^�5��
3b�g�"|��(T�du��3	,�hGw($H|���5�T���k�-[�>f�9��8�2{�2{����Ր���oh��o�#��@u��)��;����&�[1�.,0"��̱e�c[v<́�k�����UYfWS4ɘ^:N����b��_k�_�[\Gu�&��iI~e%�w��8�[,��|����t�`��(s��^֕�ΧD��0���aq9ƅF!�e�ߝ4wR�i�^����x��j���]�ܘA�#o�޴c4�Έ�i��;��:�Q�� 6�'���'�7�=]\yj�ZJ�_��]y��gU��K�O��F"Hbp�TT��'ٖ2�<��&X��T����RV\o��ʤ%LU�XF%j�N���.\m<��UNW��҈�S���$���j����!@o�j:3����H"i	|R�4#��?:�MD�'.����&p��T+;M5yIDI�x�����#"�U%}>��$?}	���m&�ƒ�f�w�S��=��!Y�a�����>��'.\jm�L�"Ʀ��s�q��f�j���	�١�8Է���J31�윇Cdf��*6��=�1��S�G��E�+"��J��ط�u/Ȱ�)�����8�����|"Tۤ�ٗ�s�-/b�H}y������R��s�A��Wd�'�$m����`~�p��B<.������Nf����9�B�& ����"�0���0��}�n������x�x9�Z���D�f^}�ni�#�NN.v=u@; E�1��-M-�*�f�H:�N0�*_#4���#?̂.Ư����;y�Pf<�����~�>�!���λ��j�h�ݡ�ȑh$�˸���1�������'K6���Z=&G��{����%��A�� �z�t�a�f�OT��c�碘�S��R�j��n��ewt~�S��-�%@a�#2mC����T�,�ln�S��To���f�V10�{@�(}��8�b)�0C�K�`?�l�8�i��	j�+�W�����݆/���.�U�g�90O���m��C���A6���%G\�-;���V��ҹ
�лS�!�y'�=�f-�:���=> ����΋żc~��T�q�t����A�8r	b����|m t�*�6/��P�Ǌ)� ٩�0����Kf���'I�p+9 cI�97s"5Z;o�Tx:IT�;y�{�{%�y�������،����_��!6��Y���;���B~�E��d���j�� ��
��� 	��{SS#�ݹ2��"���y��A�ЎиG'j�'9�X�v)j
�K�P�hOa$����j�l˥D�؏Q�+�# �U.^lNpe�+�N�{ �����B��FKjW�� ;�o���rƍkiR/������os��-zA8V�)��fm5��ZC2�ߍ��E�m�uE�n��~o��=N319���ų�n��}SjO62}"z�=�+��>�U�M��<'�����;Z#���yx`�$�fv�8�j��0{MӒ7E@ ��Ϡ���je�1��Ưm��Zne�6�1��2�B��P��)�
��H}��H�������l�2�2�)�5��ClU�n��/��c��o�N'd�\I�J�YLP&GWK6!�ߙ�g��6@R^u�8�&�C�
Ӣ��E��9� �T�����9�F�{SS�r���w���hQg��hyx ��F�1��1��`��c�T�j��ʾ�#L|YQԿrUw������yz��(γձ�-p�Ll��|�(\�j'���	i�1�V@�&���`��nƜN4��,�qaL\�.eV�V��[�&�ɫ�I�v�"��$��n���2̛��+7UK��"�'��K�0A�LR|��A��(1.ɻ"����jV_�	�'���,B����i�ʅ��n���>�yt��e��b{�8�H �K1�n�����-���]���啜��<|����W��" �r�o�@��3H z|�ƭ�R���~���@�Al�ŽB^M�dü���"s��?����P-"�KJ�w���pt�n.����?�$����v�&ۜ:�;������&�։-V�(Zf�C}�M>�7%�SLWrx�G�߿A[��s�5J��i�.u
��_G��EQj�K��73�aQ����rS��|Ȝ)%;��t�T#����}fG�~�7��%_�^5ަ�I	N��v�w�مň4;ߣJ��]JH�1�x@���껩em㧎�-�s���}��]�_M�z��9J�ʠ�p"��;��@щe"J��z��KA�����>I-����6��V
��4���P�T���Y���@Ϩg6Od�#ȏ�<�Y_j/��Ĺ�uf��Q��$1�X��, ���ߝ�¨�D�ej.1Z%�@��W+�윹�^�P��Ȃ�������9Vc���Se�no:1p�-�c�U1�Z�W�0�Ex��+�t�� �l^i�y) wMO���������F �yA��������)<B�O)��z8f�=Ew��Tg��R��V
G���*K���9���O���Ȓ��e�tQ�p����<I�}���0d���[?Z+
�Qd6
��YrF�M�Ia͞a��O�̨�8dkB��5��'jV�L�$pZ'jv�	��y��m*|�2��=i�v:}v��-u���wS<�)�i+]��A�����]���ݨ��@�i���-�_��b�ԫ	����x�/RנA*��y"&�ڽ>p���$��Q��'�t�s���� �h6�?H�̱��Oi��R��zw-9Y��2�������q��_?�IMo��}
g_J!&�����fC`G``�5��JQ3�l7gݿ4�rC��P�CT�\�|$���jC��:,�O/��3��l)����`�j��9���8nw�WT���us8��N.���D�Q��ϣk
O���D�"�3�]�"@V�YS���1}/�e����nN���p#��h��Y�k�_�z6}&���Jn[�~�T|(��O�N��|��Z�r�M��PE�a�MB �w�Xo���Q��	���Ҁ8�ik�� �o�#F�p���������3�@�੷^`��ǘ�{7�v�9x}������ ��m�Id�U� q�܀K'��d�9���;.�oC��fpu���kjW�M0�&����T��ٍI}h�X2(��5p�d�ݠ�kj�d��	�3��H\���M����߈�I0f��Y��F��^����ȰR(vю��O/~�ro�F�u��8�j�x�`�O�@��]��n����u�7"�Wt����b�c>f]�)��2vg8k�-� �;��!��Ԕ�n&E�)��w�>�z��L��i"�q�%O_Y_ԑN��k��U�24.$h�A^�7��ȪW�r�����"cq�X���zdw8�#�XՈ�i��h�;5u�����z�����,3�*�4��XǼ��5̪z��(i]Q�<��.%(��p��L<�	������xe���-+5�U�ehr�������9O=�;*���9�=�t���A��	��&�D }����:��i�����h�����UO�-8e��U/T���j]lF��ȅW>��v9�!RJT{���~������Ŋ������U��P<�c�96��i�d0�1,���M��d��ȼ,D�~ɣ��+g���H>>�+f�->��$������f˄��I^d�Uo�����c�1�o[�p���:.��x��F�&0nXND�~|��j���D=$&��:��}����둋�Bi��'CXw<y�(rc|��*ƛ���� D��,�a�0"�:z��c�os(��B�~�{��J%�ؾ���8l {�6mf]Ē�i�]��s�;J �V�p�����)@&� �����t���=4�!k36�ҝL�e��k4��0��%�-�Y�6�( �p5��YĚ�z��7~�3�O�(�����M����n�?$CP^c����wVI�Z��+to@�Z�$�#��i@##m}�R�n��M���/H�C)E��t{zg�q(=�{5���2�D��A���[�����0=��a�'t�;K�Ǟ-�Z��F�%c�Z)&f��z��ȗ�l�2nߕ�q��Lh'�u���
��{+On�O���h������9�Y���#����9��X�=��պ�������͠��u��+�|��^��_G�P�0�'̓�'P�*V���ݼF��ڙ;F�&�R$����@��K<�._�Hmգo`Feddm8OP�k&%/>�>E��A��{!�I�E����|�Gt(�Є�)��g��G��k��fmTƧ�f7��4��g�v�rB�� G��A�k	n��w"1�2���S[�U�����Uv:]�j����x����r�8��'�9ؼ�*Hq�&@D�5꾎ʅ��Z�,�
��ԣG����O\@�gg7ξ���)Y��8:�/@���KB,IxTi��~��.�ë�en*�4oO�����;Q5���u~p��i0�Q���C;G�C�EZ `C���LG�>
�Ӄ�amH�pYg���W�&piR��F'�������m�뿟�B�J�Ђؘ�P͝O�ny���<4��,�8ұBx�7[;z��A���ؽ̓R��o)����@�u!"U�������P�P��"k�$l�[���M��҂���BA�?���:Rv��v�:q�ɶ�S�֮����[�{Ү�Y��(ԈC���*_
�r���m�zb�|~�A^U#3ar�R[�����O�]��eH{���E�\ɼ�]��;�cx�wJS�y�ݬ��v�G��F����*'ԙ�U)�WU�x����������2��ڲ�]�B	b���׈����]�)�g�)�"55g��k�7w�i��=���R�Zl�c��r�@8���0<|�/O���p�t 3������f^�
l��ba�����էfy�H�r�sjH�}���Q��E��$+Ϛ�}r�-�ܮ?��� ��g}!��e���؇8�%�_wGJ���K�1�nZr�@����1Q�3�>C���Ns�R 'A��ڃ
DЕ���@	5� �нq��N]җ�}�,��f�=t�N��䡇�#��W��#�>{�8!�E|,��T�!�o"��e�0.B�ҭ��;+��Ysj��6�r����O�	������r�V��5�߮T�r�A�[u�Tp$X~7X�!_m�jK�r����T-��:D�Dѫ#�`����w�QٛU\[��܃MS	���׷���BrݰM��� �Y����"��� �z����8����o$w�l��-�9+Iƽbh����L�Mu_a��Έ�k��N]s��6e9r3�::<����N�oz�B�W���_���P@���]v�K�t�E��o[��Q1q�ɾ����Ё)������G<4�#Q� /Еk�F�Q�X_`��YÄozW1��{�0��b������q�}p�s�"x9�@ү�ke��x4���"R�BQ�N�t��YiYQ�Yu�5{{�]f�m�6�ᙷ�Z��\(���7q+	+.b�,�q�=~.Y;1Cpc츉<½i�9������pU=�������T�R2��"6FX}GR`�R�m����d���ĝt��̼-�
���̝�&�9���>$�9����U�whx]t:�0t���.�,��h�UЍw�w ��4�w�������������������E��5*���My��Ào�d���-8pE�
$�x�U�F�T�t��Ҡ~�}jF���[��3�1��>�\��v��Rȁ�vk�P8P�d�p^� 
hF��%o��K�� �#M#���<��C�d��"����ܓd!�O�A�)������Ge�̯�����o��֐�r$(_�����^���p�#�G�-g�ޛ=6J��M'p�(��#gxe�^�T5�S?&��;>=��)XE0¢�Y�Q��DZ��~G7Fܼ��T���ˇ�,Y�i���������s:���&e����*�����/�
������XJqW@�Έe�M8����Q�I�nsL� �$�,O���L�&%>����Ȉ��e�K���G7�%�R�C��^�n|5���~_קuj�?7Յ���b{�Ϗ�տ��e����ΤҢ@��*�GQń��2��Ȁ	!7�==Q�X+!j��|;�W�˼�/βT������?�Ds
��w|�y�d�7�B��f�3���&zg�jb�B�����V#r� �Ao��c��G��Y�-z#&ç��}�g��VYY�ls���.�G���Q�䰽R܃I���-�#�).�e���Djt!���Pi�J$��Q�r��C���\�(>һ)84�w�@a��V]�)ě�45#enh��wK�ոQ���|A��8�]�._����;X�QZ{r�W�dZ�5p
�I�ٍN{���mR������E����3O�ȕrX0w���*?ܒE�K������weӗyvQ��{�g��F���nx	>K�胉-x���d:�-��:˾S�F�#�G9�d��'�u�nĈ�KJ�jsZ ۷a?{���N��6*q�TipN�yC�-XЉ�{�i���1��Qp>�}nyMG�@(�
8�Mg�Uh�۲�A&�fs����}��әX�ӯ��r�ӊ��V��lN��>h���Bh�k�\]Ic�^²�����_3f~^6����]=rR :|�l�+@;�tМlx�+�o�|�f�x;8������\�g�!&��ux�h������VQ�X>��+�P�*��A�����Q�NP�s<�k��M\��
�,�g��ץ��h�^)]��B?��J�V�t7Rz�aP�Ys�C}��V�X��d���>�{b;[F�o��{���RL�g�G]P�g׋�KV,#�ئ��k �Pj�s��ɰLit�P�v]=��W�,��F�����\��3
�*��NR��8u�D$����G���Fc*'^��^�ؘ�A��(E�|��[��(�R���7!��Z��H	��=���ㅤ�&.�oh�Ó��lH9��Jv�VM���Rٍ���K��ϰ�Ms�G̓+~��h��W�Ϩ��YT�/��s�x�G�����5�@��TP�q������B��)��k�%GQ�Bp
#��W����s�B�
��~X��ҍ��x�!,�3R65�hqS��q&jSyN���?_�,���`/F��
��ݕ�|30^}2��dZQ�"V����~�0mw��kt�S�&�����'��ݣ�c����$�^���H"0�ڣ=�6۵����HE'����#�W�e�xs�QE&�g�H>k�ok���f��|�w�M"7�b�)s��i8��i�"q�b>(�q�-Q��g��*�����Ɯ�`T㎕է!�D��!:�a3gOD��5����J�õÓ�c}����i�l X���sɢȰ��#T����O9`(���"5;@�)8s��#��	��`��(%!VNU��I�aT�5Ї`�C�5c��zy�{�K<m��R>SrxQ\Ɣ�S�(�pW�{�/���K/�_w&T�:��A�htEV�hӯ�"�Y"�9���xt�u���4�#�S2W��#l�t�t@,�4~�"���2J�h�s��<݈sP��bOaԧ��#�C��5��I|����{=���)Y��/ȣh��o%܄�5&Ѐ�0@5T]�/��p(�Y����k薓x�Ytj�cj�Co'�m�*@�W�'Jpd,���-�LIR�'��|U�>�d��7P�y)#�f�5|sxi����)���� A�������AZ�T+��҄���{Ђ9��j�Ԯ��v�>��I� ��L�ⴅ��d��[�װ����*�5ͧ>*�%���T��h�iJD$��/�����8�%��G�K��䢊Ρ!LE���ϟ*KH��D	o��Y�)�ݙi4��%7��2fq(Y����1��_����١��C�SSŸL�=)�?"�Jq�0�2�P�{��܇hǾ��x��Q���LNC�/��o�
H���Jׁ>�sw�n�r��� �,�I�Y��y]rc8�=�~o��Q���L�7��i\��J��'cW�ȋ��~r�g�e�k�fP�+Ec�J����Ő��I#n�e_�ԥ8�h�A,��ݪax�Ƕ�n�P*1��.Fn;g1��Cm��7v�[A^Ze3��o��Ǝ��!����6@��6s��}�#��)=cC
�I@e_�����w";#�����5Jȷ��}ͧ13�iL�@e����`��S���lv�B-o�/<�9>���!|5x�m�G�p�������� ����1m�+q�K�.�X�,@4h����� ��3��l�XC�9'����v!w�����R0��=���42���p��$������RD@��)<y��:��E[�y*Ѫ�������j���������/9�9
`E���)����E�	�=�k����f��yc)}\)�#��r��Y�+��]�� ���_".sD����8���"�ݮ��8��X���(W�	u2��s\5i_.�NI�D�^Ų�=�\���K����ٔ8_�R��)�������La%%t6��"PF���O��E�
�k�\���b���ދd��>d�f�>�QI;\]�K"�&���.[M����'�J�!�L7������hГ3Gc����,�s��P��_��za(��Pg�3��!��a����<B;���4C�LyzU�:"���J��W!v%�0�SdwQ^ASZ'*lK���mh�n��]-Y���V*���N	�b��:{	�_�7�њs7�n9��vY;��4��G#���9_j�*^&��7Yx�fB�r��d�3��+2m5
�����{	�"���~:�F�ψ���MNЪ�L�����
>-}:F��I��?%S�H����f�HF6�hR�ZB�k�`�L�=�k d�_�At��c �a�z�����m�
(ϵp�;L� �UZ^�:��ƍ6|cj$�L�������H�`I��H�4��9i��O?UI4 N7�7�xD2�8�����pL��2��6�u�W>ɷM���`�h��^<��,a�Z��F��V��%�NF��q}�M��C�X!�y[/D�@�	XA�W�	�𢡄=@CbǊ᫆�� %���o�?Ιd�Q	$��7�v�G9����xrl�iNz߯��C�,Iu�s!WF~9�ɺ�i+��
w%�j�I��5<.�@���]E?F9�"1�C,��U1�w3��50z������/�\3�z8��rGE��Hj2�nrƦ @���Z��Ch�[��nú#o9���Bf{r����\u�@ �##��:i(��(��Jd�v_(M+�yRFm���J������~�����G8�;���N��5�!-���)���ՙ��,	I/����[��K��=�S�[52��Z��PZ���gڪҼWJJ$U�@�F�Ea5T#�B]0^NgFG�c���\�2u�&b[��%7���W7M͇i�T�����pc<�_�hrtQL�o�M�4ݣ�~1
�c�F�?!��S<�����X�!�XU{"⵨�I#���D�>�f.x����`3ta{���
Z��ӳ�t��0!���< Ѿ4j�Z^��p�lw{���b$�����yX���ަC"_#��eB|��T�-�����.Vi0�<?�U���hy���kV�]i�B��j++{�"���M��\5k���|�`���RYRc�����tE�jR�/c ��VI�'�^�Y����@dURH*�Q��.�MP2�c�ꎓ�CP;��W^q�@���/��j�������`�`ʿ�Ù�Z���#|���gzetE�s�}	�px.����Kah+���϶P0�{K�� `�j��YSz��*w��yO7�,��B V���FȥR7^W���Y?>��b����Ѝs.VM����'b�=�z��k��P���s5���n�T_!��鶧��=Cvh��j�>���\i��'C����AZ,��8�iL���������{�n����Ŏ{P^�λ�{�-@2������S}X��z�U.�:�_a��_�3ԍuÜ�[}�����v���IǶ��a��eig�jD�$L3Si�qe�*�T�Җ�p,M�6*oئB�l�rM�2}*m:��rI�	���IF�1���/l�&�O��cQ8P�ѕ2F��F[� 靎h*QFf@ԗ�)Y_�Z��/$_�j�\kI��!kI���+�q��E�A�����Dև��H���*2��H}����:�:<����b�
�o��ʃ��z $Ԋ�LoIJ�%`l��M�hc5�6ZS`��P�!{�l��L�y�]�	��h����./�L ����;�UZ+"�Vx^W�i$���P�ף{��I���}ƭh�f{]�j��M6�Y2�[6��)�1��붼/(팢}�\���oz$\��Ǔ�~w��]i��$6?��󝍧$4�G�v�`Q�tOq*74qm���C