��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<�w��Bk��S��9�h��7+|��Q*����)�n��t$��7/qf��dߏ��/H�`/�p։�x���DZ+�+���
�$�s��� ���:�H�RI�yn L��s����4CCw�	���B����)Y�
���((���bV��"�k8���aȳ�t��l��G��[NaS{<����נo�?����~� �!����=�}v�g���������{�=X*�.���c�_M��k}C�e���)�U��o���l��	3�Ɇ�J��:|��+��q�йt�1���0a�-�e��H]�~p��1~3��8)^���-�y�˭��C�G3�45�cL4c6�txbA��F�ږZ) )�U��y��k�������Z^,�!\v��T�彧k�,E]RK�<7�#��C"�r9�p��n�<Ī+|��ǋI�b	 �Ȗ}xFo0[�Z�
4j��kl�r��dy���@��DGD�Xe�%<��f\e�u�IqN���!x�l#E��L$_.����d}��)j��ge ���:N�~�t��9J�_e
����i	H����q�"*0�nID�*u�c���Ѝ�;�n����MH�A �!��(g��|j��gL��J���j�.�e-�)�M.!�̀ؐݟ�|-��-6�ݷ��o�"�ϴ���3f��݊�\���7j���?���P�iz���;}v���Gp��MHO(�GAsgpy|I�1"2���Q^Bea�-my�NK��)�:O{���:T{�H
����LE�ݜ?תד�$k�����[»��D����!�3�nC�cdP��� $L˹�a���pz���n��$}��OOS;Har�H�ҪUdr�Ө�<	��V{bS�K;뮝q(Rt�dx���%��_lY��.��]I��n�o��[��g�A����n�^�ZI8��8��
BYŀ����1�����+c���'�����T��+Rێ;B��P�`e����5�Za�����H�����Rz��e<i�6����+�ÔF�����Y�t���A7]M��};��.�\�x���4x��u�Hrf(3�ΰ]���(�/o�RFG��T�a#��Z>j�;Q\FS���6g��-����Ys �k��zF,2a���"��`"!�����R ��u�m^,�5xPHބõ��]�?�tA&��M��'p���1�,��tupiɦ5����s��A�1rG�PY`�$	�0
#Q"&�Q�dotC(�C���t�%ip��ˠ��Z���ε�z_
��G�f���G�"ۇӷ≮86�	�Mx��e�}n�^�ű�B�Ǩ�5�-=+��-[�hV�vO��2��
\�6Q`�5wa$�e�^#*���A�E�Ŷi�Z���v��@�-��9���/<Mc>��љ���$���IF$&�6+\�,^%4x9���=.N�$�Gwr��	j�Q��c3��7�#�p�2K�H����u�I�ĲPڕ-��.��}d�=�k��F_��?�7 �cT���o�)В��y��� C;���s2?��
\��7��k�����:-M�1��� zfi���!�H�U&^��e=)v<N�^��	��H��=��-y��d����H��xW���,�d�M3�\6S�5S� 3����P0Ŧ~\X� 58���ϭ��_�EV��k3T�P��.�2ܟ��MPN�W��Y���>��G�1� :{Oy2�(�_c�qk�Y�	�YVY�EE�T$O OR#
+���I�F��i��Pi>L��5��U�%����
�V�'�L�ך�g/��3o���!���a�����97,��i�A�
����Yw[�b��V�E
�~d��v�N��������h�|�⥫s�)�ܾ�-<	�?M{h��|�ef)|p������T6�!Mq`�<�1����B������n�C�׏B0�#eR�>�*�$�
��� �8N�ٖ��Fq�&@Jd��9
� �W$%�L ���7D���P��H�Ǯ|����q�PbӶ�s����"�!��]�����:��x�}�V�����{�-I�~�zZ��fG)�s��}Q`��hxh슚��&�����{�+�}�K/6z�H��И��?5 K��zv�b^��(V�F�e��S�316r���]�[��
���+�m�(�	�������Lz��g�,\��R����2\�ٸZ1��3�V��G��*]�>i��i�PE��M�?�\�<����v\<�)-���O�WS��D�B����*cwWSG>�'z��m,{;׳�Q޻��%̷�ͲKX�"`��]�5�VK���s:���).%ՈW.���aS8yvyX�F�;�y�z��5'tm������<��lXz/h�������ecv��/x=`�(����I��B�Tj�Fp��Ӝ����]t�Ea2���c�C��3v��y�m�{ ۔�=�}2�,ʩr��#8����&9��>�V�NNg����D�yŀ0%!�l�!�t75��;�1z��3uff_o-��ꆒU�V�5��f�ea�Q�/���v	������\n�8?\���Dv���*�Q|��e0t�I��`�t�L���
T��h5�l���TC�5�}�IxHN���4��BU��@s6�:\Q'PE�d�A1 �TK��x.֐Z�ܫW�r�2}�2&��;P��v�aAA��X�r����t)����9�b�����(���7�hmK�����qg������ܑ�AKT���kOq�Hԗ�W�C�0a����k�ݱI��\��HBٞ�#̗4�g�?���}|�H������
��1��N�kָ������(֌G��8ͻ��W�'k�.SB�Zocp��RX�p	W���Hu?���"G���1A|kS�'uin����4�j���SX"�LuL8���a�z��pUa�����.�J�}}�y܂K�զ���IC��>5\�7�VK���9	X���o!2��Q�a��e���u/���ϴP�7�v�#̴֪_?�>a�lt�K����>���]�ȉQ�9t��TOT�}n�(�=o1��.����ByN�UqDL����
7��y�D�!��H�KG�Y�����}���W#ſ	���&�����λ�r�6G~:3 ��ʗ.�(�%��l�Q����&x�QޒQ�,�%�����1��<'7��Yo;��z�6N���?$i�N�[�%�a�$���\{����I�p�0�dΰ���a5t��P�џ�M��
i�k��U߮C�j�/��&�?�.��gu��H���["P��cLs����kЃ��C�I�D��Dz�f�BZf ��yb1�^��q�	8�Q��SC#/Bs��D��I6�z;�,bX=�t�jW,�;	�lc�|��F�F���\.x&��d�5�
S~i�xy)yہW�j&,�].�ŉwY ��𫞨 ��Ӷ�Vq�Z%�����ϑ�b��o���G[-��D!��"]�Q+C��"zxzz.0�R$_�i�s$؍`g� �j�S�d�@705�7����uy��B��� L�_�L����n�h�H��&;fB��Y^�vu��g!�_�y/�C������zq�V�:Q���QɜeqFn�3-��o!M�@�_�a(�@ҽ�Y��Z8�t��V�đ2�Ժ�l��J��Ui�����`�:�㫒�w\�z�� �Ԓ�uA����J��q��Gi v�W�Z!�"ܡ=~r�tj�#�_��Y$O22�/���v;'3�FYPe�Dm$�*���Dؑ�/�9�fu�s�(l�o2,5Խ����!�ÖG��&��@ ��4���t��@�u�& ˫41���q�j��#�~>�+��z�:�}�!���]�����`���O>(���x�ퟕ.����>&ֹ�kw-aʪ�m�oݿ�v/#�Q�����������'G�����6��y����gJ���U+��h$FqӅFȴ�����qƥ(����������}��y	�^(Hl�d�g�9��@��b׶���$e$kx*@�"o2��	U�j�C���fT��;X�Ş�ϙ2x�|�D�O�jvu���0�\�M�@�(M;OdR����v�#f[d��]#l �+e�ڍv�a9:@�4KrHkفN"�����rY��컸۬��w��u���::�qt���1��
|�t� ћ`�A���Ŋ�I��Iy^�@���\�b|]�8��g�_|X�oh�_���VU��J�.L�+���6Fؘ/�����9�#�%� ��ڳ4}�<�J��X�B32pJ�[�`�3��cO���VY� w�r�LL���>���]ûA�j�X���_1���\��w��b^�K��s�Ě�n8�*�n�E�<2���C�~�u\f�k�i��uh�KW��Pwb�M�V�V��J�Zܵ����p�����Y.�J�xl�L	8IY��B�@ ��C�q��g[Y���K��G�W��s�Y��G��a��.t��nX��#�I�D���wBM�J�f��'S��������v����Ơ��Ph:��g��n�h�2���j6��鱥2�Q'����@����O[瘟	ٷG��#R�ZwQ�e�Ui�҆R��M�d��=]���l34R�a����
�)�����N��ḙf��E�k�OE�F�ig6<ş|x���j��� ��Μ�Ӎb��n����G�2U����9/��8��+���� 5����.�L G�P� �c�0��n��"E��)�\=~�H)Z�%�R��+%�2�I���Yv?���<X>Q��z��L��l]��Q�� ή'?��K��Q��7�Q.lJ���o�@oZ���z��Q61�N������r�Ά/\���q����ӬV�D�O������Þ�jW�X�ٙ�F�%��;���<��%�m���ݯ�&���������@�<@Hk������5���@���Gh�����}����]��gI\���dY�O��q�@ �]���*Ng� G�