��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��I�ɖ�P�	��[�&�T�u�L �����wR�K����Ҽ��<�X�L.���[��"uq�`fm��\���t�u��Пwn��(�7R���o�M�q?���������p�6��s'��%!��ğd��B�yN��}��C���ߩw���3�����5��Ɇ�T��]��{D/:��r~�w�Rl�L�W�S'�]hNs�"g����y�y�7e2\4�4a	\��v/k�IG�d	_�p3չ��U�?������qL�n�h�%�����Ćˬ�ὢSM3�X�A�6-�ρ����<� ̕kd5;��^�A}��p\��,J�G��B�x����Ӧ��k���{�'��\Yo0"ӄ ���Q���������	���4���u�5��<3��}\��xR]��v��3��-Լt�-�T���`���(��t#mЊ�;��_&�MǍ^�	�dä��8���?�����D�8	TKp7��N���%,�=���@-��)�������W�G�&1�H_�I �P+���&��Em.O	�ƺ���m�w�u�<1�N����*򼑟p˗ ɀv/D,�4stc:�Ҷ�^bv�usٮ2�,c�AI\�(�Y�|;���U�DCFT�Ȃo��;�˶ݑ�n\
nF�o��=R[��a��]_?h�%�=�	��(��R��\� �j}r����6�2�R�7iH26z��&VF��f0T4wL&3;�������(Kd�����.����Bx]��K��z�r·ɏ����26����8��\��'ݵ��6'������䆃��s���}�ǆŢ-����
��V�UN�!+=�3�~H3���z�o�&ɭGR��YUV���^do��k<���Z ���؝�h�$���T��[KT�C�P�r��|}�����LY[W���J��{y�x�;(g&ϥ@[M׊�����8 ��3�mm���{{�V���I�;�}Fm�����9��Z�ļ�Y���$�/��F"ƺ%egw7J#�ww���Bu����u��
J�`$q�9 h�0Ɛ�)i��������M�M�~���^B���'�I��Y��K��|���ѽ�0��d�d��p��JZ܁�7���}�M�7�"^���wpc�7�C�}u�����a<㸺�x^F�Z�L��;��q�I�ۋ:�'����Z���ELe������m�&I�-j�P����/*P1��m��ot��u��K�>Y!��G#�$|Y�LT�?Z;�P*'�S�q��N�i`�jA��m@fr�YꦮV�����`TN���;��0Kp�_�e�D���\%�ȅ�Ņ���$�<Zf�x7����U���Ngr���'���i�It���o�;�Q����N��-(�fd�
*�m���*�v释$�01�Sd^T����1%��+L�=��#@�z ���C^�V�rX�����Y2�kvTU�롥5���r&5$	g��kG�x�p�ي�o(�']�H�LΝ��&�?z�V�ʛC��(��v0������I�K>���Z�G�fc��ŀl��|}���5��+�R\�=�ʨA�������:�Q���/��r����Q �:��3�V�i]����	�I����p��^� ����0��%.��QY�xpg�u�Bh��Vp�<�n�����͙\�I��	��� �(���V_(���Դ��p��u��<��^݄z(?�16���¼b�'�Y< 0"�a<�/,G.�@�_*x�?��y�V��E
9�*k�p�H�W|	��Wf��kS�39��A!�����9��l��@;殛�c��;�0Ƈ1��x:q��Lr��Z������|9}w��=��zȽ1Ң��o�K�H��Z����L��NA�V��B��L���B�1�6a����U�QNp�sHǍ�ߨ��D� �� ��3c[}p���d��gM5����x�g���O�$=n��G#�Y54�#����e���_|c�k���<`� g455v��{	I������3�A��[�����Gy [�H��}�������=i�}!n˹
[�$­�J��01λ7ԙ�(�ު���z�(��	p�3���^+s_�Z�s"v��?RBZ�U���l�da��F5v��� �D�P�͠G��'c��@ Ǫz^pIumB~��o�������Oot>�$&�K�Q�N�� ��B�~�`i򾝣�d�t� �Z=B�ܠ:��dR�;�WبB��Qػ���#�o��� ���	��6��=<���yT����B�L��%ڲ�/�熪����n0n��o�'͹��j.c@�����S��E|%��̔#�Sg�i��<��o�AU��Ǌ����� ��Z?!��piP�7�(Q��dܝ�Y��c�/N��CnJ\7B�p���k�U�W Oq��ʽ�2��>��,��f�ڤngL�������7NJWh��d�.�Qp�<dN�,qa�m-��씊����t:�@\Z�?T�,2���`�$}�����N�Ɛv�+�#�;c�vmԊVfj���g�1\4x���AQ9"U��:v��kH����@L�6�|(K�f2:_m\�ֽ�2qN���4���a�I��pکW2��ђǬOT^2�$!C�G�w��-D����R��i��SW}4Û��8�cyS���N�Zd������oT@#͍N�Q�]c�qM��5V>�i�^��q�X2�����%1Z� 2�h���qp�TÊ7P����f ]sN�S�7�Z��f�f����6��W�R<��=�Yf�5-�0Z�x��,�<�z`�J>]T�%μm0���-��ü̐��)/�@Ɯ`�	w7��v�(j�4��I��:��m��V���e�?j�j�P�ǆ�m�c a��ּ�C�~ـ��6&Y�}�>�]mX�VB�BC�6�J�7K=�ݝ瀳��,����Ţ8<GL>�����|���@֮�'���l�A�v�� l�+�H;�� V���旍��Фs(k��3{F��~��rޥ�-/s:"��^x�����	��J!:�,��>�#%�A�D���м��3䖅K��Qn0���s�c�47�����[�p
i�`.�R@�#��J �����Etdųw,�]$@3؉��T�?P�f��i¦ñ�Qi��#Ɓ�i��_F�he'G�������J���3��ݑBSu���:��$P�3�JI)K���#�Pw���:�oT�� �`�����ms�Q2� b|�Fꭊ�w�Fe��[7�Ў'x֘�:ڰ����_蹵��G{�#ZA`]��A-��(��ءf��{��|;0�獥��J��ZJQTV�v�K#����>➫��R��
�j���xl�o��!��6pygS�8v߉b�Q��[$Ӳz� D}��;v�;���p��[@�wu W��3G�煾���=��tCr;��\) E���bY`5������2��J��������t�~�7_SI th�����mn�����q*욥��%e�.w�i������G��_��,�8��&������� 7߄o5ΰ�z��������[*#^����j|�L����W�0��#n�$��5\�p�(:c�W�Yb�2×���p?%���)���
� h���D"#?�������5h|�l05�;,@���Z�/"
���f�Y[Ʈ�3��g�|Mp��9M�����[ӓ�Ĉ>������!�@�{ϥ���v۹��с�|��JUfb{hxy����s�