��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|ḱ	I*�ox��͝"zܕ�=����T%>�����,<}��r&�:疃�)�1��N��oS�I,�	�P_� ��^����~\��>��[�n,�Uih-5�* P�3����i9t�wK���g0K
��%�ي��n����F<sA]z�'�;Fs�j��PuND�T���芞tE���`p�����cjV��Sd2�:��@�:�҈���2V{
��|~|ȸ��rz0�9�*��9��u��B���BB��'�-��2��)��@���G���Aq�&m7ׄb��0֛,O�hv��O��V�ϕ�`����r��(�M��4��k���=1|����5�m�CQl�y�a���d�!,�ZN�����Ph�±w��GOl�p��0���6u���f�� �q�F�:#�V�w���'��Ɍ�����G�a�؄�����T�V����8^����N��6�k�eӓ\\uN]�m�΁�����ւ
e��6F��q�fl�P|=��,]X+�w����?�s&�j���	T'�����~��E�m2���q��b�_ ZS�&p���Q>��hxܘQ���s��T�1P���Գt��햿�E���:���N|��1DE�#E|R���H���IT[)�H���"��O�l2�7�ny�L=~)�K��FT׍�3�H?e���ͱ��!>�?��B���P���ɉ�{.� U�D41}��
}���D��E��q�H����z=:��-z�>��H�f$��6J��+s_���7S~y�.$,�/�|~ ����W`�K
H��9?����g���U�閪��-5;l[�\/^�+�î����f�eh��z�qŇrd��s5�8�<�e��"Q2l���F��o���"��w[i���1. �=�]"���A�oMêX�B9���Ӂs��lDM~�hzu����_q����}2��,ӓ�*IBgF���/�V��cߥxq��ƐH�A�j\z�?q��3�)&����I�!���*���ס����@7,,����"VK�cd�tx��wq�*|���$,YI�W�����ܾD�mf������^�����|�@���:Ƥ\c���8S�3���gz�-��7�UB�^��YچQ��ssc��-2"r5��vh��G[o�C���������,�z��׏�w���j%g��%�;M��J����Kɠ���U����8DLM��7�h����Φ���U1x*���g��Pi�/��z�WK7�]~� ������F�F�)Hk x�e@�4_5��$����vvķ^Og�'�)�d�;z4����fJ?<7��N���iX]3枱�7:"_O5n�ٸ�k%-��C.���}s'�`��37~ܗ��?e�K+�O�Λ
8�a�$`��Cm��"�ĒT[�?�k�M��]��c�$9�0��_�-4x[A����f��J?�^���R/����
��մ"�Vс��t���3�>c��f/����-�*S��`c����8��������5=<�mK�Z+;¬��3I�<���|wR"����8����t�fm���3&!�"mA�k��Q�]��E��V_^�M��Jy�E���_�Ц�>����]O���9�D �R��Ԧ�﫹]s��C���z�;�A�tFy�^^8���U�J���������GN�l���ֺ�AZ�C~$し'$@�|zhZ56����c0�HNe �dF�K}��/x��Y�pۗ�<9.mD1�uJQ��E�N>��̲7~_._H�`��A�nu&�?�ͯ�x�(��,;��|h�,1�7�@]��bќg�{j���c_�/��%�2��z��ejԴ������Z�88X�'`���ש�W9�����x*�D�_�cT�ԗ�wMZg��9Ӣ���nZ�O�a�c�&�j#).����$�@�TءDs�-]��@���=E�{�1���4_�$�
!��S�=��pQq>
Y�bN����."-LE�f�5@�"��}\}H�A(�&�1'�_�_�:0[9��>'�Q�s9�ː�x�rNT�uG�R'7�Ƌ�L<�aM���]�@gzԝ)�Q�d2︓*p�o�?���� f�b��M�!��|U9&׃���:{��*���;�Y�8����+&K!X�eFO�WI���g���X����כ��6�t�����J�;����E�6h���G�+96.9۬�c�΋��=����������s�. ��w�����QT�+K���W�n�L(�G���9���g���#y�Y��Vzz;�������1f�ī&�����QfI:z��hʙ_����Ao��F� �Z���O��:��)3p���MqeC��cs[��Kc{ƒ�K
���:���@]Pf�RxH��^`��=e�)�c)
U�4�4��v2�Pݘ����N���C��~TE�a����W������Т��僱�����{��T�u��A���J��!K2�S�������¶yP�6^��	�d�����TH�=�a���DcM|3�����E��f�L�
�����D�����Ne��B<*lr�K9�����~h*�.���6w���X��2�ɶ�w��@�t�QCb��մ���k��|�y�H�`uϝ�okA�&}!`p������3��Oi�K��Xڎݗ��ȌO�@m}����rۉnҤh��T�x?tt���"�y��.�K�A�fF��"X=e�[�|������ L��Q�GJK�@I��t�Q c�"6H�x}{�iӁĮn�}8�!@#�F�[k��Rl�l#��Q���B��#�!eh#��T�G�����.Y���w+H@���c��cӆ��&���LS�X4�Z�G�3�������2m��!�r���R�,��{� K�$���xc�A�'g�����F��s��¾F���-<)��R�[���َO�q٠%5�iPˌۮS�dN;L�F�l+�aԩ7t	+^��
G�^�$c�����cn Ɏ�,t��Q������+����\��<BK;czI���f$�G"��Y�k����@n��CH�~O�	��/�
�C%bB���`r[���# �G(5�?�� ���cl�9��KMϸ��]�sV�c�^Z�#�^UcIpj�`h]x�U�vT��4��_Pb^��]%R��(��vO�T�ai�^�*+�09!:$��$�<�T�<G�5g{H@fRA��y��ʠ�<��WR��n�k�=�<�ׅ�NDD^XY��t�C�E�8�	-�)%s�rр��(��c��l��7J�%j<t��r'9n5�4�yn~)�"O�9�NK#�)����]�u#j�Po��mlw���*N@�rv'����ttH%����Q�IŕfP�8��/�n��o��� ��_��Z��,����۷���Z;��ɷ&W��k��{�����B�{��G::���B$7�Ke�i�[w/�jeIf��ƫ���+љg�Q/���TTԊS��� ��/�E�����ڢ�O�X�5��k[�C�w�'�=����ek(���x�/E�ڢ
�EǕ�� �T�<��Г?�x%2ǹ�=D=u睬ދ�lg���̴ċ 6^w��o�l�	�)#�A�,��9>������Q��.٤��/�RW W�<t3�d��b2�2a�G>`�ǟޜ���X�%�ՙ��dGT��@��(\.gU�zV���P����ҏ�� �/��M�N65�M9hvmA��\�8[�Z�c�75=N~�()�~pt�6�O�sYh(B/�xi����qf��r12c�!��~듣�9���v��ENWo2ۍz�[�
�DW��صJ0���4��`��Qcv7 ��-�.M�\>ǽi�����,U�Ì���n�[a��e��@�'�:�!��f39�dX��%@�`��5�I�C���χQ��J>K�=��[��Oickh9!��ɥ�)F=p�%�<�f*�(���6r����--�]ߣ̇��Kz8��e�W�|� F��S��AHd�`���\�K^ܐ ��{�4Ʌ@s�S¬1L��^����rs����JLgf���Ij��oV��$wLz�h�9�i�^o�^^hR��uц�����Ǔ�EѿT��[�e���=?��Rz��P�-D����/א���O\"��D7z>eտn�H֌�ݓ,��S�"wó�B=w�O��AyL�D"��������a�v1�C�]	xxMƼ/�|�� �i�e8�j6o�%Vq�?,��$�8�b�n�<�2]�K�d���k��_O?^��d�j S�6п�	�>XR�r4��huA)E�>��*�[=�4d�����	!���
P�,0�vİ�RY�f��s�"F+��R�L��X��F��ļ�i���(M�8.���2� �3'.����Euy>m��b�o�i$a��kA�ዧ���i[3��Kmx��Ľ���ߒe(��������.��d96���A�QF'��x��qޗ�����J�Z���WRO
�hdo�?z5�q`��4��rD����vt;��u.�` 7B��@�]��H�P_/�7(^�c���[eȷ�^t���\0��
C��+P9�Fl�=̥v�bm����v���"�a���%�Ե�&m;o��ʡ�:z�]U��(3��z�T�47|��r@-�E�Γ��i��o؁�]"k�ƚ���|�$W�=Z�(`��R�������zP�-���C<N'�����WL>@�=��i�BZKRO�rM\&F� _d�$�ب8H~Bl�O`y��Z_�U�Ip.u���� �JA��V8L��^��>�ZIգ��v)�T�ޙ`v�Ke㿞�Hϖ�C�S�F�)��Gq�_��5s��o�ɭ���ûs,����7)r�sFv�\	���O�B�|d}����hR�̀Rh�0���?�x�3g����q�������e�;@^�~qz�ňW^��TRC�2޷��0����%S5i�xq�����d�L��HH�����:W�7��G�G(��R��Z%�U�rp� C:��?v�z�r�E�/���ĶB�e��/X��r{2��	�qO�'j���H�D��5=�Tɜ�������z����`'���<���)�큎t%�,)�q p��ܢ����"���ޥ��_}�:�%87��������%�	 sfFq3��7E���Z�������-<n�+u�3P����!Ʃ�l,w��.����ɽXU�c�q���u���S���gwc�1�J
_���!�c��,$�u�:�0Y,�R,�vV2{���~ׯ1'7��0مz|�6�#:X��La�s+�ADR�X} �I]_Zb��Ґ�
��rg^z甯+nr+J١�yg��b������ÃϠ���t������Ɋ{W�݌@�U��>�M�!��������=<+_ѲQ��mJ��$��X�B�����h`m��sik�v窻rh���Z�W!���ށ�D_��؆�G��m<o���L\�5{�� ��EO��ش�L�~�W���/�=q5Ix�俵�%> �D���u�v���)���[�^�!�qh�.Ʊ�[���(�N&p�2�ŷ�t��{R!�$�!����x7i��WR�I�hCs�^�0�4	k4+���MQK����O�=(���`$"�8�B/�ڸi�&��8�9�ф��MT��+ :�H�à� !:��G�2�੸jhq�m�/|8�.���%�wV�K!�Q�Q�vr��/3��������W�t�K7�٘�doj���w�%�( WZ�h�uho[`�� yb��ŉ���pD�r+w�������s�i������zL��v0����Y}lx��)�ghF{Y�_ո|鬮�`] W�]��ݖY=�\��kh��q�K��ȍӦ��8ڭ	2�`�$h��d0�w[P��)��|/�����t~�>���;�yO���`���J��by1���b۵�[5�9���U�|6��|Ҹ2�?T2�v�4'�V���KR�\�:*���A�cӬ(�ny�k�/N�o�=2��N���ʆ�q˻� ����S���z{Fmk?�{Q�$G�����V�s;iɁ:��&�d��CY1@x7TH�u���1�312��u�ʣ�J�*R��ѷ'j��3�H�N6#��o�R4B���� <A����=��%A��
D�Y�4��?h�%ܧ+���g�����O��X�t-)v�y������ҵ��N^�b�"��tޖ��6L�\4�;��Gd��h�(Z��W��������.~��9��8�A��?tY���������H�*��	�	��9W	��Hc�r��Ӣo_Ƭ�����ت�e]�E�)�d�i�پ�!�������>Q_����慦��;E�+���bwT�9��^3@�6c�k{���m>�f/����N;3G;W ��\X>��K-�f�0!���'!S�
,R�,Z ܣx�渜�7:r�JAq�x�P2.�d߬Yb�9��fK���0lK�kU�xLӘ���'M`����^s�&
�8��*&��]u���C�OO����0��U�j��Z[�L�&�|�.���v����V��H�yXv�M7#��>�%�E�ğ�69�h\Ik^�C��� ��q���~���a�z�n�k���p@]4�����y�p<��q{�"�`�q���q�
 �l_��$֟Ep�N�/��*��ĺ �4���^#>k��%;g��{�+����d,k��ķA˗4=rݩ�F�B�NѤ�m�ԑ�H�5��A �zy&;ApV���V��d6P,��eх�R�1�f:� �T����j���4h;)�bf�s�G+�͸^�d�t�ٲ�kIe��&���m,�0���_hpD��3p-����R�>��=H5\�<2�7-��[��^(~��>n�*"���ЮزX�[~]u��X��������ݚ��>{7NM��*aVR�
m�e$��ףTC�P��M��@�����0���9�/�3t��ٺ���~��ۉs,윳mt!�v���.m,	�Ւj{H�2��λ5�:ok�R�m`���mD�H��;�*�<�Kp��� ,5"��V�̅��ծ���0X^�t���c��ς�Z����l
D�����$�Za"�)�2�+��-�⍼/[m..�v�s]�^�)�ެRT�!��7�_�	t�V$�����Њ�F��ZT��}�7�Jb���A2�l��S͢�Rl����u�$O��q�����C�|��%�K*�#m@�J�S��L�#Z�K��R�p�S�D�����,v�P�q�6!��pK&HW��n�q}T֟�~j_�!�{q�(qHYO�-,���!��cW��ƃ�j�9d�x�ʰ�c��A�G�⸧Dـ�x��+��`��E8�~S�2��Hpo�zT��u��:WaZ+����n���\t�xhUrW�%���P��g9�x+99=I=�~<`��8Z珞|�H�ީ'wr Ň"/c��3��%sq~W�H�;<B��Ȗ9�1�.��1����Ph�C���6u������dE^cpt�H��o��{|�(7�$��#�]�nH�-� �v�܁cI�Ӫ&ެ:�R���+�ն{uYf�e�yTH�_�� )�6�5�*��dGR,S#�~�'}��- �Bm~3�^0��vw�~�(At�;��X�='B����b��;��mn�ݢap2��� dWN���� `,#���x�&�CS��N�T�V9�EP	���-�OS(`T~��\I ��Rc��,�o�-�H<��Dֲ9J�[p�5!<��g����0���A��dt�[p�|T�z�:�|}87��F���Ws�v>)�}�0�WDm�s�Hz5�#��"V�?��qN��k�&����g������Hc������:��X�Q(LIK��@iө�M�UJ@��Yk�haH'�Į4QT��©+�<7�j���mȰ�`�����j��P\���3,3����j9�I�����4x��U��r�����z�!m�A=A&��tA�8���x�fI���V�m��V�;+��w��b+Uv����[����a�!�v��Bj��X�Ӆ�3&��<��/��X�d�SlɎ\
	�=^=o������,����G7x��q�>��b�0��x���TmvI��F���7�9�n�� ���$Y�U*�3Oo*���ݒWbQ���+��'��9._��כ?'h���g?�nkC��7�i~n�W�|7M�j��5wj�?��zx�<���������&? 7[�IxfU@��R��~� �r��U���C_<��^���Z� �J��L�;m�����F{�2�4�5L��SE��m�24��@<��c�#��!No�_|$��w�Z?��z�WF$��;;�UqX�� �[u>� �Ϝ��c�;f��ᴸ���b�
�qKPk� �b^q�G����o3OX�8��R�V>�1�����c����c�W�u����=��ȭ\��:����/�%��q"n"?�bR8�L�p��GKv��2Z���Hɒ��e�O��̀�S��������RCT<����!p>����d�]>��vسH'H��E�Po�w�X	�P�*�I�����lx��M��;��r=�"bbe-��N�)�-�s�%��,6>�A�5��lE�/����ίP�Ż�I�F�D;̵���g�+(�QAm�^#�z�j� �^�� Ȼ�#��v����g[_��vt�2�BB��@|ѨL���h^�|H.�~�#E�1^h0������n�9�Z�i՜6�.h��U�[��L6@{�͵6Z��·��L1g�I�o:�?���ҹ' ���D�0*�#�¯�/�66�(�
o,)�Ղ0�Y�}HӢ�?[
�ҮL���\m5<D���&���c�xw\ٛ��{'-��/� ۝^���O���lvk4������p�}����<!Z�L�1;��r�F�q�����^vz�6�]�+�q�ݠ�o�'�a/�Vf����ra>l>���jE��@SG^���,����/�5sE�&�XgM�f��j�A����ª<�.�C�YL$&a��G�\v�]Ld�`O<���t�'�K��o��E�����nhdٵM���1��H���T�:P˼�ALA�&���W�����jz�vr�� �B���N���� }�2�Ӹ�K���9!��g'�1�[�j�B����ԓ�U1�遜�J�~������xf2�XI�B���i�f3��z;�����������b�g�0
{}�t�9w�� ���BJp�"��b�gEp�H��+��+�Yn<�dI�?���{ĳށ��v\�OZ|_�m6�?��"��d7�$v�K�C�;�L��c@Ύ�K��j��Άu*!*9��d���%�<����EA����HK�������o���t&L���a�q�-u�ز��K��
|BR�[�Bջג�����k6p@"W��@�F�Q���Тv#�n������،עN�����q�u��z.���֮�}R�������$�Pl��$�V<��dV��ns�%��k�V&�xzQI>x�3�g�rVu�lI�T�8�7�4�rW����M�^(���y�3EdAz�׺�Ph��"3f���%�;E��32&?�rd,�6L]h9�RU�y�t
�h�pK^yBU��{j����E=˖�0]���Q�c�:l���u���|Ov\ 0�ק/�Z�Ɵ�tz�ķ���5�`�K[g�cO�FPԫ�B������O[_�fL�l$���_�"H���j��f|���6�w�eJYGe��to:��:�˯0���{�&'����8CB1��g�d˓kVd�������L̩�c��P)n�X����BF� �����p`�e�燦���Ubc<������ؙ�Q=�y�_r^L��O�k�y[ew������{����\���݇/�.Pm���'J���8��M*��y����Q�B_*�Ҕg)��~��4�ixwP�z$��N�/|T0���@��W�Y�)M�Z;z���,<,��Z��\��,��ό���6� 8Q�d+R=�2�x����*/A�[vs9X�Q�2y�~&w{�]�`�'P�� �LN�~B���C��{�NZ]�ĐGU��i�Ē�B�m	�SS���O�
t�kX,`�|�H4����~�<�2	7�3J�u����+a|�N�c�24���Hq���?'�-�M��2���ԯ1�v�\����EC0��Xe�֑(��7��!Y�V���k�o�x}�M��i��J�⬅�w���WxY$���Wʣ��9F����=��uD���9��7)ѭ�b�@��vOn�5Y����c�?LvN>Zݾ��i5��U�SRb�I���U�O$��RuR�V���w�9#�6�4��:J��u#�ۣ��_G�����t��'ܟ.��c��Pk���GX�T~����_�¾�Th�ii�dH�Z�����g>����}	����F�=+�X���N5���n0۱�&:Km�.�cH�p�Ma�]
WJ� ȶ�/�w�V������j�O�a��g���<�\�@k������`���8UH��J�}כf!x]'�ħk��vԫ��X���`\	�DP��R��h��4�p�4-*�&I�;9���u�;;�"�]������e-G��!F���U�H�����4�P2�wO�`�] z;��p�N�rW:]�N��Ob25���s�l����:fI&-Y��
��M2�va��Ǒ�������`Lf"Ջy�<bkgo��Q�I��i�Qs!������mr���E�Y����uD���X��0�T�Y���h�hd��w(��J��:�ߒ2��7�_CT���`}RYo��vLPbr��ȤQ�~��NcBo�(����,������`�)ņ	"�x�i�\r˩�FvYS�%����ڠ{����%l謏�����p����<Tn���V���]+��8\`+-�|6��Z���[�^�#�!��Z�,���&^A͈�1�{�HLk������R�5���uE�l1��J�썀؂%�S�`�(��g�u9���,4fԘxc_&t\Q����*Ptw�I ��P�ٺS��"�3��4�xg���L���w�tz.�Լ
��mf�".+9��ދ�~�q�}���5�V��b�}�$�챑�c�t�4�̗X�r����j���[�Ø�m��&ǋ_��AE� �N��{aߕ��pi�2o*���B���K�GPF,=�>T}�H#X�=n�Tܞ�sf��s�����O�'x��j�Sv�w3Q��ib��Ųz��Tkh8e&di�	k��%�=�Rf����įe,h���Zs����`�2?/���ER��^�K������)������Y ��]:�B��_�e+J栧��B����trf�7ۦ��3� �ō��O� �n�v+�&F�s˶df���ު��AL����'U��*�&"2S�@��	+�@�FM0�^˗>;4M?����,�L�v�u`?��C��m�[���"ŵX�{�",�D^�
9�jv�q�����ҠΎ<9R�N�9d6!!p�Q)"� �B�)��~�x���=�����3*l�x��⸐�BћG-}��6�KW�7B�8GpX�{�\�MX�X�O�k�߻��ǡI����;���~�ܤ�X����5[OK��҄��@U��"��3Qi�xh�LlW��`|,)���(ŅZ�����ٜ8��h��Sg�F�3��\����c���(þl|�
J-��4Ti&7���|_畄�(�Z��ք�P�.�(��|Ȅ2S�[~���h] _��qGp7m�B�EԨ1B�d�)V���ǂ�k+a�?.ђ�ΐX��9�3�G�趌�\��meS򹓓c�=�,�(��D3��IV�^8>��Nk�/mHf��g�*����$����D�6�� ��C���^z�(�64&�=��������*1G
��0�ȭ8v6���I�u�u̧���q�=D:�r
Ո�U�̟��'�k���ʷ##���� 3���o+�T����8ײ���v z8ά��3�ʭ2c2��<�ˮ�(U��Cְɋ���IZ����������Y�Rxa�we�Fϲ�*���x� �Ws7j'+NԾ��^�1:��3N"S,���+���'!�����xBЗ;-�.�$:�G�+����[qPL��'�L(Ļ#dV�'����(�#U��_sBX�\�������F��/�}{�70`��7���n _�e���P)M!��-��ԊC�S�*Vق�"+�@h��^F�$勲+QeH-H��������؋���Y����̀c7�+��/<{)bNOt~����k����o�ad�ۦq�S�M�x�p�Zp*�Ž�轍��J�ޛ��^e�hJ�OY���QS5�:�5���o�-�雿4���S������㉄Q�/B�b�&1��nc�n,>�j�1H%�\y�9� ԺӞ�r(����gC�!�Bb&}�{��^<�Ny��sQ�o�wR��KU�H��(�K��b3X�����
�6�a���#�F��.!� ��Hv+CX�D4�L������ۧ�|ǩ���/�'y`G�˷�zq^Z`�7cS$H~F5�hg����o5���n�`��WWi�)}-�3^�<3�Gغ`Xo�5U����=@=�&:���h�C�Kљ��� ��lA�I|ls�� @���ܪ�;�[r� �2+f[?0����!/>�BeI�7���
���v���F��Ʌ��&?���(��O��W�X�^����*��~03R���zҩ� =A'0����xq�2��4��GBa��>	��`(f���h���i�y
��a{���R��	�
Hi��5y����x��Ћ��Ξ�x�s�ۥ7��
v��N��P�1��qަekgL�������K(*h&$(�f�f*Z�~Ŋ�(��Я��!�e.�}"\����I��=�8��Ux#Y��|K��C�D#���y�H�NA6����}�S��P��h��]��D�kFrƸ��$B�~O�֊�UI�nl�ܽ��T���?��ɏ��n���s��1��h�-L(|�cN�f"�:�4� ��@5O�29���:t�﹬1�M
��I`Zλ���&W���Y�2��N~>'���yL��8�-H>�5���e�����#�*IKq�H���H�re-�
�h��Pgm�����%��±{�����e�	�b�(Pb��?L�hs�2ĺ�i?�c�T�B�#����űa(@���H�u�DN�Gh��c�����]�wk1c�;�J+ �Rd9��~g��SM���&%���m(7������ma�IQ�����]f٫ULg�k����vo��_\�Ҵ����.�A-�j�?~\k������3�u ��f�8���>�#���m����E��i��!�F�*�~���ɦ��A<J�G��M����n~|����hr�o��OE9�����~A^��W��ң�����$�?�f�! �D�i�������Q�FR�����l�2?���� E�	O���D�SE�{�����_����s�(A>Z* ۆ�S�9�ٱ+�-��&����^-F�QV��+�"����TN��fPnz�(��>O<��}Qx�]!�;�����Ģn7=
:
��m��I�����GT�eF �G5�̱vs��0��7m�h�� H�k�˗�IP�����R@(B$��8a o���S�¢���?�'��)��15�(�{A��X<"���{���8��-�$`��dbo�gRT�C˄��a�	��ڇ2�lZd�k!��|s�ص]����HO�:�d�R��ް�0H��w�F�!��bDc�}��A������@TB�%���r���oAr8�w;GB�� 2�~���Uw�	�̌�sh��4�T���Ϭ�u I��'��F:������S0�0H��rЊ�&Q��V��CGR�C4��v��VY��e�߫�(���;����ҏcR���nD�h�S�aԸ82����LN������'���N����':wc��s�^�e�)�K9��7$E�Ip�����,B����ѽ�Ӧ�N���ބZ������l�e�I-�	7z%��DPT��>�,ru���rlS�&)"�V��
̜s���%�*�w7�O6B��dn���=2��g��CI;o��i]^��
�͜�&���ړ�� ��q��C�`�2������S�f`�GǇG���ݲ*+%E��@^wm�H����+��U��)>�@���f��KO�5��7Ao�l��j�6T'��z��ꐗ'��";�$����P ����+�
�������۵�|��Q���4�4/<1�R���b�X�>,��zfv�D��/��d���W��HO}j5g~�q�=�����Đym���/��܍5Rf��(�:�6�8x�)�
��I"��C�@�e��&dH|��e���6�(ΎM)+��s�Rx�2",#I^(��x��<C��@Pn��n�ʑLlt'�T=ڠCJ^�����{L�I�Ce�|@ ��W5?�v��:2!_v�g	�>����9`}�wVqW�7�+�`���2��y/��̗��U��1��^&�g�-�{vN{��ll1h��٧��n��yш8�E*����ڕm����O@�QsP\4�qDN�X�}np�L��?��g%���ނ�7��υ�f�&2��si�ݧ|�'�.��l�0�4h�&����v�
�e��A"�(7�J�'���r�=G[�?�,B�_���=���Al@�އ"�]�`]�v.u�M�&kTe�2P�)Ԉ�����Q�5WԐ]Iʥ����<i��� �j��X�%���~%:��&�����J������l��_�������l.d�5���/�+�"%䮶�
���Y#;`U8T�I�>̞���g�8����Ӆ7A��q:c�;�v�A�޵�~5F��tMA�/ӛ��eȸ䠩Q6̑J�s7i��(�Ž��}�1m@�F�x0��+b�e�2Y
���b����|ƨw&�<қ0���N�0
��C�{!�<_�����p��n�t}�KL'N�-)���[���"e��x^��O�Aw(w����ʢ��lhRp��2LC;ޣ���AA����,�����\�����EqԲj�����_Ej�_M�u
��?���R�D�a%�;�n3� �wA;�g�{&K��]�z}Z�����)�� E��`����,��dfO�,	���D� ��ጓ���G�wV���.s&��!}�R���i ��7'�)�/=��Ɵ����Kb�+����u�+%�=S ��d7-�Q��}@gu���y����u���4<;�Y��'�����v��\�����n�O�!N��B�P��e�4<���)��BMgR��\��2���&�6��g�8)�h�D�H��Α�vi\MC���r�?���Qmo�N(��{oG[�=��>eq����if�s�^yxɤ<+?����P�Z��xo�R<K���T���~I0��@g;��nA��ķ�+]@r[k��xX������4�?��R1hA8~|5veV��e��D L�MGD��\!�4����@���+1�����e^���{����y� TE�$��n��]JH/��V�����4�# �Ki/0L�!�W�����*���	��/��#s�n���v�m6��G�%����JE]����~�p�X�A��4.���
"���g��[�9�Џ?�D�,���%ٜI�d��a�C!��9���i�����7��K��w.(�#˯�#�}f�LA;W�N6X�f$�!sP���:�-53J��@V#34�!��7��s�1+RƷ�	V�dP���»��?�'>��F)�k(��{� ��"����"k�Y���9�j��} �5��Ȼ�AC�Q��"#�"�����c9��$�vIhwCY�Hԑ�zO�W���+Ѻ���Fj�)���r�}O���<(6h��U���f,��/�<�+HK�`k�.�/T�W��$0ݐ�ްQ40e����>��zBG5��,��R��m����E۵�?ݎ���Ҿ�fO�Dxy���I�����\�%煮C�\������Gs�F� !`��>S#�4�U�ai��
��,8�-�01�qv���8��U�����W-��94�m��!Q������B��1;L���vb�t%��lS��`D��5�W��L{4J��R�/]"�8+�h�l�z����N:f;F�]@C��o�G���d���z�k[�r<����c[���^H�}8y�f �|�i	Z��HˏU�`���у����H ωV����r�{g�����~қ8�o`�7Ģg�d���&N�M)w6S�� j�=���tј�`#�[s7z�S�Q;�9�:~jZ�n�[��� �y����Q�o	E����o�l�����Y�ď�p%�zm:O	KěF�� ����\����e0�%�N��z����w���V����{o��2��ThΫ���Lx����t�E�Д��M���5�D��V�6%��:����n�_�%1V���BJ���}�ÐB�8Z�3�9��KZ��~Jg4�.�F��2�(��p�UH�5���YH2P�ի�~���ԩ�]#�#2��������*�<��xnF?#�6R��DQ�����[���!���N=Պ]�y��Q��C�j+��3�X���H�}�^^�7�o�/��E	�a��8��F�GTI�W�u��&���9���/÷Py���#X5��c����͘d|��V�lP5�֣��5���G���}=�y-��xN��U�xW���琒Z
��I�L��yS?#�(��+�l��."{P�H�����`���>�pa�w��4�P	�N/���/�`w�{��ɥ<!E��)��y���`��V��0�p���d>��/��ò�՚�pP��5�*�wL��>l�*SB-���J��D v�E���nD���-���;��d�����f�4�iE�CMHMK���4.��[��ŉ�ɇF[� UyA���{�=�;D}d/��$��`��*veu��x>�|vj+Xu�R�ǧz�iEЋ��U�tj�9/��,����:	��)��v�@K�c��h����f���'��Q~�*,��m�gH'(�ng��v�2[��O�ЀǦ�Ac�Ylۖ��`���"G܊�@1M9�ǁ�a�� �̬v�rM��$5~5|��S>3@����s��}?�Xg�9��>�� �;'HL�'�<}�(��@�vT�yy+3�:s�=ӜU�Q����K���A���� 	�q�P�^��9�!�o���1�g�sG����Qt��଄f�ӌ*��dt�e� �Ʊ6׋q�Q���#$�w��&�������zS�u}��W:��wU�ۑ�H�W:�1w��#�Ǒ+���|��C�6��������W���<J�Rǐ�WںS�鸥!0�
�\����~��c������E_�uZM��Rl��ȶ�,�/�u9il�z�H����l�;�H/���=��~S{l�n�?��*G�@�m��Cf��ؕ\˛(̂�������}}�}������Ԇ������~��q�����2u�\��t��Wn6��~?`�۳����=n ���X�C+҇czV$�z��:�s��_�[�w�TI#���6�修wFۥ�@�N�^&����<��Lb/�r�;/�y=�M���JR?ya�B��1j:]��o�� �����(��fz��[�����n%�/���hH�Y�c��c����<ᗀ4u������_����O���.q���y2���|� �/��	��.�Y��#&4�B�~�J��ۉ~�8��Pr~��m/��D�p-}Ul�����#*E�'����S*B �8G�u}�����c�GY*�M�f=~�-]� ��5�˽B6���{����&�z"���c�4�H��$03c�B�F6Ш*��̡�+E��l�L/��~32/�~pt�q�6[�������)���)&K�gm[�4Lmn�����ŤMO�bvMe��ce/�3���/�M�n�i>���[t���65��0��T����D1��̖��^{[�#�C���f��)��ӻ�I�M�R��%��,;��KӭAr"�UP�~����ġ�~_^��́q4�9�t�W.�n�W�,ޚ}��3�ta����H�YQ�%q��#�_���H�c���k_�p>(Zi����f��S�m�������w~	��\۰�'�ĭ
�>��}m^3�5F9�Eb��s��;���X��Qfb�)���X����}Y���n냞����j�y�D���s3E�:�m⿤^c�އ*�`;�HL��Rɖxz�ݺd�pt��]3�W"��=����l����A1�BE	�u�]�SK��A6��ƴ5/F;�ٟ;l]�҅fXLF:p���T�]1@�q�	�j��r��H�&������1�`t�s>MjRP�Ĉ%�D ���wdYQ�]T�M���\D{p�!���%�A���L1���	6��PWՆv,0;Yd0j{C·z����m����w�%J�#�p�|���n� �Λ��� �p�i��y�~����?GX~��D��q��nmzd�ce��| �w�����Ay���RU��O�Z���H���g^��qF�:}�t6�f_a�GT&A;��Co�T�v��	[�AHf����R�h�GL��2V_�}�V�����u���l���Y��L�}�cH����b�k�'��n�Et5mඡ��X)������NS/�&�o����Ҡ��[~z��PoO�rU�S�o���q&�w�ƴK��Υ��֋����G�q�)�Xx��iu�|�%�k�ݮt�'�RzA�!�h7~>7��Q���	K���~L�i�d�5�Q��o��3��񿀴�ֺZ�~���a�q�h��.&���5���Y�r#Gf仍�XG�Hz�Xzy���IBoW��r�P{��U�����s!�X��aeF&D+�G,����z���*'Hj��_+��̜S�������+�L���E�P��� igV���^�I�f��!�N���e�����W^��
�f���o�~�k�hΛ�,Ug��З�^�It���f�"�����M5�����&�%mZ�vs�Z�͗��Ꮲ� ��D)�0�U�b+���{8$��`�E�c]D
�d��?�_��&J��:�a��ve���R'��~���T&�࡛E#(X�H�"�!i�~���B͙�{u�����7����y���F��O��fde�ۑ��X���<����0������u~�(�Ь8�S��L �L{����\u��4K��ke�t�u�������F��8){Ă�'mȺ�#$n$�H�#l��S��P%�[HxKg4H�w!�Lr,Jo��E��@�v���@a�0R�����5uT��'q۩4�68pޗFf�C�"
�saI��{�)=*%��%����Ӿ��my���,��S\�+Cs�  ��3�;�T/����Iѳ����3J�����#�޺=I��V(������s���g��=�m��I'�D/�0��&��ՋnK_�{�!ӦT�ujoV�ى�Z[5pO���3�$��BTY��x��>XY�ᝳ�CC��-zI<*Tv'�TԐ%�O����Q5�1.j�.v>h�5��]@ަ���w�J��4�ҽ��J_��H�"�1ۍJ-a�!�U�@O�ޒ��;�(F���x@�g����e��#�oR�xv�2���2����%ޅuB�Σz[��:�Ϟ�C7r�w��Es�o���q)�	��E?>���^�'���^����>�"(Z����6��Lr��D�@$��[z럁l�́-mΐ�4��|)!��EX�6r�$<6�Q:9.A���Q[qZ�����s��ɢΌ�O~��fa��Cy�I����]�bSfk�^�����s��u_�����U�-���e ӗeF�͑�Z�8di||��M���e�̳)D�1ao$I��$��s�N�v��ٱ}�\��zUkÙ3�~S�wA�À�E��MK�w`z�_�h��J����w�7	�l�#7fx��~zC�`�s5�/��B��=`?�Y}�s����,yn�,�t4�>���)H6��	)z��Ղ�G;��-�/��+�S���)z��@���ܘ[Ϳ`�#�Zn �5_�����F/Y-@���v�񋈘?l�6�6��'�/�ל���'u�Ef�h���P\C�p9U �UD��T���.�ա�l4hY�R<��,���:.���~B:�;�eKV��j�o�7����{-�elhؼ[��ʢ/T���K^M|7��b�~��]�@9j�kf����)o�P~��Ic*"���v��H��2Rt�)E+�Ya ���nD�a�5#��Nَ_�E>d���r�U�� <&�탶�%�����6D��u�;:�$%R�6�pq�N�--;]�+�Ȥx�%4��Ĩ�N��y�Y�O�f@̕�=%�����l��(h ��%@U���'~�0���d���q彆���񍒉��m
:�����4�CN�
w!!�Q33zv�81�%�+���n�O��YL��;�T�	�SңX������9��vH~���;�����L�Y*��*	� ��8.�I�0��r,�-	����
p�O˿��]"d�:\��ed�"�\2�\�H��ƺ�5��߳�7��r�aw'�C�[p U�ss2�m�Ȉ2|c�o/&��j ���>2�2�¶�{��~�EFbsTU�
���z���[�\HS���eQr�_8������4�$�΍�r{=Q"��<�Q�m���U�g(u�s���d_.���u���	�!��A%���/�W�����yӒ���\�f�7!�gl���o��2��q)r��e��H������!#�_�L��R�}�������܍'��X��b9��R�*���Yл��� @<�F�kN�)��5E�������ĺ�V��Sh5GU�����T�<���H���$v�f�\s�a�HugX�%U!v�YJp������󳽣B$�-p��D��CX�O%��g����cyW�h�C���	
l����K.j�9�M�K��ΚY"���.�^��7��$j�1T�If������� A�&���?~�]U
""YR��"c�f觃��-j�l�8N2vP�T&����r�Y���F�ƾ�{XյR6L&Nt.�(����û�D��S��{JE
3]&�Xy��k/���UF�Z�Ka���Z�� )�<�R|��Cd�p�`�S�#�T�~ِy����'�i!�ʭ��!�X�2E'����Xi�i�[�-`X>��sF�u~��O�t�yƓj�4���QZ���u65���T��ZMA� ���4��c� i�d�|m�<�_���K���>u,�8ʟ��i�����s+:ϡ)H$�la�6�t����;i��8�3K�,��b8���Tc��ө�D^��6# b���G�B�>qWx5)�)��%2u��ż)*�Oٳr<i���Eg�
�j��8�� :�b��~Q	���k�"$ӵ{c��\gX w�O��O��C�~�I>��������T)A���v�ϩ�Ѷ�Dr�ȷ�A�Js
|�wG[;�=�n�3�����U-G�.���{�ܬ.[�0g'b��c`iG�Y��x��������	�T(�C��߉��ȥ���j��(�G����&���1*��NG2N^��x������t�oQxE�����*�
�w ��ˇ`�]g����b�d�)r��PZcje�u�h"����Lg���6X�$ꂼ� M���O�g�۫��V�>&�;����]c�`
�
��ԛ2b ����%ӯe�� �8���=�L��8��ῠ�8���������&u��Γ�;4��T�
6S��A7�#����Uo��ǲe��DI`�|�ސ8w�, ���.c2�])7eP�����CC}oI�ޭ���iѧ�ό �NYi�}�^�`��������ںڹ�X��q�8}����g΋OØV	- i �b:���Id7�(���л@���wl�kh�ǖR;b5z�&'f��*�fK*�#ӌ!�y�O���/��%̈́ܝ��PK�}aUk���lȅB[�N�?����Tk�F��Ec K��e>����M�3���A�
��X