��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|e����M`p��ّ���Ұ�Y��&�^�y�w������\�Hz���Xp;r8}�9���6�v�ZJ��k�j(�uK `x������#�C��2��2� �j)�8l����%�MQJ*%/�z9�w� ���:����]z�lI�����B������.%a��Y[�BKq*$� ]���}�R#SDQ℞��H�أ+n�m�V���aڒD��'��Z=l�Wcz|;���7Rm�j��&~&��\��pzl#���5c�b/�U/湐���&���.Um�'��FD�7���Ih�d�b��/��/Ġ<���73,����*�%\L(pv��sv���h�-����*m�p�x���<�q�IP �ҳ��C!pҫ�L�/�m��*���1~�_���P��?Č+��e�����
.�+����b���eh�pJAԙcD�z�R����4Ξ�lc���4r�$�]��#k����:�3t���(T��[�/���/�q�Vt�B*�gN��X�m�-I��cf&�Xa1�FJ|<��T1��Ε�לּ��(ވ��W���?���a�2��7�W�B�LF�8�k�4Nw�? *b��Dl�Oxj2cL��CCޑ�&��h@X����S������L��"=�����m�Ϛ�&��jgF�{=�"��b���Vc���d(��ʼ����ˤ1��dN)�ӰǛ�D8_m��`4�2��N/�϶yٛ5k�^`�Z��� #&�ԫ���i�Z+E���(�1F��oJsg�����z�	cO�/3vY�����\ ���u]���p�b�dT�HLj�@�;um%D2�As��yLv�>��m�z��i�� �f͵�T�Ż�f�:5ə\��*X.G������N~?�W�k�(�$U�Ҁ�(�
g �z7�mPҚ �Y4��oV�.%�#J�> �'~Js�v#���VDڳhPF�f���m�Bs�c�W9�a4JyP+���5����J��zF`��d2��7��} ��[��Y᧬�]���=X��Gs�B��
oo�Ͱݼ-_ן��O5�Ż>�&�8?�-��Y�����٪;�Ә��ż�V�ٙQ�^Q�-*G8Ľ�)�qڒy�φ?�p��-��?"����p���CR�)�:�IYpƴ�	��=vE4&[NpHr�F���ۤZ@��*7�*��^/.C4]$��`&�e�$_�1�ʹ���o�"����}�a*Gs��J�	h뙛�� ��	-���;�1c��5��KZZwʛ�M3�0jR��%{r��V�­D��$z����U6�X��?����t/��h�	��-v���%	�и�	�� �g�)��Wȼ�}����u�Z"�0j������}#���G���?��>�lN�z7t������	~�c�BA�(�;u�+��h=C�@(������2"�b�盷IW6����8�m�~`�[��Ϡ)�g�;垿ֲ��8t|}��w��ʰ�hpC��szY,�KT$Z�|n�;$��ʈ ��Q���Pb�zω6:c<�)���nݨ2�f�Y�ڑL�	��7=8
W�8��n?׿BR�S*�4�������&�D�v�!�"49�_��'|r#���n�sZ: ,�p�C�dKl�.���{9�����̢�y�qOł�2^)"���>&�j_�����]���z���u>[|e�7��/q�[�E�9��ȀA	��k�7	_�;9�V՝7�+j��R���^�l����Sd���M1ǐ��A�M��P�*�?H�<gW:���5~VG|�NFh[��|��[z��ر��<?\�8�s�R�链>�WՉ�9�nhh.F�CS�0���4�s~	�,� �Q�[U���#[V\
\�칪q���@4����|�6�od�:����]̘-mf�s�X�C��B�jT:O+�&K��b�����yL��PH�p�	�q�:�!7'� �v����������}���@��W�%�߆��3���&S) �a����)c�ӦM̗��!�y��� �`%�\��ˢ7��3l������sn#��Ͷ0��[Rؖ�{��İ���H0X�Z�u��ÊO��g��z8�W����П�1��v#-�����,io���]�s�"8�+������RF,���C��|�S�[����(�L#ۍ+0�,�z�J`o}k�f*�΢��$1O	~�ӿ2|�5��m�`�iO��*p�ej�a��H_�=��$��Kb�������e!)��GaƋu��R2��F${�����8����ΐ����B5���:�lϭזu���[r�����)����p�C��81�$|J�(�?Ǐ����jHʶ2�Ż���IK��������،��묆�6�u��8��a� ^\�:Z3�vL|��6����}�<����ם�I���`��N_|�^JWV�N�
��ߑq6��#$94NL�t,d�P�fLJ,�9(R���,OH%.iӥ�����R���.^	S���N���,y��޷��w��)�C���.�Uw4�&hs��#�?T�G�dycmg0��Z%�;%ݏ^���.���g�æ� ]s��	�R+�w]�##f��'��!�/���a_O,<pF�1
����A*{��ʑ�ORE�ޢ�ڴm�������E=��=u�sp��n7�q\�� )7���~`y��4�uB�̾3H������ �O_$���/|�6����M2� ��Y�q��禨:}���l4�Ĳ��84:��ȸ�9�Ṁ�(h����L�?~/}�Vf�L�x{Ut�28i�J���f�/�W����x����AVi<Q ��p�)��8��5a��X2�@�W,-�:�l�������(��^�ѱ�"����|�jZ� �^]�����ͬD����5��KLo���5�wZ5���H���Y�M��F��^۽|�v(�zl��~�-�۝&\!C�'��gcg��ut�9���/�S�	E�T�k�R�"�l�>��5+���ҡ0�G*�M�cdcR->���Al��z�q���P
����X@aW����`��<��W=JOwy	HKA�'�gl���bd 
a� �&@}�.�v��w6����=A�V.�{���*V��ҝ�n��	\�^*'�E�IpM�]����ef>Y��@����>t�|?/���J#9�w���0k�YC���P��N�������?`���CU�`�nڀ�l�<v��q�.&j�f^��^٬5ܛsh 	�1,�4?*EU���Q�n�D>�;�x�� ��u����Fk�8�P���0��`Ĉ�"	M�(��Cƞn�z�fDP�u�op�۹�@�%�'�X�>j���&\,��`��z������A�#%9	M�Z� �%��?ܗ�;71kzSA�)Xv��b�<0�rN�κo����Ԟ$�N��h�*ģk#�n�LGu�E���Hv0T�[�wm�NR����h*Q<Y\��9Oә�\��J�2I�Q�~��x����[���̣������3��T�ό~��N��K�^���.|OJ���	,榟v^H銓����*.0��lnk�8�c��|�������I:�3���9k��H�O�+E��vC9�y{ ܌ �
t���Z��jNӦb��k|�v%��q��c���H��df����:���6����T�5�q��ե}�_ഋv���dN�8��3��hI�(j���(j6�s��e��ֱ#d�sIW��$(��v�6 K� �_Kjz|ll����W�q~z���Cd�F
�`��u��/�]��w�/L�k�2��fqȻ1��&��a��K�g�A�Lw�
E�ш����.��C�hB���24)O�T�Ġ$�B��j������P�PU��~h��M��XA4�����#$f�t'UD�X��2ML:�p�0ۣ��8���)�X�	�_ H�JyLD]F���v�K+�;l ��RX~�R�~�*�e�.V���x�L���I����O�-��Uyt�J"��;�é'� ��9�=�8�
jGoԢwt�Ͽ�ˈ��[C�i0�����8�Һ5`Dp���^P�[�E�σM�`�������]SoN�Q�T�j���ފ:Sx-B��}��z���Q5�E�i�V+��!���w��� ^$�*n��v�����ϩ%�Ah��C��62�m
w�<�$`Z�s|^����]�����џ��m|���X-��D�&�r����=�Fe����M�%xd*j���\;f:����ű�Pd�n���4�̉�on�X�"��v�E�mL�����y8_>Ɛ�hA]k&���b8:B��x!m"}���3��D��p�����)Q�8���%�P�7jB�!P��س�j[CD�z�!�L�Z/�U��2�n��>I�8?M����q�u}T[V�x(�o��}C���窸�d��(�v������=���k�?fa�)��ˠL�^ɪ��5k[~^��(�e�)i�r���^�d����MUH�P������ �&�wU����U���}h�D� ��G��v-�Q;��Х��ȁ��?'���.��D�O=�J�����	e�B�U�!2�^�`���Rs�t5:�h�n�G%=]σ�a�c�N݃��7%�����T���#B��nd(���2A�;?:�ƀH%�χ�ߍ�G-�e���oUG�m�\	�&�.�deTPb����C����y�������.�1�[*�{*�$
n~u��Z{M���ƚ���5�Sqd4 ms��/ӗ:|zx�;���z��͒ N�Ӈ�l� �q��01w�KY!��t,Z9vͷ���E�`֔a���(�>�����:���g��4C��*�֣�
��,�߻��o$���u�E�b�T������$r.�-	�� �F&�Mal�[�vw�c����<!4]���PE0��˦f��@]n�{a�s�J�]>��r��?�=fCeم�Z��v�U����y}�ǤQ�yI۝r��ڳ���>�+����g�:%%L�D(�����v� �\9�����W�FK�����!w{��b��O?h�ҹzs�?���m5yT�Y��Q��#q��E[eV��Q;�2�0 �-7o7�Wb�ϞӒ�s�C_ �JB�f�Y�Z�#�)c��]*�EX��9�>��ϑ��ūa@�őE�{�Rlm�qT�GPŚ-�����A,]W�+��PX�Jn� Dm��e���8[2��<��=�cAa�ՠw�î�w��	�\*���ɼ1�;�(IR���
�v>��Y�v�<��)�	#Jf���E�Asz`���|2N��������,Z[X+$�^{ǣ��:v�J��P�Sj�T+�*��P̑;��{�/�Tf�Uq���u��w�tr�ِ-���S�[�t����U��m��9�މ$$� ���,զ_ɵ��cܔH�1˰����c-# �۰�=�X 9
/���?��{Ȋ��OF*K?�.p�g>�#�hh�CN�eVC����
�Y���	�n�OU?M�m��|�������>�ZD+�@Ǵ��	�(�{�vr����1rO�Z���`���EX;=.�?Y�s��z�>�cP�NO�gV/��jl�Z�n��B�S��+����X�	��1�ꚜ�8�7���2:���:O�E?׬y��6U��	nP��ʠ���Ԑ-º�@Es���e_�/
��T��H��B;������AG�Pe���r����E��ߟ��6	�p�-*��ʨE,A��e�+z���7v��;�	�(�^���-��n%P��$!u({H_b7ͺky��]�?�1�?�A�h�V���b\��D��\��2F-����>>���65��1d�5���m�/F8@^ۢ�.W߲��j�|��mߔ��R��[vA����g�[G��g�,,�,�[aI��(���nOP9�ߤ�/L��Y2�/4��<wva�'p"3X�Y�<Gt��M]�n{&z�;��l���V9�Ңv�^���p pO�"��b�+M��ΰĦ#���'�t8���W�����zNR �L]���(o6~���C	�\=%�U�u��(_f�N������hj(A��2���\-�� ��\֍P�����q�ƹā��l��:Xf���&'!~�%p�l�h�@ɱ1��뉵;��c2��IH���UE����2���0�8\��J�c��i�д�����t�Y��Ǡf�b+N-�s�(ʮ���J���hs@ka�;V��t%�V���<�5'Ӫ���w�5�P���8������8 �g�YZ�9�y[7:ΠZS��.��Z��0����;��Szҷ�(2�W��k�'�g|��5�<AnLc� ��h����؃���J��m�<��s��$���M>�.����;�U'��9�0��~M i�a��0�uT}�cd� l��sCp�-8&�O����ݥe��A>��#�*��t:����͉%U���kuf㸎����59�ot"H~_
�͊J��F��c� ��G�P��LD�e�M��=ߞ++�D)P��P�'^�g�S`6��&KT7ri��Dؤg=~RXؾ��C��#�h�/�g.5&�{����� ~��lx�!�$oA���0��C @��zJ]�'%�na�F)��P�(.�	�Y|�XGc=98���9�Y�"~.�n~���1	/O��e�bc�n��<j����vJ%;��æ$X���Ej��U��3�F�[�_(a��w@�+?�QĎ�0��l]Z�&��~R��#�H�k�3J�a��⫭%�fd}<�S�UúXm�(�eN��sVJy��\w�,I��}��CJ�Wx�5�|ȩ��1<S6���ӯ�vܯ�C��O�� �ޥ�V���_�D�D���'<��MW�o%ncO�Yh:/��Y����c��PY����Ǝ~�z���C��̕˩1�{x�����r�Q�;�c�Ů��֥��5<vJj"��`��k��F����S)#��u~!*f�f��]�h8_O7|�æ|��b/{=�Ӟ�ZqlF�s4� �2iT�*R]D��0�
<F���$
�0�0K
Gάe�\�/�=�B��4��J�;�ێos�7Z�067th
�q��D�Sϥ$ԁ�:*y�����{8��u��UE�[��0����N���)�<��E#���� 0��:��Q��.,�f���ƾq1���x�;2�3�C(h�f*Z8���w�Δ@T�/7Zռ����	�2��qh�O�׬����Jʏ]�y�b�E��a5�~d}�~AИ,�lM*l�>C�o�7%�r���[���ț�-���Lq�
������y�U���2��	�y���еȋg�U�Q��wU�%/��tIw;�@�����;öJ@�<���+&#�10��k�%]�:)�Qjl=?<���\Κ�l�Y�q���ISk5����BO��xz���\Y+��C�ߟ����޲�F��{�"�q9�V>6#������g�	?x\^��1��A�*P�rdܶF��W��Ta*�y匝I�6�R�x"��ٌ�ZC\�T\U���ּ* �R�7;?X����U]��}�
��fГ�ș(���,��-�*n��;kwD�f�e�"ߖ�����|����ڱ@�:kcg8���/��g9��p_�8�e��E��N�pma=}�8՗�]�T�����m�#�*D��]/�C�뽎u�J��zИ�&L�5�p�����4�Y��i����I� mQ�&L�G�������'���3�a�Q�����p�.go�"�P�Y��6LʞF��q3��i�K�	�V��V�
o:ms�}�:P��fG�7FMY�d k`�r>�:`��O�U1�H���ņz�5a�ƞjU�^kY"���������l��ٵX��e��$� � �J�«�J/kK�S=<g3y��R�z���U�Q8~����f�*H��xl��G�k{Sy=��v���cH�0���g^/f�+��<j�&���(�u��8�Z#n�;M�&�z㥸����p�+![��N�ߦ��X��
;5"��P�cn<�6�e�X
g�ìF�R1Z��Y��xA��O����m��ġ����%<�����>vF��H���m*�A\�d$2 ��i�"
���|�9� �$�����&!����rYA4��_��z\/�9�CH�� �eE�V~�7�"�2yf�P�E5��r����g�1�spYZ���<���'eK���y��=-�����8t%����a�mKNZ��u�Z �+ .�����.�]LU�̘��m�5��pL��""J��|���|u��٩�����˚�?�q�?���I'�g���N�M0��p7Lt�DS�N
��'o�h�V2��%�&נciŬ^chz�L�4-�iQ�NxǞ�{�-uɗ�t瞨{���m�y��#��d�t��Xx���fJ���8�� 1���	�~���fm���?"���ِ�F+����,�n����c��$ԓ���$[aC�v�>��꧙�#=�e��>�e������v�5�\W�t",�O�O�P��ߙi��߻j2aA�R1�����X��JB��<�kaڝ$Uw� �d�|7ַM�씞��elD'��#����3	��jE�Q�CH	'm�W�uF-�F����C��t�pۙ���J�-�����-3)v��)z�s�[W�˚����)��jj��la�P�U��~~#~�'v;�	�o-[��0�^S~�g~��y�	��S�g�.��f��ˡK]�݊ӽ�s���E��3A��@��mtA���pV�#Ed�V���̿1����x�!#y�y�(���uM�uWZ�Kp~�����E~LJPSծP���
�0�H1��YTʚ�R���"��&R�ⱪ����!��L�1�o9�VW�.@��r7M���
�'j��7_(_�֗8��������o�9�ɖG����0��!m!ǉ����j�.��!��=�ydE&|ɚ��V�j�-��x��d��o��y�ep��A�ɝ5ﭛ���~�ҙGfno�l�5�M
.�"�x5���
����,��!ψ���F^#3�O��_���=+�uG]�O�����5�+�� ���/�,�YɯW�_�F����%����@�m�D]�c:&&��T�x��f`�T�M�66��}��sjx.�;ݑ�n�^KkM%���Ѣݒ�2�	B7��S��?���!A����
r&�3F���Z�P$�� �&m�Ŵ�boM���<;���1���5���|��!�~������8=ߧ�d�6�N	��F�()lc���_Ϫa0%� �4��7	��P5��FSy�k��yPY���.I�g��-��7�&�W@�,1.w�۔���a�:#7Kd�	:o�ݮ����s&ͧpA�ch�SA�Rc��a�u��x�X��������ԃ�#�M9���}��|���e��`?�Ak���V*�N�K��#`Ȏv���:=DVB%3ZVQ�Q� B�F6g����Bfd��M�¾�O@�^8�����	��ْ=�rQ�L� �Q�j���y��@�O���B��|�p��b�"'�@e��hsV~E#����,7�_�T�%�/n����D�`�����L��l+�<B�y�$�N>�A0�I����*;Ze�'{�����-& �}{TC���NΆK^�Dj��Br�)��얣q�f*{$[�M�߷���dǆY�9(Z�DYNl��C���lC�&�U9E-�.������w*�[�����u������T[b<��:L"���i��l���g<R��F_�eG� lZe���\J�����$v�՛tnIӓm�����6b�c�В��R��;Uj���.��H���I�p�KejU6gd�U'=��|�u��IH��z�ݎ�dW��֢Tѳ/9�8�_���6[�u�l��}�@ҁ�+pY��4F� �wo�o��`Zz`,��%v���>�"�(s�8�!g�DZ��a6��()�s��#���O*�(EP�0М 4> �����!|,X*<�`%�Qj	�K)2}�W>SgZ�"����j��"�<�+�ZK�˴��1��7�$c�~�����;�je4��%�-ఫ�����T������j�����;1� �{3q����v��d�8�O�T�@���55H�7a~���SY�pue��Ϝ��YoP�X����ˤ�r��
�]�%�D��hIb�;u8�O�]���F�7�	pwH�X��Tϼ��c|��H�b#�>�K���m��/K3x����Z����BQ���@��B̩RJCM44�����%�ߗ`a���o6�$�����o��!�\+�] �iM�#�E�*���V�G6�p(��.�Y��;���9�O% �b��|��K������T��ԏj�&`��=�	�6��.o��3w���	*�J�4�nnN��=6��!�Q{�lU[C�?|Gl�z���#_���O��̵�E�ۆB�x~�=&���D��%�@����-7H�q]���'^�W� ����6�ÎU�����6V���2�8#攄�(�It#k�		�ʪ�rL���ߵ�w��c�m�3��06�����ڴ��/S^D��� $fC/M�XM),��a�5����=���O$�1�ۦ9jq|��y �!��%����3�@ȁ��g����E$��t��o4>�Z���ǌc�/�&�59���c�/ #ӐB�����-^�P���;0猫�-F��(F���lZh�����m�'�9�YN�3G|␧b��S�ɯ��8�/I�9�1����ʁ�f��g��r��ͼ�MxCO�n��SkgbL2��n{����Q�����O�yP��@J����|��!w��8$^N�&r�J���=��Z��o�Z߀�$�]�P���l�.k���r��Z��X����H6��n��"�8�h�57��z4t��{�try޶��n���ײ�8�"w�]�h�Z���Q���=ݏ�P�Y3}��C�p���V,�*��	�wKe���$k���R����IF=E%?���@%�vA����~����+�A��Y�Ho�PQnz��eQǒ3:�>�� |��n�y�Y�	du��oS/as�pӬ{n]�|zҞe��D>O�
����'���ջ�jR�"#&+�N3 ������Y�,��ݐ�Y���m㢧p?(`�r��/�Oo��	��5����k���qx�\�d�¯�`9i�I��ν���Y�K=��W.��y�Ed��������t,��؛�2�Q���Ň��#��&�Zˑ(4��GԳKW�C�N!����yS��_j��{㋍�RU6����X�k.6�6�d�h��ǴYԆ.�{p���*�K��77�i"V�@�)��1��έ�^F2��vp�(k�&�~�k���Yp��Mә����L̷���&Λ�i�����C�B��a����/�	�u^�Kzl+�����${8��4]�o{�A{�4�A�A����xQ{���'���14�*��͙oKz��g�$Y�ƽ�?Oש�����;��ln>��6k�Ge��L�~{6<�25,�����_]z�O�G�
���(o�G���c�=��h�O		O�Y�gJ
���H~bWw��H��!���3׹>�� 7�a�;c"��_I?�[��Vx�'5����
�upO��"�t�zbut��!摲�\!{UYk��<p���ex�
�cU�hdW�%	�AZ8��[���b��&�M�/�a�l*���2�A�]�;&͂C�y��3dbnxM�~���?��6*�\Q�7E!�Tg!ܠ%���udǛ���7�����L��y�>`3���6z���q��'�h�Q�uC����|BdO^��.uN4�A��@�#q\�f�P-��T1u���L��퓴�-D�8?7>hK<Ȫ�zv���c�K�m��c���|�X�No�{u�mJȮ�>�؝~eV�_Y�֣j7_|��Í%P��%ͭV�͹g��J�\�v���񯶫��l��4�(��0�^�&����]��؞�Ƽ��)f@$�lvq�&�'E+T�c���'(����������L_1�.L�-YL��Q���ʴ�x��;q��\]�h&>�_5{w5�v&Ř�J9�#SB=�߯��J��/~"��X�_��ORG ��`��j5���>����*UЯ�`�պ��.�$�Ɍ�m6ƒI��!�n���8L$�{14�umC��yi�7�|*=�[ƴs]�W�т;����bx]W���/��#
b�0��[9��lAZRr(�F"��P�@ulW����%�:�PEd���bZSk��P�hL�.���I��������zw:n���� ���x��\= ��1��B�
e����ًq����Lc���C�<�/�߶�!p��'�3� ���d]*��s��e�4	΂
�P�A��w6��ĉ)�)�'�O[��u4	�s��\m���5�f`$�������+k*���loK�l����	�}0�v{��\[Zk`��W�v?�y�Z��>�Ao�&��~J��T���q�Pڦz��X����|P�4-��S|�pC��� ��Ǳ�c���Q}����._� _27T&o��������&M�ϊ)��>�w��*&#� !S���/!ω6�	7��V�eC|�c��^�-���}�q�X�g���\�3lC��6�Qg6����J����&Z�(��%z��@��d�a��#���*��<�OS�uwy͎��0��� ѾQ��~�b�,̜���f��:V���T�d\H��A-P��r5��	�r�u�En2cn!��9�鎇i~�^>��W�C�Y8�.�[�� ^����$���Hpk��V� �&b�WpḎl�V��m~NPBa�Y��do:n�)�7H�)�ϖ��v1S��?zl���m1Ns�2�{�BPC��gC��唞^�q�w�$Yizy������˺k,:����E�Nn��(�eYvj2o`}^��*l%fC_
�4��4��{�%�d"CZ�9�Lћ��z�K����7��Isۼ$�z:��@K2�b�z�b����8���ٛ��t��̓o$]¥8GKM�G��4�v���+��1�N�}��k���g�Уm������'�g|P��F���RG��󾶳 � �4hY�^t��1���)`Y
��jb�H�-4+]���`�^V��-�3Z�����zv��l�vcj�(,y����v)����6��^�CsMYg���6�M;&�x|�/���ڲ��:ǸP�|���R�SHJ�T�6���7���kq��y73�RUX(ydAv����#v#i�q�jB��A��Zlqe�����<��T�A
_�>��짗�8���: }����l+��3��-��"�>�V��W[~�6��HNӮ+gL�u�N�x;��I]]�T?�c��)R������-���Nd�蛳7qx"=���|�Bq�F;��< ��{�8FzI��82�9C�9�;�j	�)�~7�Y�g��\p@%��\��Sɪyx��c�l�?���A�3U���k慮B��}:�l-�9�L�j9�3:,��O�7��;��	���z6fh�i-�%���}��~B��\M��Y]��^
��G��>k��
�9�R��3x�	&�[p���3������u�r��S��~�o����M�п%�ͼvJ7Y}������;�i�3�`�.{]��bN�מ�ծ1Re����������m�x�2A��D+�d�ض�������#T=é�d=3��KA�,6�C����&ǲ��N[B�=��V��m��}�J���Q��.� _r>�.��U�M�kw�|xk�Y�lM;�xǶ��p��M9LxRڷ̸*9���yc�����.:�0!٢D���S�����{Ǉ-g�(U�Ԏk��B�	����ր�l�.n�g��������/�! ݚ��������Ѳ43�	�+VJj�\�@��w�"U���&��Z�	ʺ|/���Nr<n�#cb'�,�՗4 u�͢�}O��~Rֳ�����8����B��x�N��sNCf���5�Ο\hI u<w+N���$�o�9�!��������M���-:�h0�"B1
�Z�%^��"��a$�AP�/���L�<�8 �7$�3��m|�����\T��9eiiѤ!�n�pJ岁�,��nP����-?u'<�Vj]�2F	K�P�a�F坭�\��Q]�3���yD>��G�sٞj����"��_Rj��GrfOi_�s͕�{���*��n�,U>&a���+;���;��r�_����0��c�s'�
n�[N�>�9�sOq��L���<*�#���^���C��)�ۉ�-�-��sq��^�\]��S?�(�h�������e�7����DZ��%���S��"a��2�
q��Bx�-�p.�@�5�8��7iͥ ����y$Sz� ��j��;J�`��g�3�G���F�� ?~�N�.E�Re H�UM��jJl���6�-$k�+S���J�қ!���5߈���~0��� "l���^(��pUjFb�.)�YV�"�]�lo������[>�*�� �K�s��_8�&�T�W��*�����B���E�����Ze����Ke��D�ǢG`��.�G[��1�_�3����"A���@z~��8K�yf��r��*O�v��B]��w��B��\B��"�s+.�����a���5m��S���!�2<,��;�F=�l*�쐹��}��i���+�p|.y��X��"Bo0v��ɚ�o����5����Cr�gs�{��w��Fo� ��ߘ -�ܾ	���5���8f:����~	H�p������t\� v`��gyK��])�ÿ� ��V�o�������S�ݔ���uCs�vZ�ZT�3����<���^~wo[�#�`��(�*ĭ(�Y�?ś���v����-����z���NnEA-��^1��;Yd磶K��w,��ӔS�,L�3=�G��E��'7f�B�+��%I����$:T�w{UkT�UB�b��Xv���iY�D&��Q��[n�	��-^X��=j*�(�#�%���l����{�E��2��>���T�3",��l�Ն��E��+�K����%���	a$�Ne�x�yd	�B�8?>;Ϩ�V�Œ:]B��Y�j��-��e��J-!�l�ʮ�,�!e+cp�늴��,�����眢�y*�3�U��ڇ0��%��� �JS�	o��s��l?���KM�'Q�H�s���rs�&$�ϼ�,gա�y]K���%�g���Q�t�)�G���G��ΧR�X�#�����>�3����p����dy$Fk���/��iV	�I�#[l�A:�KM�:EM3��i���
���~�Cʝ\퓯?���
=5\���Y��6�/��X�φ���z�M����褲.?>*[MF�x�d���#�T���5N�˥��0��"@':z���@6)�������l���]�Ok2�j�"8�_
1��?�)�7�{�Xl�R��"�#��?�]��Z��sn�c�/S
�؏$f+k�Pm<������25�tKϘmM#��
�p(�<��Hm_{�c�3UAl,a������WȫYNZ!$[$�0,dQ���,����N;A�9����\p��"���d�r�֖�<�}�;�Fp�dT�H���$Mɻ	�JʂZGr�9b�lC+�]͵kbE�U B�9i���Ql�����@��������H�[���9��.B����d�4��.��f�P�R>樾eg� r�"+����P�ќ�mՑ~����'�[}��C5MGwX����z]�sݦ������F7m ��J�t������,��)�\���Z��5���{E8�m��3�'�aC����'�7~�Q�j�?-����J�t>���c��ny���J{���B�߯�\s�ظ�x�-B���q�`��Fyt�*��U�2�_γ+�di��m�&L�M$Z �U6K5k�_|Y_��O�1�G?r�ht�_]l2-�6KxBWSH�߻J�Z̰MB��uB؃���u}��`b�VzAT������!�&�?b��ſMo��Ȗ��U6G��x.XA�r&�ME/&� ���4y�� �Ά�هLɽ���Bt��^g1N�n��Ŋ��-�طb����L��Ê��u_���6�kˑS�Ger�����z�迃��VAy���yE���Tgj���4 MSI�u���~.�"ܦf���g�~?H��U3�1�h��eƺ��JV<���k�|T%��7����T��������]C�}/�T�Ϭ��I6�����u�P���>͂GҸ��o;�aۑw��kN����rn3b������l�p*sK-D\������ү��E�'��}���UBu�5�.$O"Gx�L�'[��2Zyp�/+fDE�UxO/d-2�?�~�� �fC
��c'>��+�p�G|g�^`5���i�pp��o�ɲ"i���%�|��|Q¨�ԝ��	�O�ȅN@�d��@�L�nfP��y8�<X�$r�����N������A�?O�a�W�W_�� �LY��C&H��{�ev��L��r�7z���"K�M��6G��2��xB�3�ʩ�q��_˛�۬\Xfdx�p��-~�ѿjڛ��TH�>&a�[�.��{VI���O�~I���[�Ƒv��$�l0�������D,�]�����_��j��+RT�	Z×����\K��nY�$o{t�,�!Z�Iz�S: WGKYN��ݻ���>̉�(i�l��h�����}o���*�B~��}n�{�ڨ�ϩc�l����]�[ww�սaˣ���X���j�K"�g�5�O�������B�L�e7C��J�V�n8�V�Xe&�+�n�ZTN%��t��-�����ӑ�o� ��;��A�خ�%';��w"��b�Ԗ��"���pUvC��_��u�V��Q6����<��w�e�\�x�O8`��}��w�$C}<و�Pw�@���[�ʌ;�c��w��2�W�L��2`��z��g��������!�1iJ~��i7�\a�:M�r"�w=L@�)Q�~���#KF����+:V��0*��жǛ�`(Ϫ8 [fS�O��q+zF,�[���x�������Ri���S]9���˭��I枉w�jP���x�Xx�B���;ѩ�>p@���}��i�+�e�`m1�]� �ʊpl�>�2.�E��Z%e�c=��6�Qo�N�E/�1��w}�gO�A�.i�
��G�g܋ !�ϓ���E�p�k�h"�o�h��c����ܗ辳�6�h#�NX���,1�7 �\��rM���r0�v}uKb݊�˲�j�����P
c�[昉@]y4>�#廊ĎA��(=����DR4����=	�Z��jd��N��.Y|���������p�p���X'���מ�q�(�,��ojͿ�K,�=��*���h���b'j��I0�	�q#W��эN; Y�&6�H5t5�J�Fnoda �ᆙ�Mnvs*�+U��|���v����O�@�)J�]��m4��.���O7�D��!9�|?!o��D�k&3Ax�ͼ-ܬ c���t~p��4�v�/�2�H�D"��u�;R��0╁y.�{��%:w6��͟��V��K]饀dq��N�O�4S�l,t�_�����b�:`+oH�Z� ������da04�@}%�m��'�!�\�h�y{3�avF��<%x�2�ΐ#fl��`�ku�)���=���s��Zm�[�8�>��{~A<A��t�"aZD�[��$4���n�+Æl�Dh3�s��3���r��b
f5+�_Z�����.���r3�;Y�s�����h�T'���������X��[�o�фU�Z��p
�!X����e>�;�P	��a�hq8C�3~lTZ&1�
��'Jхf������$!ko��`:M6�7��Q�~�~Rd��-�n�0�yvd�V�ɔ��x�qhyV���z[?6&�z����'���W���34u,���m>G�Y4[�����	�W.3���u�E]�U��K��u&����Mx�l��u��b?>�H�)����hS�0����ayA�����M�7mJiU�d�
Q.*�k�������o���9u����Z�M�9Xlav��u&(r�<���rW��u��L,~ѿ~;80�PN���X�&�G%���_4).Q�&.}�K���� "�t�ݰ�j!�o�]�B�z9����`Ѡ��.IQ$.\Z�*�re�e`B�}���5)hzJ?�YS��)�۵ws��I�l�/��������o�P�!D�_��:�O	���W
i�Y�
���j�0�l�N�H�tC|Q���8'�7�l��0��x�jv��w(a(�Ȟ�����G����gvm1"���8t@%���O+@-���cǙk�t��FC�d{����u���>	��_1��ZCG֓�ˇ��bĭ���L� ��u��x*�ݛ_��޵J�4�p�0ߋ�BZ��e,�=S� À:qx#T�K�&����y�<�K�F����|}3��=�-��q����.�46Ӥ4b���V��W��ؼ�� "��Qϝ^ev�	������=J��`"{���a4�F�)��2���yBK+��I���g��_Y�#�v��	���䖋�];�k=���3���{ރYb��ī��y��{�}-c����7�50��jU5pZ��F@��G�!��\� �����Ek�"N�uT�VE� \��=�Bp4��c��))�;)6U@\u���\���"��UQQ5S5���([�փ|��O4�Ȥ-o�1�;����5*�'�W
 �C������X3ʏ�.w0�(������ ,0:��$���^���(��W��[UGq.�M~Z�_�;v\�OE�Y2�mg5/��M-��\1дZ�s�
�_�f+�3���Q	1v��'*�q ��QU�0�ͮEn �&9 f�Ci��y��Nw�4<o_����8�w�3XWl����g�{=��>=�(N�(䢻�P�K%Q;F?���Ѣg�uaɋ���\ȵ�2a_��m���):�VN;='	�u�J������	o�N{<l������[sq0�z�X��Y�eD�@h��x��fF�T�u��C/)F������������h� ����3�?�>�����]f����@�·��"H����ŗ
�?������zev��K�ޅ~��ѝ�	֚+`��~��v�����=��i���k8
^�%���C�р�4�����U����v�զ�����5H�z��1Gذ��wv�	6�B����g����\c5N��o�%V�r�C�\�S�5alT�5�\��=�_t(S:}�F��t_$�����*cJ��&��hyprP��v�!j��9,s��%�j�O��k�C��ǖn�b�W�76�����R�����q�\h�I��q4�-/�8f������^���:��REY�� 9��8�?ڢ#�yc�m�%|n��'��z�#as���R�aյ��Et��B�զ�~��{�!�_�A��%��4���is�)�}ChM�K�]����hH���0��yɼV-kN���+�������1\�X��9��\���a�ʑ:��ѨS�+�]�Y@G�^���ꝕ��d�,z���_�<BS�m-#�c��/�.�$I��M�
��;�d��Y��%��7�a�qH"_�����,!�h���G�7)�:ב�n���2w����ڍc�;0(�iG_�A�o��+nB���ny��t��yaw4e�
�Ku����e���P��B��d��IyJ�ٙ�U�/���9�l�c�����(ѕ�34���F��E�O��퇒2~��`���y��8E�����?`��t�9�ڽݬ�?#��U�q�P0�&-�j�
d�lYW?_����v�p�7�ڗ�.t�Zj��z�|*�iߍR Q��KV �~�;�h�v�c��B���� Y�R<�x�q��졤�4bqu���;%��$(kU׵�2�l]��Dowmh[V�����%��ѮS��*oQ��b�#m�f��g��gی7�j:lw���H�z�e�.��pHW��ne���!�1�ɯ#>f�e���
=u��yנ������c�R5�'p>\O������)x��._@��X4���ب��f�UuNK�b�p4�*2Ǘ0t��� ����_�ބ耈��N}�b8����؃���&b\����Y��b0�c����|�MJ������ ��R��)Ӯ=z�)��d�P�gktm�7N���HT;[W�*0��! Lf0�d^%7Kcd��>�lb���	7��ȇ��￠!��_7�ᢸ�V�еwy����Ά[^Zo��Hy�_���P���_�]�w�p,��&��3�'�2��;I�2����t��O��Q�s��a&'���c�c���3h'W^�3]�e�")ג81��B�*��)����gϞ�At�^��P
�^_�d���O�dǄf�
�D�¬��Q%���m�1`�pF��a�Nԁ���K����Ţ�	���ch�}�v����ۛ��Y���jA�>�C3Z�/�ϳ�3(כv7�gr�z���J��ZlUN�ݸ?�����	S��>Y�S)�k�P%��q���ڴ�*�9��g�[��Á͖!9��yR��O=N�H�У얞�X),+ �r%��.5�g~u ϮJ!�&Gl��2H�Vem[��|h̿�#��LL�e�����/�e��7��P^БY����xZN>XPֹ��P��MwN��D=�\aEV�o52���XӔvJЮ�d��:��r+��(AE(��o������՟���/3���)���в4u�$��2�FSØr/<� Q�mk�#�a'� H�y�q��$@���v:&ە4�{t:��H��p�°�9c5��0�W�Ƙ���ni���L �y�L���Ň��5y�ANl52�w�g��̿���ٜM����{w�ݍ߁�#*t=`�I���X��s����?�v'��}�K��&[1OeiQB��1/-�"|�疩���|���"�[A�˘�7["��̒E&0�'��K��%�����V��~u�ػ�t�*;A���(UP��wr���9=1��.����%֏�Wx[a.���7@��2".�-��n��cp:zL�Q��grK�A�r]�j'�'�>V���LL'��<Vj��tI���f�$��팩�͈�K0D�|�{[�"�A�BZ�2��--6����^�>�N���\Mh���,w[_%�l�56=jY2�,��83�������;����2z�qhM�FrrJL�\�~Da���S=��h�!����N��e"5\:�I�~���AB������hѰYbS�o�	*R�wF;��԰\w�5���筵�@�;���_�V�7�)�ٮ@�j��}��j�d�ɭ���z��3�A��q����M�]�I��ʹ��H�O�3,�.���b�~���i�O�����F��l�=<A��w����)��RA.9O=�n���k9v�H��@*����
eTT�<��R� *�S�W��(ϑ�,/����7$!�5�^�d�{[��1�ߩ���+b� ��,��d��FR��՚��`����^�$��x�+�<��f͞~v�N�c�U���z��%�(����e\����J����g�����4���������+�@�6�TQ�U�U���2YT�Bʰ �f�$Q��­$JZ)�m���Ͱ�'S������Mu�a�k�w���^�f�I��,�0d`��u�f�n188�ک�%�!��D4D��&{|�2���s ĸ�k���^����ٍ=h
t���J�Vg�ѷ�8�$����?|�
tyZ�q݃�}��i���g���ė�=�焤ڿQW��A�c�C�j�u�ej���!�v�X,;���b�V�Ol�1���P��tN��m�0i��q���f��z��$K���+��@��{�/��v��/&���;�5��1���ȼE&���f�c�R<אR�z��B����)_*�e���<�8r)4��e���T\��SU���Vu��FԬ�-��$�ʏ3!fe�w����#�r'��9};��~eP��q��A}�U���^bf_�i�q)p�m�Kj���R66F�s��]2M�$��~.�K� s�=)�ָG.='z��;���5���By�QPa�xG��rU˦�����$�@h$�:{飘*h$�X�&:���c��S�uq=���n<��G���6�Geb��]��ϲ���\�I�a����|��$@����v��:r#i���$<�\X{�er
���*9������kʗ�Kȑ���u�2v�"ݺ�w�}X�8s�x��c��A�D~b3e
#���u15����,\
.h/ { 1��}\
��9Y$�#�����s�q\"ĔV���w<w��C	OX�X�B�n+d���I>e�lӴ���V=UV��yj�"�Ӎ�=6E�Y�t`����^'e�QU�3a��n�wh%>�)�/F�:���wWt�N"8_���É�s���M�'p�y(KeZ�UԺ��v�;� �]�me��/G�ϓ�Ҍ<?��dofI���שׁ"��F��Q�CP�=t�a��QA>��4Ϊ+b�'�SrQ�Z�{����8��$-���� � ����~T7C��?jQl۷Y�'�"��s��w_ww��T�������|+���mdt�C%�c<�<V���@��1�E�ݩ����Z�+'9�j���2o�c�E��b3��j#��He8�<�{LO�w�D�y��N��������SS.H#���H�z��ܫ��~pN���k����L��}��*<�_��",��S?�$p\���d�P�ψD�쇋��-�0��Qk���'�	�y�E���F�m��hrn������a<\:ܕ���f2c�BL�����x�����k����E���ُ{J�44HjA�l�������)$�{�L��zI�:" Pތ� �V�D2�c���PG7�ȃ/�^2/i}7B�G"bedVJ4)8���μ��c�W�C���/cY�p�h��N�����"��.���l�sM<Χ�[�O�_S6����&�"=� k�����fĄ��v��vꙁ��`���9�{��(�"�D����pv��WS���Vl��0���72������2�|z��zC�2���i�mj4��w�MQ_Y
��S�L�B)j��:U�,w�J4�^�8�(W-ǳ%���&�=?�Bl�<k�m
8>����N�E��7.�{h?c{��;���z�����T��IJ9�䜖%ZZ�(���k�3^�y"����T�Ǫ�R��j�6x�;�;�nc��c^w<�J�."1Y���f�k���w��+=̽:�T�FZØ9m5> Q�����%OƵ	��� ����]�s��ʽ��FK��aݎ�p�K�ي)C��,0�~������i�5d%��!��~ aR�����4�;=�''������1�1�n�6��N3��])�e�� �R�P�Cz �Q`��t��8]2�s855��j-��}�%
S�Sh�Nń��򂳐�FQ����Z�&���pq�'�� R�	�q�f`�)�8n�}�iT�>JQ�I��{c�����q���t�-UH� |R���xڅ}���K�k?�_��Ņ_'�*vu���1��#���O�_�5�'(��P� �:�_�<�w !�ݷ�9#˒RR)5䳴�#X�DD浇XYP1̢��	#+�L4[z����4�?�r��[GA|Q�ʵ^��؊iR��	[��ڵu�NbW�U̾�Q�ҷ�����6��ӑ54�|$��fnV���fy���ٔ�X��(h�`S�؂5iOJ��K��^��J�8�J���i����`�,��׸���-%�G��f��A�-(�, ����S�z�/	��Z�跊8���#FzY��_	TB����+�����MS�����3�o6�:W 3�,3�k�3���e��5�e�8v/�qe��C��٭�gg8�NN��X�yJ�iE�[e�;�1�}0�4	LG��K!���y���l�K�U�Lo��<�\�/��w��jxX7'64���~���>Y܂W`qQ�	W{{�FO����:�c�q��h�uq�d+�(����CMq�b MPi�3[���Ac�}naa{s�,���<@�P�h�C�5�f�����7[\
L�3�)���I�S�A�:�����b�ڟ=�~�~��F�e�D~%�G�\{~�׶��a�����ҤD$Z8Z"D�5�k��wæ�H�{��*$�z `ꀘ�o���a��i�K��:j7IF��2��Ȣ<|��J�d�}�)W��I�,�r��J(i��go�mȬxA����ZP�')�^�1�xX�$n&kHG��F�A��ͪ���|��vh��F���MZ[[��zX<ɜ۸���z�ƐE����H��2��~��ev�Z�}�!��D�g�z	AxF7"h�-e~N��,�f�������Q{FE��$����ڕ$6Hui��|~��{�O��gZ�UQ�`JtյI7�'Ԙg���'�"�5L�����'�(7c�	H�=���N�3�K{tR�:M�t�k�5H�R2�o�[�g2>����Oj	�Z]ڙ�����p�;�ȗoxe��H�w�� |8*HwL|a�4�J4�m��Fcw���)bɳj�e}���Y���Z{��i-����ĩ��)R�<��E��5��J�w�_�	��!�ٹ�M�r�����t]��2C��K����;��]v��L	��3����2?7�<���[u��eC�?��g���#}:6�I7=<��o�/dtkpl���fgGz޵-�ۄ\v�0�Z�z���k�`zr�l&}����>�Xa�ޛ�����exG��Ԅ��j�"�15S��<$?��86�/��a� �y�|$ϓQ�4��=5�M=_�cځ`0�q�5���)�J}nE�^�ۢ�������6aD��K���N���k������X���TK���=�D/<�����:*�:h;ߵ��@O��y;�H� K�h��@n���Og�C6K���~l$�������I�ۺSAD�^�$%���VceY�#&�V����M^/P�`n}��_��-��T6*w��`=4�
.# ���^D��W�{yUΐ��\ۑ���1�����A42�8?�O7{�vZ8*�*b�,�U���62��T�7�[Ht���Ĭ��ĚN>�O︢[a�Xy՜J��@ܕ��	J(���o��݌�����J��)|���^'���}5KA���S���SNVU.��ܷ9��	7��8bMq�T�K��Sm�!�����J��\�k��F�o ��+sK����	�c^��\�P����ȇ4�����{�F���:�c_Ęv|-Ս��Uḁg;<�K��$b4{>kPX���~�].~Ј���#�r; �~[�Kd7�<�Z�8�$�.|�Kldp�GOQ@㊓�!��+��}���+��S�����B�=\���Q�e�C~��K�W.�
˄��i��c��FVny����S:�V�(o~s��^7���|�U�0I%�#�����z������p[.UG��GJ�&�����rį�	~F7��׽�Z\lJ��Y��6�]?���a�S��OŢ͝��X3
:9*\�k}s0���O�E��W��{�H�V����
B��o���[<*+pS�^���y��67[��@��:o�3�X��Y��B6Q���l�
�D;���x3�@Z{�����$5�w�+o�M�&����9�=�������;��