��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|/K�^!�� �Ϊ�I.F3�h�]D���� �1x�ϓ�k�K]b�ec���9�̑�2�۰�}EW��E�aǧ�b��S��+�/Aė �d��׫�~^^��y�4�4pjTK��~<OS[�EI|�ݾ�wi���tW3|��.�O�	��t�q��Tj�����E�u>�ET�Uj�a:W0�{E9�0#v��g��_e�I���7���eW�t�Z�.1`��u'�8�7p�b��I)�XO���n0����߲����7ɬpÝV�%�T�g@ ��bٺ#@���&պm/X�b��XU�PаgEn��8(�4kT���(F)C�)�@�ޑ�Um-���T�56Xj�}�ڴm�nCO�8���t7ྋ�ߧրkǎ~hc�U�.sТ���?��yk�0���)��I!��I�>��Ўru����}���T�-?�"����$$��%B��/��@� ���}y�ܞ0h㷴�<|����G�֢9���n<��|��X�?k(��x#�b&��ӽ^�,ܴ���X��jNȺx]�^r��`sNC�GVl	x<9L�_4���أ!���m�So#�r��vK|W�S�a��Ѿ�U��<����=�V ��m�r1��&�4n�>{�6���!���֎ϑ$�1pQ�I�'�<��>�N�R?E�U�e�.�\��n
���SI�q5�;���3�?�n��Fh�[*�3�`�pՔ�Ya�e~Ù?1�&�8��; �+��v���zXǡS&�p�wK��.v+E��F�-�g;^@7낄cqif��s��p,�'��L8K�^%Tp~$+4���f�����7��(�� �|6?V�I��w�n�/~�ې���׿I���z�y���h� Su�AШ�ݴ���ٔ�鑇)���K}M"oS'{iV�|�ŭ �i'T��O�͠h���c��#:�!�~>���+��RR�����g�<�A��?�P´3&��T�Oai����ND�Kv6����
f1b��m���01�ٻ&�6��'݈.B`
�q<<��Q�$i�������z���Z�K?v��?6����}�1�K�&�xj���z��-��Kn��ˤ	ڢD=z�xIc9}-�wG#��?�3�|z]��To&!��n�����6�/�{��ކ*� �m@܋��J�$����N���%g#��18ƹ����"N���~���l������Evd�!�g®���WL��H�R�`+`Tc��@�l�۵2�cSE^C8����-�UD�z�|M��3�m�6,` -h`�Q|Ȫ���B*��B2�4���8�šN;܉����C��rHMA��ZZԞN�#��{gZ�;�	S�/�� ����p�q�W@d��"-|���K�"x4w���������T�TM^�*��=�wSǯ/P�I6g?[{��n�ף?&{����ϱS�暣<�a;����M���;����F����X�i�0FMr{ZX�r���,�հ7ͨ�J��mRH+X�2�ۻ*"_I�d1�3,]�{-��u�D$=�ub50�;��(Ӊ��12��ZU�Jf��ɻ��L��0�HR� *�c�F܆R��Z��^�>]��z7�"g@�VPsDV,@��C���]EF�ݓR�e�����m���)�֦n!�W�\V����78� LL�0�����i)3�謼y�*i^�����^�hl<:�L)�����(P�j���`�q3�i���I�[�G��J@��R����$m�S���@{b��)R���C�܊ -7�)1�F�w�HG�A]�_�T�)��6�T�w�B���Z����<DSWf_*���t�ֵ�8����ɩnÇ#Kɘi����އF���O�(=F�bǚ�)���>�X$vBO�|�3�J.��nM��U�z�r�<����'�J@b��Y��by���!ԧA�F}�+mz3���F���S�7|!��
m�b/�~�C���b�ᡅ@%g�O�Q�b�]c�1�u;��uHNً�!z���8��c`=?��w37��'��r:5?�.!�!�;~������0HTs������k��-��="J�
қ]��((;�������T`5,���x�Kx��r'8,��+X�������	��TV�H��|-��Mi�=����,7,Խ��d�5�i�MO��H���ɣ���nG/ �*z��n��[��e1����OT���DL� ~�������g�*�*܏�����	��'����K�����+� ��h��L#67�A�޿���2��/",�YhQz�q^��E��Ʉ 2���FY��2����Y�[�H�r��ֲ������\8ĵ�;u���nT��&��f.��9K��0���}b�ї��MُkFN�hdmB�4e���Τ|+ndH��a�޳��MX�Qt6Ή&�1ZX��Y{H��Y0��҆=�ߤhh;�-o?�x�J��&��FǢ�f���e��z���mx{-:��>_�H�-��7�O�U�<`���8�dt�%d,�2�4`cH�?��>ē�p=a%��L�C������]�d�x���GtV\��x�����7iTrkBm�I���ef!d���rqF�����Bj����R�/�ɡ� <�#����>�E*y�H��-~��:�+=�<[�ٹ�&��TH~�y���%���f�n�;��������l��}�k��ą�L��]�$ �^a`j�nG�=���UN.�~��ܥ�D�,
�iD�	m����\�=���q���ܑQ�ԑIe�_N/6�Ҋ�8�[H�yl�먆ߣ�0��(p���ca��004�4��v����������꡻^U�EO(������\p*���#�������n�����-~&�w!����K��� ������U#�9�YU ����Z�f!��GPf{�tg&OH8�����(�3��Ιv�*��>��T��el9wv����Öa��^��,Mǀ�a�?G��DX��ɷ�;���^���FwT�����5�Ĺuo�G����5O���?(�E�1i׹��4��&������P�3QR����������U*J~��l�T˫��� �IÀ&Y'�p��d=<鐶���\�{�\�G0�w;�Y���&�U:���ߑ��/+��
�<��J8V� A죀MEK�����eQqe�'܀)k�)�+�=H&#�(l�*nm��X�)��uv�C��B{M�E�F���{�LRz��a4��L�����Ē6�� C�c�j��<�:,#�A�/��$@W~0"y�:�-��Y��������r	��n���$���� Q����F�2�no|��R9�V�n4��Ue�u�R�Ϫ���ӭԿ ��������cP-�|nnl�k��2оC���$E;��4YMȤ(�R�����b�*��og?aR$RD���/k��\������l<�g��L���]bnI��Al�K;"���O����?Z\�Z�1����e$�y6�-�����'�bݍ�&�B��K��Os�=�3^7s�w���6� `��U�-�0����ة�A�y�abX�c(xs(�\�nR���+�������I���`��h�`�N]tK+��wY� =6�\ͭ\mfsL����te��A�wM�ܭf6�;ny@�H�}��uY!���Z�Y�0�pɼ\n��p�2�l��@�ӯ�y���z�n>DW9_�%�:U)[jm69eN@ߐ%>qز:��p �ڱ ���&��_���k�]v�[U;��A���L��Y�9(Y��h����8]f6��@�R�H���0ť���&͵���sNP�,�P3�/�WPHQ�.b��p3�$��WB��u�.쉣���b�^�-h�q�t��,�s��R��
��"��o�dPo(V�7ڰ#9da�]�9�Q����Z|;|�>g�g*�@Ǥ
�����v<�nQF]��,٪-��D�M���j�U��G�j�<��b��h�1���!U^6S2>�����q�-;�&��R�~�+`����Ƞ?�(��ʩ�\��ۅq}wE5�k��J��>d�{����T�q�4����3>^s�T���P�U�xW���8��
�{×�/����|9�+��|��qX�W��Z�z�0ʉ��eW��\X���|9a����]r���	M�(\�X�nB�gE(���̭z��B
�!�Yp?��e��NH?�&q|��l8s�
��, �o�*�F�W�z�˾n"9�ک�����c�-�@�]�yC�/O<Ý���8��ޞ�G��v"��-�A$�(b��K,�q�F�6��2�[�|��վE.�$Z�0�)`G�V�v����:��S ��5r��m�߶G���gM��ő��{@��z ݦ�Ru�7�:�_�����l�j��;� #�f_(�KW�C�5�SӾ��3�I���J������d�ݫ�xbx��qݑ|7k6}g��5=����Qc�H�'������d�����@l#*�"�c=�=���֤w�mH��>�ή��K>��f`�(2~5m9�&�ݥ��f�$���{���L�UMO��eo�2�Gn�FE��o��sd�
k�j����[�!Y��$�p�E��^��V2�Ss޽ܷ�K|�I +{%T�6�&��&!��fq����I��'�o��j��W(�z^3��ĬD��ډbW.�Sv�I�뜳�QJ!��;�1�u���!+4�au+�⠻��%�	@#�F�~��'ؙX�Z�0�f�������g7�F|n�V��W1��%Ξ�ȬrP�+���N����Fb{��G?�Ъ=�M�
<�ĻT��9��ۈA��UW��qUc�7�vR��\e%�!�H;�p�dNg��=g���k���Oc�c��*	YQ���I��!���:b�h��?��U0��G��r�X��Tsh�/�d�k�g�F%����S�ay�C/�������aDJ�&�kM�<i� ��fҬo\�d]h�%A�J�I�G���Id��1�����PT6I���
��§��[D���_��s��X!8�A�����<��OƆH�z{�#�����'.�S�,��0�0*��g8J�*�	�		��YRc琋Ѐߣ�x�ؒP�9�{N%�T4���'�B�r |�����s��?j�
��I���m@V��:�~��1M��4��kl7Q\\� ���>�WZ4xM�u�S%~M71�uH_P��7�x��"�}>����d�*���f+�>&���i����.�sU��^b \�'9<F��ŦI���%�*f�CKI����mR�J.�?�A��(�6���_K�ƣ,�Q-
���9�H��SV��v�-F�lc�d\TJ���q_ӟG�ݖbPܛ�\��'he�e:~�'[&�4'��|抮91���(#{�$E�F�_��j��=��n(2z˾$���8���ޕ�4!<BϒCR����+{5��gI��3��|Sx<��_c�t��l����^|��H��2@Mf�}�%��8����(�?��{i_I�~Г�F�{���l��IY��9�*���L�\�ϭ��Ş����/�n�^��_7H����ϛ���J����2/p�=�Nm�l���=CĤxbf�O����� �~���=��=��[��(������t�0�`�~7�CT0,G��U#�y9	l[�v���鬯u�):�F^}�qC�x˖����
����kP�(Ё��1�`-�I���X ���K�M���`v���Ru�4|��σ.�q�רƘ*�y���e��N,�� ��ׄ����ч��u�ōr���Z�)I��E'p��ϞL��bLPc"$cB ��hؠ���T��2�]tjiζ���>�@ߔ�̲z	,��.z&#��M)����E��Xi����(�;?�Kg�4��*^����h�Ȫ�:���k���cd�o�ϲ��_�r�@g�<��i�f����J[��U�D]P��˫:�2���hx�a���F�#�^6 �ߵ��gn���	^�P.�)�~'m\���xޞ�i�G���>A���~o`Gr?���&~x���QS'���d���,�9!��~ifu�%�to2�v�JOC~��4OC{-8�.�	S��V����S��Y/�Y�]�x�*���j�mfC/f{HhfC�כQhL%ly��Y��g#h�׊�帚g���s�����>���w;V]E��Eg���+�YMQ�A�����ibM��R��Xή��i9nT��EJ�c���X�</%f�1$��1R��(p��4a�`
�?ה�*:�7��1!���E�Y1(�g��[����a�^�X"���+ I0���4��l�H������7�д�v��V;V�ˡg�_05vJ��-��������O� �V�,��X���G<�)��	 �����p7~,�ylk��~��=m��i̘�{�ժ �.�'�mU�zi�wb��S����ʟ��^��T��*�t�"j�PR�E�v۾�$�-�3��s�3'�k�B(N�a�O�W4���JJ�x��j�[�&*��߯�su`�j���i��B��A�k����x �S��'��3d;�{,����\M���Yfa��7��u�Z5���l�|7�q �}�����s��nM�MS��8`��u��d�`�����Z���U4����>���۝�.��+@E�E �����&vk
�ں��X�=�r���t|���0`:�B7����%��y��jC�u�C.A�$���2�x�`x=��c�7�7 ������m��N���!g�N�����k�3���?LKaw��?�e����	�^@̺��vyƌn��V�@��Kq����6���$h�bެ�XÜ,/�� %*:9��Ԕ6�_���*���z���x�@�Q���SVb��,^��o�*t����c�/yő&�Oj��FÄ�YY�V������fIm!�oK]�|m��r0)�� H��o\Rń��أ�j:���X��1.����iak:sZl�16���8l!j�����G��a1Y�?Q��%A��N8aȯ�x�v�Sv��bv���_�@k�_�bn��+���)Ne�I�=? ���D6p�NB5ۮg����2�j@�(�s�	n���=#�]�p�5��
ǚj]�[g�Ր5���։��R�,��+�kv��(V)=��y7��SY��;�E_�^I�)�C��T�y��N-�W�Wb�+�}߯5��ު��L@(C`��U/�v�i���s�����P�ڽ�[��p��1_Jwkm���iUF�c�F.=�Si�`2�y!�~�쟥d��򍏨�5m7 ���F�� Zr��)u_���/s�`Ъ��6�I���46�zV�11