��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�8k�)9�k���J�f ۘEN�R��>�Ug:�&�1��ꤛ�R��i��&᤹�e��G�!�3g�}8���;{��DÄ]�\/6�6��Z(�P<�k����⟇Ԑ)��i����������Q���o�(�����	�/9�B��*N޼�l"ͫ^:�J�Aܞ��aH5�^*,L%��x���	��臶u�p]ؖR�P�z�	����%W����D?L��M<�@AѢM&��RH�� Տj�}��4y���t��}��bm]��#�������튠j����?%q;��A�^� �r���C\�ÀR����A��'��kƞ^���lޭ��I�ۡ<<!�tޔ:��sd�:�h�h6�}j�r%�O��vu��	@1'� 9$_�;���o�C ��j��Z��&�|�ǿ^ x�ڝ��������Zy��r'隆���c���<���Y���ʆagį���̎UQ�����v�����љ�^���L3�����s�MF���o�\��j�h���]�G�Gf��Uky�4��I�8����J��N��9�kd�ew�"����rN��|�cư��𔥮��hC�W��sn�Ę�S��DU��Fx���ݵ���x�x�T�����D� ��{��WUo�L5ԪwI?N#16Tv���Lᬈ5��	�?�L�x��v�%YA!�a��o�r�F:����7��g��"s(���e�=Z�f��c�Jv�o��p��|9�������+����;�,p�9�(1�˅.����Y�����*��;�I\e]7ֆ�|����f{���we�h��n>�A�2~>��Ѩo��r��ZV%��5F'@�3�'���n8p�aB}��~b�g�I��g(B>����C��#����i��ݔ���.`.��ґ>]�-��f��R���mY�!�nJl��	��p��w�xZ/G� ��T;�����w(�0�9:Ș�Jwg��|�,�/B��fOj���D�@ԯ|1�9�qT�7����w��u�-�>��S?;���{mн����-��l�b��t$	�2"�1,���D���l:)�At���$�u�g����g���yi�|��q�i3��|d���@���;_����[�$f	8P4��v�}H����;5!�J6�Q�A���CW3�F��uL���"��x��ퟒ{m�EB�>[al�*�B]��Aox�v�B+K����b�G
�F�Y/�P�~��Zf�X6Mp��Oͧb�u�c[ɽIh��D�@k�+k�	�n(���{���M1Ja0�y�+,��Nl���k��L�����G�x�>%�!v�u��\�٣�
ߊ\mں�� ��K�K�dJ2K�܋m�+�3��G�_��y����|j��_5���F��	���N
���%�i�.�^j�$
eXUy���I����%��p�RG_7��� ���O�s����˩����,�� W�B�q�`wHOX�����``@C��ݴMzߪw@?�,&�����|kht�%���]"!,r� �-:f7�bT�EN�/P�x���)F��3��F|��,���3���2�ţq �����:�*�az�n�a)}���"J�O��մ��ϛX��di����8���_��u_4���������%m`��M3Eay�������%ND��3� ���z(yEl�en�����Ϛ�B3bDyÍ4��f ��4�G�� q����T���H�+B�<+��{K�^6�\�,�w���!� �I�/���ƪ~
��P�H6�U �34�?Oǀ�㿌�`Ī�:����7�<��D�y����*��'��a&�1�-�`I���&��)��$R)(v�eb�:K�`:^="�$��E�_q�-Ѷp!���B��c�%Ù������	�g���"�!"�<��~���(�����:mX���O����2T҅��u��d�]b.:����_dd�H��KT��|���������
�����M\��C	mW@��)��E�/ך;���K���o�Si�GչƗ�!�M&Nl�v�-=c�T�Y7�n<1�,
!��iTr�
��˜]�+Q�bYm	�j�R9�ǋtu8aڹ�������REc���^�U�߂�t����9:.7��4�$��m�n��3���FTH��:p3z��VxI�5����\��5;��E���	�
3f?��!�2.����)�j�B��q����b�y��g����������䯪}�<�-C	��u���S�j�+_&tz]� Pbኆ��l<aT��M����B�VC��p�#�y��G�T�W��_��_�'��e��CH����V���BG�
o�(��qh��$Qh�,b�w�9��x!:l�=���H�!���2-EN��Fc[��?P�
lg��5G���F8���M�`U�`+
�C�R��ݬ������a��1���y	h�K(�ړ+hD鵜�؛��r��e7���4ǛB[�r���6TM�0�������L1����.n%a�~uܔ���8��e�i�.���B0����l��������Ҽ� H�ԬX�ŁW�*�޷��R���`���@�*��<��Ūw����:úHq/�v/d�����9	l������1Xgc���B�i)hM�a0d�� f{R?�`Q${ �љ7{��ZJv���욺&��!��#�b�x�����#s�t��A�9�Eԗ�u��㫮��0;�2���WO�@�%L�WJ�^�rH�$�ԍ����Z��(�����S��0�Ul>�h���g57�52�}2��s�v��L�B��f Z�Kex���N�D5Cq���v?��<��l�B[��?`����A�����k'�C+S��͔Al;u��-��+���B��>���u�ܙ���5��d���������z���Y7�#q��1��A�µ�W�����kd�-�Я�C�8j�B�Pٝ��.nV�+�X�4�̒=���]ȁ&�8���������Q$:x_[��};�����G��4����{ِa<B�1�����9�֤{�8����l2�B]mN�U`+K�b1�@�R*?��4W.?�'����)J�=vu��B��Q`v��^������m6j��w��ؠ!���nq��sLT�*~U�+o�uޡ�1���̗�Z@`&�y����׀u7�$E
b�[� JNp: /By���� �*{�����}t�\���5|Q9��V���"�G�t��CVxѺ��R�M��l�'k){�V���������@�@��������0���R��%����HR�G�b������{5�5��[C��IDW],$ ^��L�wvBZk����6�O>��#��~�"������RZ�N�.l�_F��6fY�r�>�.�f�[Q�E�@?:[�jKf����)��ީ;�&J*�h����ʽ����鬃�\������b��\3����,�|�sʋ<��+'){��+���3�.�XXg&8;�|�O�{�&�L�t���G�?��0z�٨��@�f+��ڰc���;!��ʎ?�|_�����+�����s}�����Bf �&���FOܕu^5!od�\D����pw�i�����1"-���|=i�~�a�-d�.��v MZV�nIW���[�S���n���M �/XR��0�`�lB�#���7�{��8tD��Ѹ
V��+��%�b���̤��ٹ�:o�.uJ}%�b�1q���y�qbGG�}��I{��"�����j�4HE���ir�������'@S!s+{��[������@g�$�Bݮ&�2 ����n$��r�F��zOyz�^fTܷ�F�Nܺ� 	�@v�Ӯ���Hrx7��X���An�Q_ϥ�g=����q�B��2�9��H��XwPT.Y�e������ne��ξxѭ�L���x`VF����\�(3���Yρ(�ԝ�$�����h�'�:�Ԧ�rDX磲����\�0�����ǫ�xT@�����On
�L�7�US��D��K�y]�{���zv.����>�������4�sgg%O�*�M���]��|vl[�=7�]M�[��޸K.�rقc�?�	�󸀴����&��T���qD�6y~i��Z�����G�}��Q�3һUg���x�ؤQQ�j��j�<j�K��S���@,�U���GPT5	n���	�>^�6�9�vٍ���y���T�E���$oR��Suk��dU?�v�v���i`�~�C�0����X@��;�۔?;$M+4"�TX�y���)�H��[�6���qˈ�Z��N&��l+�c�G|�9�e��潅wp�.�*L��T�%C�K���	�t� �G�|��a��U��%�:�#r���Z�C�������Y�q�1<�0ڇPT�!����e7���f�H���������5׵�(�������;��L��t.\�L�B]��/�I��8��:y���47�Q����[>�!���"#A`�	ؼ��Na-qq���ށ!�J����8;ʤ��Lp<���(�:��H��N/YJ��w�C�]2t�nd�Zg�!W�vlYy�ކa4�b�$=��(��@D����t D�(_̧$��T���A�����ɺ��b�9H�'>�?y�xC*r�p�G&���ӈ�=�Y�u{Vi'`�����$4ߠ�M��Y'Z�	bF;���v%=-�)U5�M(��SI����&���%�޾S��m�6�i��܅](��6mb0�����;��E���H�M:��믨|Y��]��r��$V\�a���KyqՕ��j�QA���KݼE	�Q�����-ќec`H��@V|?�ï���� Ё�ż�E�	��Z��sG��X6S�.�-��K0�S�*���{�Y�B����f��� �h��--��hV����J5q���%�� U^I] ��`�%����G��Y"@xڛ���;�|S�[�l�K_Yp�P�s~�%&�&��c��󍆳��3vg � LG?z�@�UX�:g+jO��x�x(V]&(+k������&�PqJ�u9�p�{���jzR��/���2bm[J��Q�R^ZP�:��)�`ۏ
��aC���[�$��T���.fanN�a�.���
h�����B��Q��R��t�kE�՟���ȮaC �k�o�c)���q�f������r�����U�|�(�KoC0:[�L��ռ�5��Uu�O��IvR;�c3(Op`��?��>�֥v+$�}�[��d2 (j�"�9�������/M��V��m"Rٖ�����	P��'8�������3bE��
'��8!F�w��y[�����x�N�CJ99$��)��N���Uc�1H5Qa�g�6�rW�?�Ot�G�z�ߝF@eC�_K}���mA���OO���L��9a_%0%C�c�{�l���Ͻ�i�ޱ�~0%Y��W�κJ1���������6a�f��`�
ӮP�'��f�L�0?q~e�%�q6���0q�B+��S�'�lG3�¯��<�
��P���������1���T�;� m���BBԱ�{)�~�h0��p��8�^�&�� �z)%�*���c�JU�,�1����6����Pbd�Q�hͨ����6�2^�$���BRl%v*z-�U*`�7ꇲ�y����p�(�߰�t+ЈP#/
M�0LA Z�1�<Q���+B�]�ܙ��>����W�b���-2o��(�q]Gw����)#d���u6[�Nm+Aw�_] G����B�U���瞍��AP�B)Zx�~Lw���<= 9y��\��Vn:E����@��!��ٲc]�v���#��7���$����)	��@��N~?�O���e$����Unؐ�гoG�.��(lL�� ˎU����t�0�6�n�gz�q��t�#x����UR��s��Ȣ�.�UOX,A�gT=��2Mc���T����M��[�dÙrf�ɧ�^�_ե-����>Z����Q"�U<PZ;�7��u�[nA����+�������Z�(9�*�W�c,	�Z�q��� �!��Q����bo��R	�P7��u�?��Ȏ;��`��!Kh-ED��F��dn��^�:D�)���7��梧��'F�9�=��}�c�'�h�	��\+l� GԮs��(ϼB5������S��e��OP�7Ojh>��^w��� M�y_/��������[��������S��X�u�GP	6v����wJw��xn�E���`�L(Υ �@�GhI�{��땀!A�w{7���U�#A;ձ�K��?/Ú$D3-�v8�!|=��rw�j]�򁆩7��GM��oّ8M�v�L�u��%��gx���.A��@{��<1d��1Qw����K�;���J�I�� �:�a�h�crth�K�� �D�����"��Yɴ��@����_sIu19�>*ܯbq\�M#Y����"�9R����r��øh�8�|�Jxӡ2���韘J$��ER�#�~Ѱ>4n/�Ty�����R����Xmq Oa�����dD)�8L�vW����@��Z��$*a]��'G�9Y5��W�������5����k%�	�&���9��Y���2w7��K�p5#YΫ4 Ićc��:l�Kx�m'��F�����|1c%�O���{ۃ~�^c �]�s�u�W�r@�D�񴲬�������lQ�tX�迯�gj(�@�U��v���"�%h}¿j��&�,?x�K������li|�[w`�9����j��0�b��l������|)I6��RXl� t��N���e��(�?�>i6u8a^ �u�|�:h.[�@+OJz�%�ࣿ�����C'JI���\*ɸ��q���6�O~	1h	����lZ�L��X��D��_�c��%������Q��[���N���3����Ѹ�a�s�"��h�1Bj�~JO/u�����i\SK��x?�K���)����[Q.T�ӛ{98�fD[�MN
�������-�'�9�,B���郄~K�7��n���ڵ&�I��,A�X��������$�6Ի`V��u	��i}�P���n�4�ɮ|:��ֵ���F�X�(U��p�Gg�E:{���Ԙ��:���`���1�ұX��f�L����3:DW���g����	V��{sp秼����t��H�î��	��]��X��eN��o4�`�Um2K�ˬ˷�� &G�)Uxsō�0@�R������,e��St۵$;�}=>`�*8.d����o8������=2�ߏ���߉}'-��X �'�1�C,cA�W�W�8�c@��4	��� �!���K�&ڔa�)�X�9j⻬1�sh<b����������'q�.liθ܏7H�r3�X�6�=�����l;���VA��§A}�f-��윒�{�z�O"s�����V#i$�).9c�j�
sZ+�J�N�P�u�ċH'��,�D�K�j���餞N��?��΀3����#��T��Z��_55>Op��9�$M�%h�SB�P6X��~�P+�,��&в���`�~-g�y�o�Nf�R��F6:���ʈ�<̒D�g
��5�*��R�kkz�&:��ab�p��~b�`כO����a_=��M���]\MT�Xj)s>:%ޅ,�k@
�@$x�湮e�[9��,\�}ę���*J��Q�V+�a�N�/I�Ҷ���	�X�H��U�vE�ML!�i�^�����.�},M$Q�{�b�F9���|�TN3#ق�s��q�S..���I,�O��R�&ʹ���@���@,185�d,~����:�ߕ񨊩��Id~���?��C���r�Ü�����f�Y��;Z�)�����72my��U� �i���G�Q4��݊��n���^5'k�p�-�`�-Q�����qMq�K��������\�q�{�^�,�1�=?5�B�+���ay1�B4U3�
�+$�6��u�UV�:Ä�̫�6]��
s�Vb�m��U Q+�=Bz�Nw�4�p��}���ɾA�ɋ�V�`���7Ԟpڵ��)��U�S�w�\�0iQ�����%ʁCi�o$�ޱ5��)d}|:^1�8`+d6��O�1���(A���@��a��:�0R3���`�Έ�wŽ9��"�����X�@�l���*`�u&�:Ћ�Y��'��  W~�Srt��i��qy�X<���跜l��������3?���r��C+�:VRހ�h�C��cꮑ�J1LQ�!R�IxZ�5�#ד5=:�x���-�G�v����Z-v-���~�9o��=�y�8M۪�"É�1�/�&l�0���X8u�Brl���,�����E��fa@W39R8�O����>�J���%��Aq��r�@���cJ�)F�)LW�}̐Q��4n>������# ���N���~��0�����Z���"��Yv�A`�>Zչ�P��0��S��ƪ�!2���`�uO@�B����S'}W0�?�j�⮅/�Q7�����Wg-Z	�,*2��o�.���nq��ג�dG4Rn�M�$Y����sT�Zk۬X<PC�G��f���Z�����3���EYκ"�5ċw�6-��F��W�GOw�x��.�1b��mfc���SR����
['i?��������Fz�U�Q*сX.��-�t2�X��6�u�b�!b�;E� =����!8|u��N"��4�O�G
���o�p{�w�2*�Z�d+��A6��"�~é�D�p�n���&���9H���x?�IsY��?6�^�d8��&E�tL��\�y��{����h[}YE9����c�V�4l�t�K�I��9�]p&���8;�bI�t��ִ�l���Ui0i�_�k�ʢ�Z�8C���=��b�����;7A�G�q�+i�4��TƉu�(�>�u���m���ypJR����'�9����L�]�@����ѹx����aE�q�R n��B�g
�M#�7�r6Yڇ*]]f�4�?� ��#:d��80�e�S`�O�����x���]2ė�%�n��B¢��Z�Ww�笓�QE�Lӷ×�u�3ֻo͇�5���S������t�o��l��1-P��{H��ߙ�����.&�����tH��,��χtso���,��3�yw#q� 5A��C��sņ��6b�t���d@��-4K�"l�3	�)z�^PR�P�[@ʎ��[f�l3C�{��FP?�����8Z��h�m�Z�oa�|R�-HE՜�#���R䋁{geHl����}�0�*M
�;��%0��U�"3�˩�g�!I��t��|b��Ma̼���9���LǦ�+\�x��)I�fÓnK�m�<Ԓn��b�V+�i�YK�'{8 Ʋ�.y��?�b��z#�nځ64s�q#i��X+:Oc0W�X�"M�����颂*(9Hsc���ɵ�fZ��=/|��I�Q|�Nas!�҂��Pl�l ���M�=��ފi�#�]��q�
���>��$���2��NiX��Ϭ0��E��Z�[���W�P��q��.�C��?�� U���{z���7�w��!���x!ṞPb��1�Z�UN�WCW��.�<3���Vuh��v��M�����,Sj�
���/�pu�*k��QN$���ΙH`�d7EI��*J����I��B��%�u@td�W�&��O1�;ֈ�B|
�c��=�U�I%�?�k�6`�T���jRh�\6(I�Ȁu�r=��	Q�r8����-�'ő���$j����T��P������z�,��!��x��T�n��B�2W����_}D��qA����y���EMH�~)$�p��bb`	u_�u�U7]�b)���`�*�X6v��A*	
�K��$7�8�����A;�K�	�Cɀ>�+�o���T$���u�0B����F�){�׳�*�S���q)���>Y�H���~>%�:���k�v�LCq�?��ӟ�����B?�������L�z��:1����Wl�@A�
괭O��^�8,G�4�BL��?b9�������#�Z߭ �m�Z2c�ϘԷ���tޔ���g� JҾ�v�Ll���b"�(��Ȳ����k~���-��?�Ϲd8��5j>�@��n\��������n\�v���g�=fR��u�r����G��Zmҧ�����d�|�DF������i����B�����X󰺄n:DA]�k�.��gy�}˩J7���ts�pf�L����B�*��.N1����:>kE�%����u�Yd�յ~�1Ēo+6�*�k��[��ϨЮb��,$9Hz5���h�*Cm7o( ���0�L.��f�����^�(cL�G5��7���Zߊs*^1��מh����fԲk2�4������l:��8�N.�0}IP���1������5"u�2�!��|�aL���^2��ݒ�͛���;�~�:��%�"q�}�h�� g����o��nC�9.�.�Z"�ۀ�.k�Q���v�)��7z�L�d�y>���o3���Rnt@��)�6n�ݻ{Ŕ?����E3-�\��\��Z¯��8���ho�'��~Ǝt�������Æ�~h�'F������u@i,,�9�������&*+cLsP���i�Y8�r{�B|��n���`e/:�_S��!�K���Zh+��q��R�D
ГKf�����G�D�Ug��2w*d���a�36�e�6�]�����'��U�J���{�{o���%�rÄ�����)}�ߛ�+�X� A�v��E�}`���8�/����	1�t�h�5���̟*�k���@1*�Ƴ�h�;�\�����9Kf�/�$�W�!�#�;߷��݉tT���f��/���*\H��AFc��S-����P�0�W�R�7���c5���{}�r�2���a`���Rz�8Z�3�QݛE�����/T�:���H<ŲBM���b���ۛ�dsj�q����S`��%���eM���pV\}:M�I�|�,�����&]����hb/��@��2�u@K'��L�jߜ���9@x��DI� I��w���]�/��d�f���0��?u[ĒG_�P��8�mQeTd\����eg��w��R@Aġ|�l��J�Gs���(����������dk��F��h��ow�#���{�E��� ��LI�aE�!�Qџ�M��R����NE�bn��omJ�^���+�f� ԅ�&�1�EM�y��9�������q��)���ut5Ҳ.[1�f�K�^�ho�G(d��~!���+I�[%���6��ȫ:�o��j��r2X��������6D��Jo@g�U��F�������4yH����Jll��P��	hx!b����y|��m @Z�v�uU5"HyZ�'���8�V�.Mήfڌ���bu��ic!K=�M���x�2F2|垒x7�8����;)<�7&܃�S5ؒO����O; P��Q�¼.���Tܳܑ�������VӜݦer��r8˲A�^�>Z�N��T�rs/q���a[��0�?[�^[k�:O���z�q�����䷩�k�}7�ӪD�˾8��`�XM�u#u�;�逩��k���w��G�ux#7ҫt]e�HOV���YL1+@J��*�1e(Z��Z��A����:myٷ�Jsm�K\���9�kt��2�����{=vRoOR�������_��!��@V��o���~�&b&�w������u�X�<���&�Uq5IO��+�f���s�@�YlK�,I�U(���A��65��-�
��{g���w���s����P���~����,�e�v�0qǌ���~�����#|YIDC.t��?Rx�+^��_�`wh�U����4�8�ԓ�L[1<�|����Adz���0 T"����-�o�h��H��� �.��mX��4���8�-ܢ� �f�d`�i��G��R�lH�.�tNu���@����5�߽��Ȝ�Q?mV��J�D+Uw/p(T-4�H�|ux���oe�lOb$N�WU�G>�i'�6���ԒT�)��Z"�u -���if�H�������N�7WFn.�y��C^�Քn�V�����$~�M^��<l�{畽Cp;M��o+��؝�++�urO���&����Ⴋ�s�H���V��@o���W|l�&{7'8�D߀!/Ѧ���0ժ*�G':oH�?4�[��fn�� ��R�?����Urڐ?���&c��ew� S޺��A�>��Y�U�|kĞ�X�S$b1���+Bw�����l_���<	j9y�v��Z5)�2�3Bj��Òm*-�C��vg�l�����wU;r\%h8S�Ԃ�jk����h�P}m�-�xd�Q�'�Y}��y��e�ƤZ�� �h@�N�lvw�3QX�����l0#{�� �'Tmzx`f�g�����V쮛'���Rm�+���y���Uk��+D�=��!�W�e�P4�{V�Ώ!�]�K `Sh�F0�`(���|�U�l�����/PWw��
�x��h�v|��;���FgH(��>��� _�y�B]t�Z��$�U@c)�3�'n�Ի)gH��>�G��1����ݝ��V���h���^k����7�߅v�%�B���4�h�t,{��j����6�!�pT��x��8s��Z�ΰ,�FF�A����!����� D���2:�=���� t\��U������|:������Tn�v�r�<,�u��Y����Dy�����gfb9����