��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<S��!O �&_d�
c��p9Om�D�ܱ: ��S��"Tx&@Say]�\���I&��R�WLd(y�Az����YDYi?ѱ4�ɻ4/��w����.��R�";=�Y����➡\�i1�C��޵�T7���D���q=?���/M��X�uգ?�XXnN_�b�S��k�Npo�Gt��m�,��,W��	��[�j"�3�g� �hI4T$����{j��{e4���m�Sq&�}���W��ԛ�r�N���w;V�К��,e��U�n�*v\�Pi�Ε��KēC�-K�k��ZE�BnJ�Y���[@��HJԽ��#����$��t�y4~�-�9��)EV�����>%gQxWW��`;n����ɏ�7K$�dA�G,�i"���.�jwC6�h
��E���vˎ����m��ՠ�%��Z6�%l��c��y*�C��@	g�c�d��-��FTЇ�c��*/��އ��@��PH��j�ͳ�ԋ�|�0�BN+p0���:��D�L=�i�j!t!F���<���"~..�킩M��Sv�\�&P�M1gr��b�Y��9l��(�s�a�T�*M�m#T�,rw4f�&;#�[��Z��1��{�ņ�f_U����}z���n��� |� ��C�Ȼ��@N ��%j��<!���F��dJ��OK�aD�U�;ߩ�rY>�QO�z�tw�Xc .B1�Ֆ�-��Q5
DY�W�c����	,�h��8E;��2�&�.�P�!x�����}I�[Zԩ��?d�ZdtEhÎ��s��S$�=���*��A��0Z�����"%"�P��ކOWQ��=gs.�8�y"��c
FL&.��$2�����v�A�����LmGi��
��/iHpSR�r�X�&q�Oq�,!̭�];�Jq>��z0%ݵK�x�te2�;l��6{2�jSz�����v% �G��:�zȲ~')t4��ɳ�%���'�;�ʌl�A_���W �ǜ>���Y,N���KSl����\��tSS�,k,/k��N��
����`0�s��H!l42��ػ!4���:�Q��P3wр�\y�J��h^���֜F~4��$ե��ؤ�K-�K���>!l�͈�͛�N��}<���r�{T'0Ė%�<�~��X��N���͓�Vv�/�u#��Q�Q��Ȕ��������6�5�7p����Aj�2Ϯ������y"���P�	�R�=�Z��1�J Y7��a�uP������4 $���^ȔWX��CRxL��]��#�R=�k{��#�_��`���yv���(��R��M�S���Q�2��7E�2P�J��ڈ78 d=���0��$�\6}�2Bۦݾ�	�7���Z�| �!�x�q��:a����-C4f�s���Q�?��؇�i�����T�����w��߫Y��G,���k%fzѫ��s��Q���r�1E����UÊ��=���F�f�3^����υ�=F�2���~���@<�d;|ѫ2;��U^�(�P ݻp<�OR&x�Iމ8-�z��$�V����DbH������{��x�%7���
�UP�22]@Y�sE.O�Ƅ�<t,$$b:���(;��:L4���0\�fx� �^.����\��s���7ls�{�Í̒�]���I��HWZm��M!gU
�
�2���	�2��$������pȠr(7�/�	%Xw5Sj��)uZ��X[䝍�m�#m��B_���4���G%x�P6� )hO֚膟F�CawA������ܙ�»�oC�m v!�8e��>jJ��hZ�N�M�-��7jQ��Kٛ_���%`�(�����+��<#@0��x��������'�K9���}�{�0��[Y_���cz�u�}4)C=@����8>a�e����"�&v���\� ���XMG���#t�xO]�?�g_Q]�j�|���cr�[:�M�gȁݚ��c�ӛ���X��y�."�OdJm��b���j��B3���ց��k[5s/��)���qۯ�28n�	��)T�[ۧ3�H���S��u��D������#h���%6�2�|����Q#����N�Hub����*4�� �f<��Mf��X�TUO���[;�R6�\�[��>��pA����ѕ����'��l5�)�ɿ��Kh܁xkc �02XP�
o`ل������6xv-�����dَ3y�F}b�z'<����*)���6T�,^��x6}�0��?��
������X.~�a�D���	[k@�Ml�O�8�c搇)�.H�i,P�&7AW7����*-\��*|j���E� �U�5����ct:�H�t�AՒ&��(,&���������	��[s$�S��잂(�S�鰬����x�����
���pW�H�$�I�m~��>��C*�|������=�Y�ٷ��ķ�q�D�!Tg��$�j�4�Ny�o��\Y�q�,s��A�k9y��Zg�}��fO�ڜ]��脋��.^;e�|�\`5��	�E�\�z�U�I%�Z��z>�<����ou��d�^���{x��M�iw���K�&��	K^~�$�j�S:��Q��yN�R&ή���k�b�E�R!��-�*L�w�}^�<O�ک+^��N뵍�C̏Ϧ�r�]��!����{�߷�5��ʿ%��m�]Z��F8�چӷ�$���6����C�0Lhm/�G����x�π�<�7ȏF�2��ԃ^�^q]`�EQj�C��s���U�'�x��R�N���5�n��, ��-�Գ��⏓�G�%���]bI�yTG c��l�_�����Q���U���8{������("=0	�3a���!�$���5���y��������5G���j�{h[$��Pk�A0��0R�}1���(^���� y�Եlm.�I�R���lsy�[�(s^F�a��=��N��X�D��t�q�G�q�Y��#��$J5G�aB�k���)�&��(e��Bei�͟��lBu1���g}�4�!���/���K��IM��z�x��y���j�b�ߟ�@<(؊,:���'ܷ��
|&Z��Y�RJ^��+Α�^��C�k~�tӽcK<�!k�;9�*����[v
�ݎe�$�����R^E�����ڎ[qRB����Ƀ�,л ��vPd�q�c;�:u:��2]�mtM|��7U�
i�e��k�`���t�����������^h�6��dktW1��^Y��Z���#ה�'����FѬ�cŨ(��'�|r�0цЍD,:`���qEC�^�����0�Nх+�G>̉Ha�Oji��+>��1#�����-7tt"S0�!��>����ӏ��3�C�ʅ�1���AB��Ƀ@��1��"qJ����g!���|��IP�BM+� n�71�O3���)���}a�Y���� ST%��-ۨ���ڪ"(�D�&Qx�4��UP�T�
��δ[ t#��	-s9�M��'5D�?�ܸ���":Ӓ%N��� �;�R��R %qH�c�j���*/��9�Ѣ���k�Y�"&b��\�.��d�XK�7��N��,�!�$�]�mG���1a�j�>C��J�rȻ�
����6�ڗP[�G���g,N��ĮD��آ�_e�*��W;a9~���b��\7%*r���՚��݌�8i��FB}��~u��@HPp�(k�� ҍ҄J"�o��~�( �{ـB;\R�s6]sA��Q��-0ԫ�s�ND�,�R.���0���Q�J"A<l�j�<��i�Ln�t���8H��ƺ��c�s.;��M�	~ӷ���|�tW��j�x�FDy#!SD��̛���I���ʊЩT����0�>C5�Z���Ֆ[OӤ��n(��y����C�H�P��
O�[��W��qa��T-�ޯ�a�q��'�&ޢ�Ґ�EUF�$e����vM�fĈQc{ ��]-�JL`��O"��;fj�lY����CjTV�!j�C�i��3��e���H��yp-�҅�d0�2�8J*]DR1��jk[`ݸ��C(��o�Q9�FN���ڪ5�TUO	_a�z�i�é6�,�_Q���aؿ�B������p�E�/H.�i�G�-�?!M5)��Ys]���& �8���us�_�b�V0��]5m!��Ğ����0��qdΎ���ϻ���B���������1���/�S�n��v�2�ڄT���K�G��\C�\I' o��L�YN�	�	�}�.1�Xuf�($Rcg)�y��3�E7�9�߃���������@�k���0�Z�3�B@(I�Z�����)��{������nӇ�a�(�.�8��t;;W1�8�[����Q� l[�N,���:e��p�eʖ�!�o:�S�xx��ժ���;��;��H�$4��&A���T͗�|ݞ���>��k��DHɾέ�Ι��K���}�\�\���W�q���)u�
L �Dl��z͍gq
�$��u�|y_.�u
_��r�<U�w����ƺY	_#���tnC���,bf���q�WG��N?Oj�mT �͎y�$�<.{۟|��/��-�Z�~��Ϻ��x
�Y�O[��ڶ�o����{���g�6�����p�	4�y�oϢ�L�n�j�5I�ѿP~]7ӻcvEKռNs���(�'/�]���o�A�v�����*ΐ�-��0�.V�����`��Oc�h���;������N���_B��J�'�Ě�(�@Lu���B���rW���Y���*��`<�sp��[�g���q�^y�b���W�T[6�@	i8�tpI�jٹek���\�t(7��/�֘��x�����?��Ͼ��J������ H��'̯���NG/����0"�EcgFX.���P�\�0`����lxf<�>>��ʥ�,3d�HT�Kp�An���cх)�!�qp���,��0��K6�Lo�5�� �T>y�)dn1�|�1�'�R�����E��|�L��Laqڣh���ߠl}W�F�J2��!����Q�w嬶���DLV؞��}���Wg�6F�i^'枲vD'r�O��oU�����~�ݰ��}��ja���g�W,9��ғ��u�J��d������
�Ȝr�t�K����7���6��4 {�y���驙)�|�	������N��I��ZPj%���N��c��'��t,{CS�]��K�^�ٛ�e��/�XUX���o�3�^
&���{�>[P������{/Dvk�����5Q���1�X����7r���D7�Ǣ�m�JN����'�z���e���6�OG]Nߍ%���߈[e���v�����n>QTz��7@��f&{Q��bT'�Ǆ�Ú���{��Z9��^S�Ƿ;��r&��=���S�����k�簳���*3=�.S�jo���ȉ��'�oa��o+;M��xL�k#��K�l��Uش�-��H��P`4b;�wf�C��C{<����Ҷ�=7O%=GBU�5u[�J��`�NoV�&��
Z�g�Tz6{���!b�7t�����C��5����ӄ�:=;_���mOS���7}n�WP�������/�
��rn�羋V ��V��6Y/`ܐ6���鉿5@�q0|����5��f4K�[I�&y�5M��\?���̓��Q?�+M �v?4;�q9X	[��74o.�:�>���V!f�HK�5z1͢��Q��R��U����/爹Q�c�5ⷅ��r���2X�+YE����5����T�R�`*O��І��Pn�}o���g�:uN̞���u��.����<?��fT���1��응Sg��;	�I���6��aԌ� ���:u��H� m��ZdI�e["��LM�c`�]Mݰ���nm���*�p5Uw�5"rF)�T�rr���@�ȗ�)��$��b!��-0�Kr�cL�~&����m�>�&��x�[�\�� ]�M�f���G�'��u� �g�����H}��C�b�E��?1���c�5e����q��6�:�Oys�gv���y��7��T���y��<��m���w~h�Ao䓇��xϛ8��U�����Q�{�+l7ǑZ19�����k����9ɰ�g=�)~����w���U3� Pv,H�o�dNv*�&-��1�h?K�ML[��Vm�6�8�om�h��P�w�3��^05�h�ͻ���佂�7*��Wjƒ+🇶�%iW9��~?���]ၽʤ��|Ъ��+�``���,),�#Ma�Ҍf��.�����/��-k�ڮ��鰽��p	I����o�8�(r�I ,�\)6��H�j\�`6S�6*ak�j�M��i��76�|�.�^��.<�ͨ�$���F�D6&����c+j��3x��
5�%;���u����gqǱ�G�����^�p��Y���aX�Pf][�\/e����@'&��.�a�	�O�}D˪�Ik������ Y���v���3�����>}{#"�}h�,���H�j�.R������ ���� p�g��a{gW	�)I�X=Z�������/�@�j"O���X���o�<�GEW�)]꩗�U�^�P���mT�Zf�ڮ�.��)(�!l�}Z�������56zזj��_���,���}�ǆJg�SNI� �3WSV�V�l<�p$��Tc;�����iD��>�^+�W�9���L���a��Pj�cx�-]���Y���:��`G�0����1��z��]�n��t�0�QeE���5�uX��hs`V�\R�ҧ��2Z�U�]��_���� ��z�~q�I�r$�m�3�G�v�v���~C�t��s 1�TI��!�O�x��~��j�����^$ߟs'?z{@�ݮ{��	��Q5R�d.��2�ej�.y��<�B���m���#Jq�U��okT�&'�5�uǆ�h��
�u��+H��=��̀��]K���	a��݈l3�-�Tz�\C�<�u�/�;�c�'�q	g����&�N8��f[W?�gG��A��)�K��2OX�%	�L-b��!��C{�2�8�r�����g��R���v ��!d��rs߱�iS��}�i��U`z|6�q^��6����о�9��*��9N�F�&?T�Ji��a�Y���e�����a�;��6~֚hLD��~���@�B	Xlg;_��i���H��){�X�-��Yi��n����H�-��
��|���~hW���m�|3�ԃ�n��$@wD|!آ����^N^Po�PUw<}YR�-�빗U@��*�蛞"�Q0o	�j�ܗ'�_!l�z�	"�S5�5�,��nڦw��ӕ�m\���2Bby�+�
E�r��0htT�޲=���ܵ���_��o�#�nޞ�5�j n@n�x�Bxnz҉r����16�Gi��F^C4}j?ORx�3���$w��3!@M?𹼙q� xI@U;-���a
�&�IğV���Uc����ɉ�&l��=6���A�y���I/���H��&&��ͻ/m�ǧ�?�Z���F�J���>�ä��?��`���۾���FM�w�vB�-��x(Y6|V2��ᴭ�y���̰��$�����9��:
�ߛ�'�˷�F�/��M4tz+��1��D$N�/��+Uv��ı�� ]ɖ��4,�.?6��>I�r�3�[bN\F�Jl�I�|���~��f���`��x̵�pTY�D��*�#�Ƀx� ��Ly�3�I0�W����9��`�z���毰��vP�P?������ D��y���,�	�1��u䝽U�S[�YBвG~8v������ݬ�oa	�I�/A��a\���n�1S�yDf���YtJ���s������ �B�ݣ�ľQT�*�2t�At���z��`!Qw52's�`��Ѐ9o������(��Z�.,[c>��j��ʰK�3��1���,v�9a���/�phAt>�=�����+@.�(����	�q�2��f�!��7��g��Ʉ6�3��b��ύ9��}��`S�� -����]Ǳ��?rs5�&���ڠ����x�7�~e�t��h�"�|�Q;�Cg�`�6��8���!�VB8r�A8���-�F�xG����5E2PT��
�v��$�ȇ�ˆz�@Os����RV�z�W32� ��W(�����D������~gIo���m�%H��[C�]��=-�TX���ҳ�*U���h`�`�����`?K(�)N���N�62�ė߬� Y�����cW�n����eX�4ئ�T���',�T��ț��&ȷ�� ���~e�?�fLYr�Q6a�E��\�&a�S��
�^=�1 a5���d�ݼ���vĭ
�铯��#��V�L���!�H�Ѩi=1dK��u`���/���!t��F�M����M�AD֕��8��ya�5���U�a;�*LR��^�K9�?l�}�8��/o�xsAQ���ޛ�Hg"��傤�-��9N?�ϳ+�w�Y��1"�(-
��B�S	��I����Ñ6����1� EP(2`JN<nk'��]IA�~����� ��L�57���u-�i\�M	�M��QWA�Cp�����=�RL��.�V��C�h�Hy��)�(�7��V�(�Ԧؿ�G9Ck�R�j�D�6A�4���~�<�Z"x���03���%囱�r��,�c���q#1~���mὌO��=樦�*�EBYBM��-F*%R��T6�f���!���]U�Dt�/��o]�9�+�rG)��5�m/	��uh���~���\�,j�汜����WMfџZS'2%W��h�����&��*	w�hC���Y�+�kmQ�$]�o�_��I��#������]�Xb*e��N���hU;j)m<l��N=F���k���<	�X�U���R���i��5��	�������������>�c�$#^l�fyo7�m��)p6��:�N!��&�R�c�&0�tC���b�y�~�s�h}2��A�;�3�#�O�\;�ŨH� ��H�L9HAr�;ΟH�m��'�D]ZDF0��6P�ʰ@~�r�ńp�bƏe���(H;ZC	���K�>!@/
^t,���:'p��d�
�`R�)����-������S��#�k�tf#t�2��
o�,���یM���}^Hn��0+Lb�j�Kߟ�_�h��Bv���*~���9wm�g��/E�p���c�h�Ⰱ%g�q��z4���Q������f"l@M�Dꞕn^2Su��/g'JK�ފ������(]���H�tl�a�p�&+��9��D�h������6�w+K�xhr˼D��-P3� xH�R��ɲ�i�&�#1�����ѫq H��2.4C��O�3���+���z����3�?���$�M.�́'�d��hZ���a��Ίvk����L�}��v�~�8�?�Q �+�*]��}���j�5���u�.J�,lf�JBB�VOJ!���#�6E��=��)R�/ذ��l��s�1z�)��<�X��Hθ�	�k�2u ��Ws����o��t��ܠ�g����EbI��0���+�z�`�o���<�˿��񀔰�K�ď/���b7w�0�T��MV"���.��p�K��ҽ��y�]�_S�nf�&�V������)��!wkՁ��ϼ���r�K�Q�p���'�8W'���h��'R=�u�"���ȁ+qr�1!���}�@�SWռ�DM�<E�OR��������u�q _�����������P (>�c���	��Z����y�jI�j�H�l�*C��j9oK
�����A�B�#����%��e,�+��.e�c�)��h8@��2mt��A���8��Ƙ+X��b������i��Xc�48H�.�����r�C"�uM�rN�X��de��Vг?{W8 6��G��l�`zEa�ro$0�����ZvBt��e�Q����X�b��g�l��	{i֥C�#;x���T4�􄂵�s�c�9�����+%�~�k-n;$]���2U�Nn�M��i舨��J�Rp�7J��L��t�5-vn�Į}X��z{oԏ�,ψ1���ж�ix��~f�,O��AK�ug|t�N2�&u���y	�j��uq������:�.���>��-j�E ���<?���"�v�@�v9�������t��Q��R
�"Xj���w���O���2ď~t,�����$�Z��z�m�4����������O(�u��B��-O/��#�+
W��NU+���r>�����tz�ck�Ư�4P��Ŀ<��/��"�a��r����*]?[}��_�?0��dֳ��ټ;K�(Q�g�K�̊�1
�+�e���^��Pㄺ���i���ď��ɶ�q�Wt�렀̸���fϤ�	>~L)���w�M����r7Y��nxN�Ev[��Y�H��KA���i���T�45OhD�_�)��R?֐vͼ����4@���A c����C��Rd�b� .)Rml���W�o�69�̝�%�_p�(��I	n���1k���얂����rh��eo���k��e�N�>A�^5wq=�p��R�D��Ni�^ =BQ)Q�W�k�I�/��Ƭ9��Q"��'�&�"$d�Mw��{n,&j�+݋�3<�Nm��U�O������&SJ��D5[	5�\�
8����4T��D��C]Ә�A̧=�VX���o�̸dj�*g���j��664-b`B:'E���Hӌ~FM �/����J^&�]��Q��ϲ	������Ă���f`x^�Z<(Ƃ�#�b�H<*�ñe��6�ǔ�ș.J�ۍ����cb���im����:��n�غ�q�u$G4a��V����Wd�ۊ��q\z�N�2�U���I)��@Z>�s|����"�5��°���r* 9�%e�K���}�h������\v�������N�_���i�����D�`�F
Ohd�PE����`=?�A����ܯN����5�Ǯx��va�q՘��+M��'L�H5�W6;�c�F7k����t�OZz���5�Jg��q #�|x[%A)��� !5q��E��t;���83o�H^�݌�tjR[nrш]}S��n������Xx�EY�X����H&�_Zw��L)Iz+s��Ť�&��}�X���&2�����ώf�$��P�顸;�� 8c�[�GX�u����OLg o2�D�,�0�*~��\0PH�)����n�O�� CKʗg<��BW���I�|f��S`pfuX2 ��m��=�,\�؟�F�h�䣏�y��i��l� ׃DI����Hۧ�y0
Cwp߈�hna�SJ!���:���l�+ �/�{�7��;6���E��hg{�zf$L�㴴R<=8�"Sݻ��59̙�zG��̉�^��x��xa���V�j�R�㴄PuL���a����I{��T��� qҚ|tI���V�/�d��-��}��6��J0�����z��{�B�G����.����e�[IL�3UIP5j��ф�X���,����iZ��byLt��}tD�(v�j�Bj�l���Rn&�r�P � ��:���"��cm���x�t��7^4��j|ĸaC*���_(>�`��K�b�Ϗ����E�K� ��i�\@j���ҸG���i�	�����T���bA����/1Ę"G%hxs�!��5��)V���fa C�:�,��0j����c�]�b����Q���T�,S�ȵ�s���3�:��+��n�1���n� �gi���;���g5��w���+���i��N�σ��dX@�z~+�K.�)�2]�m��_Uֿm�3����w��Sn��q�����Qz���jYi��1�fD�jN��\NIƔ��*#�B���}Z#�B]�C�Z�	��?2��]��TQQc΃�&�$��x�n��w���������t5m��s{&��@�)=.�[y�����4��Ob]�lԧ�!�δ{�$�T��*�~./!-/eH.�X
0�����s$��u��PI��F��4X?���y�����C�{m~�4�*��l|蕜6ENQ6����A];+c���
�~��Bi�H:��G8��^�����"*��f�f�Ǉ�� r���uCk��V��n�DL;bVAu�v��tT|x^�S�r?�R�F�������A�g�ez���8܊L�ː=e�F�2ۜ�D�(RVf������\1%
�
7H1B�J�蹱�|��]-,�3QI���u4&��j]
w�>��U��h�~����l���x[�����M5�4�L=oQ]�� �H��b�����T�%+u���^���ۣq*�����X��V�*��^7(�6��	$�nG��H?��|X/��ĽRt�v��_,����P��|v|�^��ޔ�Ac�RW�N��Op'�t8�QM� 2d����ϒ���&�ʫ��v$|�A��ڵ����3�V&Ĵ�ǭW�����B��v�k����*�n���f���H�"��+��}Zw�/�o�i��~�_�Ǚ�%�g�i��m�`xF8���8���f���N:C��zG���\e��Kx�ᮠf�$w6�o@A��~}��=>�LrL�߶6���*r�=�+��I�U\�TI�owpN��׻���Llq`VQ8 ���I0 LU�.�s�f��d�
&�)�&�e�d����+�1�ԏ���)��q�4�FdB_b�>Ħ%/�K��âIRz��lh>���2=�#,��p�{B/A�1��3���Ic��:k`���Y�Z4��O���1�~�l�uNd�:@�,����^���2O�|�Z�B�H�A������W�)��B��#�E�[�h�+N9E�N߂��_%f�i@�+������;!qv�o��H�|�C"ʨ��.}����  mx+��{�E�ߕ���1�Ht�=ldK��8����2�������P��x�ǧ�AM����b�Cz`�hM��tkay`��r���+�A��4�����c��f��������E�M#.E��f�zW�����l�a��z�z�yg)ZʘtZ�5˰\�-mI�]vD�Q�>�����~} �9�b����$*�Z���Z��i)ԇ�J��5����!��	?�O��N	jA�	�'�����'"�fMd1i��smE��R1���fsU��B2��S�g��Y�Y,3��1�U>c�p�<M;,CѼ�@7�,�-3V�)��
�)v�,U���$�)}��E�^$G�p�ng� �F+_�3C=gO�ç,��YT�Ȕ�Y�~��l#����"���^���*A�~���o�R)���ʖ�־P�[��X������ȩXشĝ�O�G�������Q��B����*	�!��))k�ه���
u���PtI%3⪚�n~���=��Ԁ��]д�&&���a=<�9[�y�fU5����9���s� i@d�j�	3���	6�^��2��'��Z�/a+�ݜ��?�y��K���]�u���7ܴ�5f~�6��+���C�Ptv���:Uj�g�au��أ�(w��j�E�~�{�+uW�D{��'Y)����IF"'pT�gw�I��e��jv���U�R����ħ�;g�N��|U�������H�I���5���!lA��k��F*?2�:c�6�^��mY��sf�6��{�:�C~i��~�(kRH������q���R����T\˭	�-����]4/�^!aYDdC\�h�L"�G�l�&�Iz���-.�V��rvi���?�#�3/-r���ܻ?��ُ��������Q{{:�ȃ��Ȋ�����<Q�A4� ʐVd������]�Zp��=�_}���mV����es{T��sh���~LU5��!�Q�|��E��3$3�˱����7<i�XQ��l��2��1��&V#����VZ�?�b�P|�.��_x�A)
�r��s�u@>bĒAt'�I�eb�%pԪME,U�۸��]E�8^U4>��G@������6��3�O�@�F/��&�v����a�Q��Ɇ	F�sa��,Q�/ۣP�h�O�7H�&T��E���kv��FeP��y�»c�̀J�'xU�S�����p��d:��&�ֶ䡈�I��9@r�b){sT�x�}��LG����A�s�� ��X��7�]�DkB�����n��ۄh��C,Q�ur�!S� ��5 ��ۄ8:oUȅ�[@]�P��1˨��?��)�t� ?\�]p� 1A#�F���yQzy�݇#+hcٶr^C?x�|�9%m���kto�Xq��"\M1�Uz��5��u�Y2�a�.�����ۼ�����mg[�x=V�e�N��SkڈT���dR2��>T��: =A��-� K�`�4�l�U��lJ�`��/_�:�}��4��`]R���"b�7, MJG��!�d�ם�V��U�T$�����>0�v�@�7G3���u�FW�t
��.��[�_M�u*S�͆��F��'���{��u����M։�R �l�Z2/=���X��Vz�ݾQk�W�`s�����,f�8J�J2c��x �����&��s���7�X�@������N�L���a�ƛ���J�g��� �|�ݮL_���K�A�����g�.��HJ�S��J��>v\ݗ��F]��>�]F�pfܙ�<����K�0�q�!pd|�>�E��a��|nц$�f�o��G� I�a��P�H���+q0F#@��}��gY�e���z�0���X�Y��*i��n����J���Gm�TUrd�H��쒵�K߾
�@��l��ۥ�4gH�
�ofb}��~��ӊ1D�5h4 �*4�J֖n�}���E0�4rN`Ar+�:O��<�1
Zku��n�5��c!�@i�O4[j����R�����6&"�~�D����K#ؾ�I��)����=��X,5{�|��Q��c���f��qe�4q�Y�"V7��d�A���Cٵ���4�?���,�9�����:c_��̽��l_���VP@8�u�MV�v_��E����������׀�c�;}d�'��Z�$������v��]��VM� ��C4@{��s�ԞQyQA���{"/����g����ʇ�2�JN��-j�B��3^�jJ�k&�p�ً-]���TjJ�]��\��pc΅�q�	��`&sAF�ˀ8��g��Z6�΄-��}<�W����"GݵHM8HR��iG�	{���n���P�ǰ�t�M�)��3�
�+����˯�8ʊH�z�wǷTi�~�Je�������ɱ���%;������*�b�A�~��8��ɕT<�<g%z����ツ���"�����l�dD��afD��8U���{H3ʘ
���neQ�������,t9��U٣��x=��SϏgW,JW�ӤL�.1�����J^ZW�f�u�4*	U��|y�LL�'q-�o�-6n�@�n�Y3+<��d�����|��e"�ZQ��U�l�`��87�a�mR�ERAn���=g%�.Ѿ^I ꠫�(k2�����mIظ��5��'ďq�n�%��g�굜��o�Lo38v�z���ݜ2s�)+P��&S�Wѕ�����<�$͞���;��Y�X$���NԬ����`��(�2��j;����l��W�Ky�ȇ���I�v��P�1nt�1,�NG��G��`�<��:x����	C Ma[d�>Ţ|B�����JN}�
�S��$������������r��Q%$�5���S
��}���7FAꎚ�O4����}���&�ᐰ6��i"��B��,b�ВV�P���K��[G���Pq��Q�� ��O�ίD`�T�$�[-sk�[��|�`C�*�������f���C*�f6���.�c< '����S�U�|v�PHsQ��i�b���h���3�Q7O�q�X]�)����Y��/����������h(�h/
��DʫJW��l�-4�W�	��#£����n�,�vt#��������m��
[C�)�A[����2��.1��q> E{ yͩp��ю�����P�&�q���!֌C�FR���y�q�Xa���E���^5Y'UC'����������>�q��2�?}��s9xw)
�kUJ��/sU���q�y=L�%t���6l�g=�[�	Q��Z�ް�I��n3<�ӀD
�)�g�O}��bĭ���)��Z
���+�_!��������D�f$�$J\<���#��u�$�<�ۡ��
��1�n�����5-���1a�M�'��CRا3�ǚ!��.�I{ V }ny4����%����N�0�Y�EZ����[����J�T;�4��]�O���=w��ZWLU�4�J�=�&�'�6�Ј`ز���I���G�R0�w 6%�A�3'��9\(4T��:4}d�:V�B-\�vq��X0���MU����y��ś�.�8�z���z}�Z�֙��;�A��Hȃ����,D0Ԛ�j�&���}~�U�ܜ��@CQ�ϛp��&s�t����b��y�!��<9� +l�H�#�;����"���.��"(�+:n��I�Xd�Sw���=�(F�NVi]{ݲ	���Wm�L�͌�i�lI�����Dp��'�zo?�eҭ.�$�]��jg���D���x��]�I�ӿ`�U�+�cM@c9�J�;2"O��5y��)Ug�~��Q��ܳ���K��:�����.6�4�n4��Lᩆ��O�@�]���#��T����p�i&�5�&4�N�W����*a}%���kJ�Fr���s$���s����(|���|�����JQcZ�7�yl��H�f��'��0�� ���fjG�b�$���pxtH�r���kp�E���"Xw�O�3����8e1K�>�NC�P5��93�V�gn܉֜�ӔqOT�X�̕��fL�|��d��_�,�~q)K��Ep�m��A�����?�j��>�.�iG�m���=/��w��ˁ�9*�s#rl��.+]���qb�Á8~���|(ӂ?'�ϵ/ۧ���]m$8�̶2�}#�vH��S=p����g��\�ʇ|W�
�W+P�Jz�TS�ME�i��R�{�#�<Oж�Cם!��H#v�}ص��lz�?,�$`q��Q^���B�_� u�t����� �{7M��j�.Oc���?�)/�I�yy��b�*��O$���yP&efS+�R��\�礸�wjҢ����P�w�H�����o��&Ƒ8���
T�����\�M�V���s�8IDy����
��R�=�O:;�O ���):��IVE T�^U��w��˯���-J���6��� T��t:DDZ�2���(ha7�� I���ݪ]�T�V�������.
jRw`��3��Bn���mlګ�@�fh�T#�Í�r�����Ay&;���>�D&�{�����(�&PԄt��`��dKvIrt�J!�6���
��ׯe<�0�BP��o9��b��AqyHH͗�M��FKz ���
�z���y~y�]��09by�����6���k����g���#Ob(^p���;x`q�pϥQ-��k��ȖĨuه��:�Wx����բ��[q����J��R�6?C���M�/֛�n�Q����5RH
���hm��4!����}��3�h~��it��lM#���pn2r�Xu���u��ͮ�ky�`�;7���j��E��	��3�y8��b�ܪy��S`�(`�r"W��ф����W�Ԗ1�׳kF6ۖ�ֈ�KdU�}N��p޲�PL��/�Kk�*�Jj�˰��Cd6����u��������)h!.`�+�����wQA&��D��a���w��wR��'���K���`Z.hGݾ`n����'�>�f(��_��7�8=��)C;9_$+esԩ�j��M�D��4PNϸ����ܔEu��b�y��\��ή�|������[O�YcR�����$��F��{V�`�E�v�iU�\WvŸ�Q�.�g��r���7�����}�:�+�Z��?�W�wݘQu���]=�p��2�!���1�a5̗�2J���QNAٷGَ���CxQ��2�/Q�3].�=�:~C������B���8�D�ݏ@J�4��uq$������B]����2��Ӓ�^끮��3��hp���m�������U�/�������H� b��2��wX�O�c8[�<�/]�@�;����� �	�eD��}ɇ'����"WMn>�������������CL� ��"�p�f$[�� F58��R���!xKy@+&rA?Ǽ��wi��/�V�~vѽ��A�-���@z���n��|nO�$��ΪZ�k��N����2���zu>"���]H�?�W&c���	�F.PvM���Aƞ=�>ֺO0	���>(�������״)ܬ]�k��}�		�u��������J��8P���Y�m��`�P|���I��C]���жܔ.�x(M���y��F��5G(!+@f�`l��|�s���Rz��(��C�v�ԧ�s�H���sB��Y6ՍKu��'1�؞�ݬ�<��zj'{��N��]ۖk1�q�2߹�lpcǤ�~i[�V���,���V'ܹٟ�߿� �e�.�w��@�����x���.j�D�|����45���p���G�?8�񘲍��
����Q���։	 �a���@��uFR0xC z9be2��|g�X|A���`~����9��8�;�e׽Nfj�I��`��~f��TÙ�i�J.6Kr��L��<j?S+RG�)gR\"��/���w�b>�)���6��aT)ѣ0a��L@ꀀFU>����8ܼ)�e]=��eu�E5�g�G�k�J,]̛���.c���j�3d��zzrԫ��=6�l�<��"4}���+s�.5:�R�Ϩ�g���DB0>���j��_������̖�%i�������R5X�btK9�/��^��"]��B���������G�LI�eF� �U��}�[GH�K��	�2�t�>�?p��Iu�A�6��6���
p�8@
����W{	�羐���aR���;1U�{���v}��ءfb�wM�܍É��%E��.��NU6�4Z��u���*h�*n��Xoh6��F��E��E�৷%zK޺GTR��4�l��ϻ2c�����7B���?HP�H�Hw�Ͷ��ф$�Ai5�Q���y]Q�M��*C֑��ٌ� N��S�����r�%u'n��l0JУd.g�̓S��9�6N�$9�hU�B�"M���B%W ������U�q-/&%Ui�H4�Y3O������#��O��ir��RC�9���x%UHk'��V��#X�6�]�i6w���	U��[O���L�Z{�U�B�ڀ�j�-�kZ��0]�љq�_���?\� �a����e��X<������q���ȧ)N�� ���z��Ŀkκ�X�^Ũ�7��ДE:�޲�yN���}�́,�| rx��_��G�!�5lPj���a�����ْ�����i}���˻l^�m��vu���6�j+-�U��|)"f�e��*�/ɛ�Bښܳ�6DYġQ��M�jt�Z-�P����Md55��G�ݿ3D3��U���8���A�m��i�5�b�54�vr���=��	��>08xQ2ƾ�p�nM�]�QI�B��E������� ���m��2�nl�F���nyy����<�y���r9։�g��`*Wa��@]�,O�D�#���!Q}�YMC9Ti�'Z~}���vU��GL)����#���2���t����mq|gu��������MO�uS�U���[��u$����/�n\���^�Q�7�Z;~�����q^*J�\���3��:�6�D�T�U	��p�b���/o��jo��#J���l�~sd#��1П �ȅֹ�4�h��RR����n�N�ѹ�OK�77" ��R�#�֑�_Ws�)V=�餓.�k�uţ�_���Y�O Q�u�\-�l�u]Y�ઙ�V��6�U5�*Nr�� �9��؊�}Ȼ��S��}E��G�@��y#��ޝ�{0l�龜r^���Jo��Jj�9C��d��LD�d��=v�U���G�r�/X�mY����k�Qc�:lS+lI|,�M���<����M��U#9C����4���l�4ѽ.7h�=G��iI`�̗v��K�i�	 ��,n􏾴�d=>F��4����M��=4a>DCl�;��>��cf�T���1����D���1�2T{��1I��TsN��ܦ�b��6�,%��O}�	{R��+��YA�n8��/�V�R<O��$Hi.���}JFr�vF��&�}V�h�7-,W�v�n�s�ymZ�z���]`��-@������GYE۝�<���GHE�� o..�o�?�������-ZK�B��=���sh�Ğt���@��>Y}%�Ȇ��%����98����c�_�tF�|�d_�%�n�`	��B�`f���O�v]�ԕ(�z#�d{�#���\�h����� X�{4�2v�?6�0*C����a��N~�s~#[ ��(*KCYa���ɬ�^Rl�5UhX|��M��k���;��%�`��E�L�,.�[x�dc{oH<U<�?������Ɵ�(��<��M��Vf�Z��O}w�V�>�Y�Q�`�un���3��J��5mH�m��ʎ4<�	-��x\��k_�m�}0d@t��u1�h�'8���U"m�Q ��B���F"r���aOҷ�z�P�ՒdA�`��p%Gq9J�e�58�WY����NN�d�*�A���,��(��a�r��Pi3��<���vӢn���bn&vdyϟ��!�~�w\� ��h�i��bL�,O�e����b61d5��j�P�rko�ņ5����r�ynn�tP�zo���S;2��n:��]���d��f����):�-�TDH��#�N����A�H/l�@ڴ�!�_�z��S��+p*w�.Z�7�Ծ�Cd*�X��w 2�bR�$b�E�h�8cG+@?<�6����v����Nd,�ca`F`�O~�Ci�G�m��X��7�^{�m}�vTy������`v���/~��.�Dz����3x^v��-�듍�gT'�Gv���\��ﱯV[���r"kc�~�|#������Ȯe�R�����(C���$>dyVp�M���3҉R��1diL<h���Cm(K���c�N%b�JX�#G�5�.Ɏ$�{B�]CR��v�tJ�Mw�r�q��2�:�a��o����Vथ�9���+��V����L�[���Ѽ���a��xm�s���%��4�Xr�� ׸���@ylk�21�����@��E�s��Ċ�G�E���-��š ��a}L�]�����j��� ��c�lA��3��s%���&�h�2LI( ���v~�8�#��Q?��_�E����՝Y*�tj�=ڱ5��JK	���	 ��o�lP�y�(�(Y���NR��ȓr��I�[w�/���Dd�����'����M�>\v�6�o�v�e$�)�X�I�s��Ӣz}��k��`1Ɋ���0<a��q\�J%R���e\�M�>s�M[p(���M�
ІLn�S]ѭ)v/�\A���[Ct�C�%T����]�E��|t>v%�F��`7�R�an�����'0 �H;���pi�|��:ӯ�J)�F֐^� _}
}th���N��ۍ�P�l���1s����]�/��u�lx�w���v�K�
 �{��M��P��&��_�03�%�ڙ+�6<�v��Nź��3.��`ȭTo�J�����	{_4z=���e�[�k�1��?�P��S�xͰ3'5�� t�#��qL	0""0�H�W�5�-�.\\�[yw����j[嶼�p��a`�}���+����W�W��aHk�6i�U�](#���A��ڧM@gn��n���ga�ί�K$[�O> Tbt	��l]�i&v\A�
��FW-w_E<5p6+r���O����6��N�Lg�ͫ)H���Aob�+�!�[1�V8}dH�o��n6$��AYM��5�A�����G�ʮ��Ƽ񵗵4g�-�0)W�0���#2E}	���eRJ~��7����5�$�}���V��'LA��4��j�4aam�n������yU��C��{�d@5�����d(��J�������چiG�������F�N,�"���t��d_�I[9�%dw|8ˢ~��aL���sq���R�@���)>,�O���Y��BߌF������L�F/f�o�2 �����ME�UA�ob�� ��@�l?��Sd��+F,��@]���Z���]�LvЋ�2��|�8�7�����TR��ѽ��~(Q<x��~�@��יD�[��oJQ�X����^�C��dM�X�a���7��W�]�l0����GB��q�R�9==�p�@�]�
��$�]b���/&��XW�Z!� ���/�o�I�n^�]�3_&\�c /b�g��4s)�E��g"�ȕ��qV�>E�uA�ʻ��3��[�x-	*�!��ε⇢h2��|s��a�yV���|+�$��db�����ּF�k�<�����HZ�X���Z���b��]�4�:�	F��}��8,�V
W �>suFO��ݕK�y�����?v,��d�2Q�7

	���,��;��oڭ�����l.�������g�u���I�ンg�7],1��j8�v��`�P�P$�Zu�4�� rK!������s�H�^��{��;��\�3�����|m�T�E��c{���9{S���޵u���=�V��e ��ƃ�4��?��K�	KZqg���r�B�I��_��N�5���D�z�4s��@{?p�������7}��C]��Z�h����7`vq��|�y�s�S6[q�KC��k�b�T,Y��*�r��ls :������lt��B�����Ζ�=ռ��'�{(=VE���cj�h��� ��S�98���m�m8�Q9�8�����]��DNû�]ob����yܢ�}�۹@)�Z�`恘HAX��~zD]�d5K�-�a�G�HR	��t�hͷ��*V�9Z,=ݨ$���nE�r����)�@L�H �Zo�c���%�YCY1�o���2��W��7�B�tm�f�a�78����$JGAT�=�/%���b��)/.#Y(��$��f�Οt� .��Լ�Ҵ���{�'�v܉����4���Wul�W'�G	�����e����ٽܛ;�~q�J��أ+!ͅn�ކ3y�-1p�l֯F��?�iYL0��$ֆ�f����N�4�$J#��L/M�d�R�""�Fx��_�S=
,�b�m���Yߟ$a���^��ފ���`?��o�g�#��W�%�(H�tw��b��L�r�K.!G�\Yd�;���������Y�e�
�T�����|�2�ra�+>t�.��8��d 6��XF��?��w��@Xx������U����p�;��I�Qn퀘)�� C��HDL)$Z�������I��]��O�[����'HU��D"o����.���.�XǄH����^Cow��n�`��Q���������c�N���
�O�#8Y��Cq�^�g)�\xO.��+��Vq���G�m���uڿ��ؒ��6�q��<Wm�s��L�����ŋ,��͍�kn�^+��h�ڤ
.�j����rW�󩼶��V�������S��^���sʁ������r���&N��W���D5=/�n��ͻ%+�hj�Hs���f�/Q������C֤����\aL=���ɡ�$`�'��������z�ֳx�g�-~%��f�Wٸ��>F �&TO(@�t�H*z����ߜ빵���C>���y�6'���H�����]��n����/L�~��*;�|PCË���)N��%���~�p�l�6��y*�)3sE$�<���[A4z}[v��A#w�(V�Ս�$)���U�nV�A�4��`��d�{��/���RĎ���%�FxP0�2�[��;��bm$��X���6��c!�O����{�#�Jx�	f!�8����?
���\����74Gu�7_��H��@�����̅�-"b��9;ɮ�dt�*h��~ņ��A!���c��Q�٣lL���?5��]�KEC�f�����:�Ԟ�܄\��6�n	�R��CP���H�&4,�$Vt���[c��ی�u	�z+�����ou�b���0 {�U�s�%F��N_g�0��v�$�(ۍ�a5<n�D��~��Eo]���Ɇ�^��]�^�hv�~1�yLnN���Q�\�H�uj��`��k3��C�#���,�bn|o��D(Wz!�'-���d̙�ۨ���F�N���q�u�JΗ���M)/CMB��eZX��R���{��p��]F��MN�^6�k�x�<�7�*��6�zJ�9�^�z	L=�'���+��ʿ?
fÉ�M72�NM6bz�UQ#��.���C�������^��V�!_7>���M'6(06�nQ:�>j�V�w�ȇ��E��520��[)xIn��q>�?� .O��OM7�nDh*���'��(^�.��g�
@�~Lì��c�M7iQ��V��bu	}�V���w�h-�F��;�K��RŶ,QR����:�'��j�u���y�-�JMb*��$R�$E�+`=���E����=�s����D�1�5���Hׅ�13��D�2���6)z�o��Z�-�e�E�h#'�&ҟ�/��``����Q�;q�=? $c��%�/�@��������)��de(l���@�ڽ�wf`÷f#�$McT�=��j����<%�@ƺ�������=��O�8$�V8S�|�<��C�q���2T:�"m����U
��&~��[N4Է&^�ѽ�2	� �k�p���j5G�X惯��R�;�+!��U*y6!��X �EiekF��҅�auf���h�b�w���sŮ#`|�Kt���Y�3[Y�;�YV6�謁%d0��
é�j
8%\�?��	�ƶp���1ӌ>�to~�~�ܝA��@RR�o߇������fH���j���#��7}��u]����Ӑ�R`�c�F�dbyrt��O�X��/ǰ-���1���f�H����Mf��\7��~�X�J�7�cȀř�XD�̶��W��b�x���o��dšَ���,����aYEz���|�K��G`�4��G��E�$��-�"Ț��� ��bk�����YU�i��ko?f_\�B�k7GalS���)<��� �k�zI��b@��gP-�A�^o�6�83u���rD�q�����J<�宆�&V�w+
.-�ִw�eoT�o�Jf>O��b!��@�CF�Y�$:`�Ka�)n�Q�Ao���3� ��/�@w������Wf^!o&m%������Q{|�/�����d�t��<n��� 	�C�%яg9��k�o��QY��M�-_Q�T��um��+��v�X��cX.��f�d/��8��.!�Wnvq$��oK�Tq��I��"�oC"�f�uT�!�e o1���6���#9iyseW�?'��1�1:0"���{vê�O5�-1��`{&�d\��mI�£7�c�P�5�`f� }~q��/�Ģ=�榼���柢��E$�X_��S�ۉ~�{빙��5zm!;ƫ/�@?�h�1S�����U;.���Þ���Ʋ��a%�`��������O�Q��v����1��aph�c�$�9Ik5��<]m��b�&>�ZT&tl6N���&[s#���q�ݥ��r�㥔\��B��[$p�'§
��1�C�y!��9l:�̞7!k�m�g��N�7�o����R͙W�1�_춒f((�ۻ�G=�e�1� H�Ox��N��v�����T�P"N]���<���Wj~�B��!��m�-��ӻ����iZQ]�N���L�2o�������9����|�-5k�t��7�^<�/�Gұ���Ѧ��'z�'�#X*�3��VIG���~[�p�U�]2���گ��	�v2]�2�pOȚ,1j�B��v�~92|��@��������	5l�yjXR�G�tI�@5����-3�����a��?�G�޷š@�^��K)}�-y9*����A<�&�#ن1mW�n��@7'_��B���@��a0g��<���,�N�kФTD��>�	D�?Hj���)����{Rz���f�J��,G��a�a�'5��W��v�ZO�/��'��+�!�-�bX��9@Yw",+G|�^C�y���X3C��S����T�f��B"�7ֺixq8o�ܩ���.)�l?JЛM:	�܉�PW�'���P䯣Y� �:��p-ԕF��K�� YO��C(:}��!"��W� `1�ܔd�0�n}���\F`�Kt�AJ�h���+�Ә�El�M�q���j�����Y����A���+��j���s
�S���e�X��W�LjU��YZ�.�7#�Q�+�|�I��Vu�[\(ot��������-y�+&ס�/�{y�
+���5r5=[�/M���}��ɽ�s(��n�ٟ ;ZXt��� B?���'�L�w���4���[��[�P-(��P�g%�����K#I8�W��Ϙ��_�}���dA�0_�X�&�'Qx6�p�`du�;�G��\׭q�כ�|�,�}��Sx^Lj�T����6��abJ��h�8�n�/������*u-y�S�(3�RUHv�ؒ�����#�`� h[c��`��d�+3�����o[�nA�[�^4m^��f�#G&t�E��L�����1p�����&��|���rq�zoH⊅��R_d�.��@����`�s�7O���HBUG���Z������5��X+TV�����x��y)��O�O�* #o���.φ��L%5\_�k�
�U(�h$���ã��_��9W����[��60fc�T��~t��U�'۸ٹ�J�H�����\�;cU���͕%���!�nMǚ�U~�����	���]S ʎ�*��1�x(��C&9wl�Z4����Ә�'E��7x��,����`��l�8y~�F]^�I���+�%0��עZ_�r�掹  �K�/P��W��W�-m� �u�������4�Q�$��C���*���<�E����4��s��i�s�x$ҋ2���Py��Y���+��~�}�w�	�q�e������	�� (C^�$�%�k�Ī�#I�{�O<�bgm�2x����w��Dq��0A�4_���"(�$C���vH�P��1պ֟�)F�_�f�捰/S�T=������38㵊�h��ѥE4�ه��V#��6S�<��gR���p۳31��X��T��1�;[��Yr�n��m��!Tj��7�o͎�����u�Fj�Κ"uP��n�D-�ݷ��p��8������y�������5�m�uL �?|�G�Ib��w��8��nF6���)mX�dyQ�s5E�wX���#Y�֚[��m��Az����9�n m������Ph��K�3�R�'�5*�ϡZ��R=:07�G3���5h�W�1�����0��-)�fz�j��~�Y;�Ź�𡎐��E�ܛ��]���9�E��
G�E<���GNY����W!�k����&���!�z�_�I�p�L�n�<��|�6I���2�~] ����s�F�_���S���U���ڤ$��E�AݘP$4�9��d������>����w�Ln���|��2�
��uU�fF����@�u}�)X��%\�����@;]���XV���N�!4#�N~Õ�*v��o���ם�sb}�/�c�A�K$�a���0��Va,Z��E�R�"J3�T7��˼����[-(��?�'�n��y�Nš���.9ne�4��#/��r'&o��</��e��ظ#/��y#�>��j<n��?�De�pg�S��J����(�,�;Ϭ���x��W!�M˪aT5h=�^�bm���J�إÖf���Br	tw��\�h�Z�p�Ԑ�&���ͺ�rL����!�Y�te[��(�(�x�9rv�n�p�#U��*Hmg��ظ��Yag�P�.8R�Mi�/��o�M��~�&fސǙ�T, �^<k�B�!���{8��ХՀy�2l+EyCP�5e4sm�Re"�t��ڶ����q}�;=��Ҡ`�x}���gi��jQh�"��I���cL_�������Q��o�G����N.ӎ �̊ax2���`�W����E
S���i��>Me��li�S���q����,��f(Ͳ�m����{�K�a���� |�+�HB�����!!,iX��/�>C�z���E�h�!jAJ�c�,���)g�J��Z�P9=^�Z��>�����D�39����(�*AMN���|��Y�= ��r�n�A�d@�L=���"_���������e��\ZC>�^�7�}=���@k�� ݡ+r�����I�l�*��ujtz�����R�A١XL�x�p|9�	��d��k��Ƨ��3���5K
��ͯC�&}?dhf� g aKBG�-��x���um-7J'���}���<��	����%�r�C���=�v�}�~�o�py��h(��"J��6fT���V�{��[T0�l��c5��2P��[i��ap��"c'�`f�~=����B�߰��^z�� �w?�<AqTt��u%��D��}�c?����-����U� v=m�	s��E�7vM�Tߩ�w�W�.n�:��V����:�O�ܭ~�\cxC	&oʒ�sVį��u��h�h���C���5fz�{��װ�jM���#�K#HN���� ,�9�@�5�$����� ��D���7�{gX^�|*`ɝ���V��u��Kh0*��ԭ�����c�S_Cn�ʯ��52���$.{ �9?��!��ݱk؞5H�	>_K�_ϴ�[�L��}�7!�.��_��%�왝�Lo��N�"��x!x.|r�����`Z�_Ts�s2�m��O̵\T	��	Q�T���:��6<����,�����6��F�<�Iu��ԝv+���T�1*�����#��B���f�Ѭ���[�V��!j&�R9Fv��f�{��Bw�����]��!R8iv��+S%|}���S�����݉�9"���ֿ��V�����)�l+:��qXpA�L�%|ǃ�m.qt����=��XG>��RBv]1��L9U|ق q�Z�Q�F���V�=��������S��9��*�B�X��LTWhZ��^�J�をN��ݧG�P ���yQ]]�E�o��"9D$Cbyu�PB���.ب�6�4	6�=Y��{5��Q+����O]MsIv �JD?�A��.�6a_�	r��5�������'��z��>�r�}G5`
��i�sv���z�1��D5?�5������PC���D�}*s�0��J�4V�}��̿��$<x��q�A�*��`�M��-n+����$+���8�b�X�k
do]&�2�-{��~�o��&�S�ߧm�Kt�@��?bY�+�ʠw4�Q@�N����ё#R����1�>�G�L����p�#{����"�x�LOw ����3w�I0f"4�[�9Q�$�V�����<���Ng� qo�v��xSt9�-������ԙ�!�84�V~gF?.x�	�l��[ @���,HS�)�V�_�/|4!	�eF����3�T��b�A���k�vF�{{����'d@����n�|i�S��X[_����a¯�6�\6�n�za�^2`��WE��x�7H�#5
EVLYW�=�cg#�̑U��-��N�}�����6#l$�xxCx!��v��Q�8����ф�/�x��1m���n�[0Wyn��x�V�3R����<�����=�e\'�E��k��?%RZH$�&0�����ʵ-#ӌOk��u��D�jc1Ye�ȉ�$Mw{5E����0f8-���,�O��)7���x�헣���>���4X��,�@&Hl���?�'���u�i��!��������u�FO'c� *�H���Ʉ��g��T`]��e%]�Rz�p�Uf�^�D��kv�d<�Z�Tw�R(�<K�4�u��ū���6�G6���<��6���'��6�ڶ��VA���W���c[+�|�I�߱ˊ��*��q5�{��Q��v�8RL�nV<Mɥ6�X{�P�d��n26�-j![v��&���[���w�Ru��2�Z�g���:��}[>����\q�QtZn����͜�'��)��ʢn?��@E�x������pBײ'Jo�S4-ޏ�WH���'�d�~�>P���d&N�L��k��`{�݁�:�a�4���.ȞWz�P�J��z^QW�6j+OH�tZ��� �����f�������a.���. B�����A�ے��&������a���Ax�s�35�7�iA3���������I�Qy�P��e���8�K� �OeC��q1��9��h �o`c� `�@Ǩ��˴�~��E�9��,�hj�8���oR:���R��pH��r� Q։�!��,*#B��k���!c��BOw՗�5�6{�G�f�	ݣ����ףR���3���=��M�(���`W3�P �������� ƜaW�����<�⡍��P�]���;v�W�ˀ4ʜV B�A�W����\���|�m�_����F�H  e}`���1��
d��<�Z�b'sM�[&��\B�-��L�	}���ύ{�)����&�\I�s�1��;}�Db�����Qz��>��zX�e;K��ϒ�Sl�kA�L�z!�uiF����Mho�[�Km�rU ����0�����T<�V�}�<��xb��G��o���l�Yu�!pK�ɏ�[��%iA��h���p���&7ɴ�L�|�= �0�"^��}�b�n��l3���/=�S���o�������o���]�F(�.�� ��q�9�b���Yi���\����z�g�ͲVC��!k'�(Q4���aQ��s��_���,��aZ�ш�_����|(���^����1bze�zz��8��_]�H�U�W=G�Bj����LOR֘v�:�^#rj�ɣ�@;��H/��(i������}�ɁF���Q�,��y#⭦��s�J�����󽞯0��6?��v�V�Ymv�`:���`�\;nR�3գ���!M�x�\_fu����P#O̕͞�t��R*���~+UE��w�ͼ@���NV��P9��S��G騰��B�� �~�T�6�g����S��R��3�j�����v��.��������.�]"�K��/��V���v���Ȳ8۶��D|� s�$M�!�����K�lf��
���kk"���D �J�_�p�
�� ,ϦEi�Q +���G�r҅��_z�����/�g�Њ�b�Z�Rg�؟�|���K#�2�S�b�⯛P�J��߆��s.�,���a˴�C�;�MVGۚ잃�KCj �����[80�՟Q�p���3̔�:�=����߰I�����%z�&{m6(����:۬#/�t<e��-��I� ��OLڤuZ@"t#B��y�b�`j�[a(��VjD|7B�Օ1| �̈�Ïy�,��L����u����&��}n� S�]3zR��m��/��Z�QzXw��1R����ưI�9fI0|���8��Xf�+b�c���ǲ�UЄ���9m�.s"鱧�j�f�8Ă�KǶ�;��+�����ef�q�����G�����!�g���჊^7��5?(/��-L�"n��#�뭗��@K�K�1��ֱ�C�AC[�@�L3?B�0�7-�P0,/q��?!�w���n�G�W�u�{��Q��f׹5���:��^�y�qU)dC
�>��[H�G�kg���c=�'���yiؙtn�Y�9��V��NL(��>�]�.�>�|���f�M��R.��p]y-t��C?|�;�2((�R����`W��
�w���C� �!��������l#�Oñ#�+�.Ҡ��d��5�+��-$f
���vy;67�$+��T��E�j���y��
��������B	�+3���f�-�ܓ�f ّr7���	8_Ќh��Oᶭ�F� �;/�Q�Y:����q:�	6����)Ù*���)��"�)��*R�ݗz3�p^o�kh�c��h���d�k�dǜu�R?	����h(?��PQʂ�������0�>X�躾��<��2��ho��~���[s���:�-��X��)!|��0���s���p���{D�-�!]��޲�Q3�<˹�H�5��j
[G�B]��d�*�H��A=����ʣ��N�i�O/*30�Q��,\�#�.�8@5M�d��"q�^
�u�����E�.o�1�g��D�@;$���Z���
��w�r.���$ty'I�[R��I�)� *��̴�X��$?l`��@�A��v�%Ձ8,[`�)��$�����S��a�
@O��n͙
����y>�}�;f�6���mSu�ΗhX��g� 5e���\� E;����8e���A��������N�sS�Vz������["�F�v�0��r
\,�Vڔ��Ϧ��A��Z�����Pb�ЋY�M	CD��<
�;H$�ZD/�c�qւT��O���k肯(ʣ��Z��Vw( ˳J�+�f�ůt�,����T9�D�v&�z�k�i�(&���VR]�t[�F9�hI�=`�
f'N���QG��v-3E��8��ɫF� ����/J��?Py?7�\��:_dL߸�k�%�%a*%F�0�h��; l<�&:�zM�8�Ǧ��`�.z �=����oڍv]mL�<��h���J������ݩx�>]��S6cýʁ�vA�X�\�"�M�_���:�*�u9_؏���,vF��y\.RvzDE�4T~�|Rd����<��A]E/=ٚ�bJ���Ju:���s#ҝHUp7���R���k���v������됓8:��H�3/U�s���#����C��@T�!�Kξ4J�2j�匢�� �8�
���!��_��AJ��U�a��d��H�Z���+	P��K��L�k�5:��#���L�b� k�r$��la��u*.���d9�뾯��9`v�%���P�,�7`:�}�x;�ͳ�	��)�uГ�e���Ju �We�a]m
��B���0w��~�ܨ�K��1q#�����ZSڵ���h8j������Z��`��vO�$� ��ݫ�h��
�Z_q�aO��-Hs��T�ؑ��+O/}t��t�D���;�Y��nz��Ԧ��:��g�5V趻fd����X-5񵇈� �U�HY���m��Z�w��5�샃�c`�W��%q	�%�n�[JX,�e��2ۑB�,X�R����lhu8��F����Ⱦ]�=Z�(�By�R��S��������z��nd-�b�N�^ ���4GdR-ZQu��~�n��g�dU�AC������C�wN;e����#߬�
���Vw]���\��I5Y��n�*��‾���(0;R�5�6�z���ޘ��&�yN���u�B��*7)0����?�G\��a�#a#��;͋s/�S�gz�6	�g+MT0pS*�ܐ�3�buv�|�W o��t!�"���O�1���{�~������*D��v�uh��AI����P���M^��*�
��Nw��6v��B����C�V��cg�����+���M���)��ۥ��聫І��v���&�����p>m�>���|�(|�$�<��4^Li<�6���
��ɻD�,�.�U��͑��i��hq��--�ޑ{Vl��J���ck�qôEAl�l�*�2�����e�{{�: ŗ�m�(��� ,�`��,�E7��Vo[Ԫ&8�Xg?v��R쐆Ǽ�6��%y�T�m����=��#g9���U3p���;����J:j짗�v�5a�ˊ�*�ؕ޼��Z^�w��]^*���}�8�:^*�95��9�rtm�|����0�)}��+Ǔ������t l�u�DED,��V�K[S%�[*��~�kt�!����b@�2E�pzQ�xm5��?������}	�����7�Ld�P�"�,�)�B�p�j��x�>������� �A�U'��j�!'�u���r�O���-!���G�Zԧ���qv����l/��K�j�	���dΊ��+nv��'�.Y:z�����#�ϺD	�ԄC�଎���c^Z1���T�F���_p��oŧ�z��Hu�-@��}��j��bq���$,��5��������kٺ�Ch���� ��X!Tr���{u�Ue6lջu�P�Q+�?"t���ڨ��9g$���}�qD8��̚fڡZ!:Ζ��J�>/�ut����c������7:~MQ�=��'5-����)���r��C�[�b�^�OLZ(��w�&��Ь��a���U�؀�P�H*��]�T�i��<[��.�����f�ܱ�O��i�ԩ>��� |2�
�1�se��Ô3�0�"�x�Jd�4b�Z�H�d�{�/B#겤j9-l��k*
.У��h�	rh�,�  ׌�"X+�����T�֯��ob/P�Y������M��¡>�7)b�bXx�l�x��~T�w��w�9"u�Y�V�WM��Y~0w�f�j�i����`ru���ء�1�'���;!_�±��DXӖ���x0C�on	F��!�,��:<�\�{��j�ۡ';$�G��0)|5�h�qP+ܣ�&�/�-��y�!}ܓ��'���j��,	(ڰ���o>��{���8Z��T��yc���.�Pݧo
f��gYG7��b�џYi������4� �=h��I^K�E	�1�>���5�A�q�6.�*K�rK-}�M���윩��X�F �9!g���^r共�XW�T���`�G
(�8{�eT%ݮ�v���
�tfi9;���A9����g����Ͱ�J��}6��+��S�*��xoy¿"��h��z[�^YB����b��?��@7CB����; e�����{�eYr]���f"O���P�Ku�k�vC�/���ʒ�AH�@�'���WF謡���ҡ�体z�%Vk��L�������V1�������0���T��.�1���v�����o�)3c6����2W\�[,��rl�z�[�aQl���xa@��n�a����d� K󂊺}J��7�=�^��	g��=����>�!���oJ��ɜ����w�nW�իw��8��S-',~����_����뜌���www7~����V\8)s�\�������tG���������`x�T;'�UE���d�J���!w�5����b(6�Ԃ�2�]ǂ9��E�sz����hT��$����/JH�F_�H��M,�	]�m7�J�19
Ϣ� �%�4�lIV�E��_Y����q�ĸ�,ݢ�I)d��ĸ�U^��8�}Q]�
��J JJMve���9%bT���&�nM+�v$����P���S�"�*�!��M�q��Oeau�ya�AC�p�`��!�[<�����\��hC��ʇ$���ERZ�Mҵ)U�	m����i�_���갣�;E��w�38c=p�%�ʕgf������r:M ld����PPP*���5�T�Xì�k�0�H�]N��j�ҟ�)�����]H�.�S�yJ�-�R�r�Rr�3S��	̇}[9(9i|��Gh�F�FҤ_h�G���58��Py��3�u���A{خ�B������c������u�.����&�ԙ�hJV�셠2��.0�$���<�V��PІ[�����SPN頋�qQ��XV���>�4�!Zq��}b�b��h(�&K�
N6I��~l�*˰�t���l���[3�	�=��u��g{$��x���i>��`����ڊ���؉&�U����䐋�O]۴�~D�.]�T1R�WN��o�lk֭���$a�>�a��˸P#P�����?�!Ejz5!�����;y�*7t��4��BŁCw�L����� ����m���r�^���長�VD�U
44w.�Q���<g.�U�@(땂�$�S���I��Ř	�t��g^94�a��y;R�ԅ�G� �fc͋�SV�`w�Q���\vPL��e��mb�ϞCV~YJf3�}�EMn���X�K�d&uȺ͏��?St��`O]N�/V�`�@g"G4b~��Ѥ����;�Y�������eJq}��I2dR��ɜ`��Q)���7�h��Qe^�(��G�pA{j־���ŀ��+1�TǑK�<�$�Vf���P�(޿O=�nخ��8�<}>�/xW�2G!A�pD%x���z[�{������L����(r�Z��B��oQ�Y5�S�
�~̸ �:=�;
�D��H��F���l�2�τ��|�� #Cs��kG����4I�70ߔe��c �`ԯɗ�9�	��g]B��b���>Ż�cԪ�������c��r�_$?��W�s�dxy{?����=:6�$�ǎ\�|�u�#� ��5(�᷑r��[��l�u�R�� ��t��L��H�ɀ���iW��G�%}m�Oh���J�jdb�������G�ѓ��hO=���R���<yT�˷����ߩ7���_���d\�09��hBH�P����; ��y�'�5|�(��a.��w���K��-��A��:�Rp(��Z�*�m�
�3�H� }��vb慖�<�W+�[V���"5_ڻ���ox�[��w�R*(�i�h0P�������6I>��Өp�p�p�'f���H.��o:$�6#��)�%���gV#v}Ch��Sv���B؃�[��w(����/d��Y�&�Ʌ��4G���0�_/��iD!y�F�`�WpX	ID�m��An�j���)�ĺ�'�uġ� ��}.�]�����N5��R��*s\(�Q[{��� ��y�O�W�l��C���{��&Pn#����ä��ƕhE�|��R:�$�%��������X����:�q�}x]z
�Rp'Y�.͆P^QP�D�ī��;�����[�O��*j�/�u�YkUh��qU��6�n���ԥ}ā�gKYW+N��2[��s�_�k\���.a#�2����<e;	�q@V�i4����^�V���0r���/?�?���������+��gɧҰa;I���<4k��2iZk0X�q��Qz6���/�_��*�V�pA�P���Ί�`wrE+�j�;���@�A��d��w���Ʋ_C���6���ȓ���o�us��AU��\qAv~[��}ʲp�3���r��=d�Ks ��t�'d������������v�@��$Tkٶ��Ae$�It�"q�H["�٥uK����-�coi��?��߇�:3M�~�-$�̐��ĕ,�>�6㋐��	�r{lc�q�{F/�%�d�-��|��i�䑽<����O�E��{W@��������G�lya�V9%�7�����;%enJ�,�ŷ-Ve2��|�TF*Pw�����`n4�^8Yl�`�����?�O�p�D�ǰ�J�nE�%ɵ&F'A��,���/���(�t�S�pQl������xH�Vݨ)�����d^�Q�[u�롃#�9c�$�=Q�̖�F'���	M�^�Rx�>��̅�w��|hnC:�����6��>S�Ʈ�	fSJ=��憘����z�����l������?%����,���E��\D�?�	W_א9i��ˑM��9[�QpT��\� ��۝���~IOP|����� aNm�&S��I��P1��?�J~i�;=�|�܋}�3L�Ocp&J1���$d�#�Z�^��;4kLc{���8�9���x@���_#;g��l�SY�(ѩy,u}�O�s6(�<�[b,4���XE(� 	m} M�Lt���8��w�X�ihZ-� n}�!�JH H�)ǘb+eWM��k[��Q�$�c=^�-�����넗�� �Ө�c� X����sd�7ʝ;�cK
�)�LT��u�Qz`��]=�-s���ޥ��0d�s�	�*�L���W�N�
e�f�xf-�g,m�(^��^�J�+��,t�a�kӜ�X�%%�ê��;�/�<=����L��5o��l�+�!:%�V0�1%����퉦�%���ҙv�N���t�W��C�����׬���
t�(mѾ�Y*�;�>�Ĕǆ*)��A'��X��b�r���|�jb�ӎ�;��B
�k]�;�����O�O�a�c�}ADŞ%k����2�����䓸b��$�s��> ���^A��́Bi��b�L��˻�.�#3�׹.>Ŋ�J�E���uf��i�/?�%���h�^�XHaC߶/IATI��K*d��9�`�M� ̢wu��L5NϦ�>{L��Mr��@���kPlg�k]h������02��gW:�:?2��ٸ������ea����H%�j��W�����1)��SQV�ު=_u����^T#|&�cs�C�X\��g�}#X��g.Q��~r�~��5zֆޒ��&������� �GV��o���������á�|���a�$����
`!�u.0��!�4`�E۬��(���űoe:�`.+gAhC�q�x$�Y�� ��(�� q+�ީ�(lh��y�/؉�E���������T�o�'�Hc�@����lQ>�Jt��	�-�n*�OG���9yJ,� ��qnݣ�,q�w�6�"d,��eW&X�"�{��x���lg�m��r/'iZ*�D:9y�*�ez���.�"xZ^]��G2k��hD�).�r�z��%'A��+�����-� ����a��o���-m�U���_�@��I<��"֊������ ���EK��$�K����ʹ���Eb��S��Y�\k�A�EG��գ�5)H1� ���GMt�Jϑ[vdԽx,�` �Om���I	:��ug���3�CԡL\�p��I�ǲ��b2�C�9?�F�ߒ����Q�s�C�S��fĘJ,NV�2'�RT�v� �2DN�If��8^BhI��2�a�G3��i�O2�vQ����=��� �1� DE�1�2���Z!h��6��'<H"x�.#���S� �|v�\*Y<i�Z�X���4������8��W>�M�k����]�����K������kK�Du��Q�z��Q�aKP��r��Q@�����5'B.t�����\���b���I�?\�O	+M�*@$�)�_��١֤$�SȌ�ϥ�<�}1 ��)��UCF����a�s�K�������#i<��5Ňş�V1PM��7��s�9�B3Ė���A���b�Y"T�oa�CM�o�3�����_ٻ��be<�VLR^2aI�c��'KpF��]�_�RM9x�PtK{|x��{�d%{���z��~E{�3pР��c�M�W0 zYEQ��UP�S.%�Ƚ���j���ץ�K�������c$�A�uN��;}�F�(��l��|!*���H�HSx��ܞeN<�J֑,�N��c��1	
���3�C������q̀����d<h4����+��C'��P��J%{9aŇH�������U⍌�ʝ��X$ω��|g�3k� ���d�^��H��fSE6�+df�U{G<��~
�S��l(7=��:��smP>��0@�]�f�)�"��!E��v���H�IV0$9㌀��8�yT&�F`&�g `2"�����9������P�6�},#u�E��~gN[1\�U~�صzC��)��ލ� p�i\��ʓ'��B�.,H[SW�8<����� tMlT2����(W :$x6�>"��mz�ՌAvW�����W��>s;N_$��/Ͽh���p�H'(�x5��U��۫T<�l�!<�]߆�}�@8���<4;�����~����tB�3�`�-��ܞ^��+q��c����@x/7�	i?��&��@P'qOGb��b�G��}��F�EV�1z�b�m���Ra�Dڑ)֗G�o��oH�kxCv+�Z�0�7�r'��S^0<n��d�����KX���ZH�&Ern�w�s^/|��[]E��w�k,ytL2WHL"~�E.& �,��˰`�s�i?¼ɮ��Dxap��!#��m��o�.b�{������d7N�d��b&5����f�3_m#O�"�x�=�-�U0���u_En�Q�>2��v��t<�sg_�m�,1��<�p�Z@�����!m�j�<d�o h��:i,��>);�% <��\@���`ۇE�vж��`稿K_�y�v��2�]E����,�����4 �:n�b�uAچ)f�z������e"���?@���:�J[�:Q�P/m|p>~5@���ud<��GeBǿ�ۙ\]�Oc�&��ГO4uI{`i-���P�	�a�'SZ�&E�o���ߙ>����Ýgo0]�(_,xN��y2���M3��]��:�u� �ݵ}���i���gk
�'�;u(M҉ ��p���Aw+M_�j��Ey[K�=T�Sja�k5�#/�}�����m6�5H+N���S1�w�r�]�x�d���C��w��w�;Y��ۉ���B�ڱ,���ƭ�]�P86�:�4[�((�cP{����䋍�(���%;��G�%���P�����}#{U)�8�h��=�a���|+,��#w��O��Ԑ�B^v����j����:Ų�=�rAљI/�p�/��~C�r�����eY����w�~���s8�<�J��}���ϡ��f��m�?��ڎ��R��l��/ǘ��~�{k���`j ϲ�i^�O��]P��w�t@Qs�*������q��Ӻi�C[��l�kyc�ۿ3�B>/�*߇JpF��)�v���{��I�>c K=�,��pSz4&=����	v��!��v������a9�uϠL��%��w�p���3��f/E��S�:j��P����@���$\���B�0�!2�y7�Nr�3�����8�=��KL}P�$  L\�]=����=���#{�:f{v{D�NFC�!�3V���%LA��wX���܏������n���Kg~W�J,[��~o��=��r@K�P�)6�	�O���bt��Ż���C��&����0����^џ�*)�b$�P���z��n�ء;.'�]q2�x��#��n�V�j��"1Y�]�����6�*�������=��Pk8ۛ�J����X�C8�&���5��ka���<�a���z��&((��퓧T���&X�Ϲ��u����Y�A��8�o<�����
~���S���3�DiUFP����Es�+�5���B����X����I��-��!��l�]�j�,�vɛ�Q]?پ��jЗ}˟ӥg�%wHs�Qz�6v�f��q	�8<
AZŵ���Z{B��ۻ�Ĝ��s�%9ta�3�P�d,�C_n��;���r�/�y�W���-��k���dޗ�9Ҹ �"֬�~�A��yt��3贪����������7'-��z�w����]ۋ~�D�jR�ޯ��8�bԿ���~9zu�K��b|���������A[xE�Z������0�wޥa#?�s�c2�v��t,���`�z��%��IЈ�{�	c��s钱㙿�-�@?�+�x��B���ꂞW�/D�����QM#��<U�.%���o+ѬKQ�i2�o:y�:I� q��:0���{��5V������IF��⃀��j|n�i�5��w�^[�\� �+�A�����-8t�z��N���;�ٺ�B���a�����[��Bn�K�]��/ �K������E�?�7e[����ʹy�Og#��)�h�;q��*�r� ���m3��n�V+�M�ц������t�+;e��uKr�ti�
O@.:���#8?�ۧ�N�w���.c�T��;A}(�7i�H��Is�k���&��L�yVߺw�"��E�3��U�1#"BS�c6Z �'�\�+o�f�fe�1C@�:��b�����[����9�����5OrdR��_�5��j|��w�z���ƕR·D�t!�[���f�H��H�&<�/��HȻ�/8�.�{|$Ո`�w d�>H��R���d�R�����!MCg�­,�i�]u�2M������}שF��/$��#j��@ŀi��y;��k������yl���Z]w�����hIR����{����Ut:I�i=��l�h`�*�!Vѓ�9A����_��b�e�Um�;S���W�"��JV���/J�}��X#=o���
(!�812I�?��~;Gb��^�il�h��F�������Oa�*i��Dq0Cd霿�?�^P�d��� E�2;Y�qR�9�I<�Sn:|g`��Gٞ���,(Nua�>Ϟ��3�-PW�����������{f+��|֌u�����r�٨�?K"�����C�L��DO�I������o���5�f�;̧�~��y��em����p%*$⨨jg�����m3	���e�W�@8����Ϊ�O�so�\3nQC;\ȳ��ޥ���13k�#�2P#��GF)N���@1�J��H�����XƬ90qTRhBX���(���U��R�5f��mK��ѥ�1�ٟn��VtuaM�8��*�s6.�9�-�?���M��sg%D�?�$���^�ٖڿ��Y+[���R��f��MEe'�ؖ�̍���$U8��5�7���V�8��݂4�ج�ۓ���$�py�v��l�[��>�Wb���v��-)- ��q���� ���m��IF״����o=h}f��>�#X�0��?��QK�~�q��	�M蘣��)/eQ��1�� �<k�*�Y���:A�uZJ�D�����MS���ij �F%����ͮ��"�g�\55F3�Y�o7��P��׻ ��zm�KL��L��?����-���SXv��K�45�"M�4��x����	�T�8�����^�Sڐ� ?&���:\:�@�s\�����v[5�~�K���7)����?}���t�1(��9��f8����
z7�^ۓ�m>,���*ː�=e�!c���
�Ͷ�F�V�~��D��r�`:���B]��4M.5���3?'~�2b�Ɠ7�r)�\��I}����m�T�x���������M�j�}Ԣ0d�	^���g.�2�P=�m��et�s�k�I4��"O ��ǈɯH?#� G5�e.��Q ��O �W4��oK!G&�d$:�^�)~�����FImw'����[�&���Y��0QU:��vD�9P�V��⡰���밧�l�@��W�U��Y�c��ЈL\>��9��㯯85Kn3�%L��(DL쌘%v���\1�4耼�qq;��;L�Q��zl�gX��ީm�u��WAx�[s/��0L�-��3_^��E�_��ý�"�w��]���`�Nܭ,3�]���0&o_[W!���ؘ��pC}�iDb����%z〈s��D5E6���3~s�]y�C������btuN(���˺�f�H�t�+����V�����v`��/l��el+��E(9rW�h�+,3#/���C>�-i��Z��(`|0�Q���w3}u��F�n���:�^� F�
M7��'���S-"�.��>w�p�c�IR���!�w�=2n󇳢����,̹�u��%���`�_^��JFF���}A{7�~����ҷ+\��<fH`f7(�Q����:�� ��o�I�e��rB]D���Ӗ�-�����?�����*����"�Ң���jy�$����뎠zIY�3� ���M�--�'��eU���?_ۻ3��f��u�9pr��������a�YGo��Q��ރ�E�9Do�]��"��e���R��ד~�1��df���jmQ��A�WR�̌�H�GfH�	RI^�rP�����D�]ZoMz
?Y?m��2����z����qm+nuO?K��0�E�j�d靱ܟ�Z���e&˹y!�S��?�^�� ���Saʚ�̣[;� g�u��_u�G2�+�|�<��ʣK���"r?wgd�����$�ie����3�ի�$cV#hT_.��D���8��P�A]O��Z�k9��P�qV���4�W����E��&�9�S�-u��H��#p�LF9��C���V�����x%���*����R��G��bM�f��%�D/�y��f�7�������r����O�G�� Й��o��{�9Ć�s��PPQ���� �a$Q@OgK'w���*�������.�ݬ�<�J#�#.^�,�N͖�L����T�~0NXQd 7�Y�֪r��	����t|^i(�l��,�c�őE�1s)���?$�J�Fk}<���W�D�4��!E�	..F�ź�5.��=�?�,�ի�o�i�Mu���Z��)9��D6�<�>���qxVN�j<�㉾$�	���{�y�iU������a�TY�d��_�P:.�@�@�k�Nz����}�ͣ���_~�S7,]$]��:U�uSĬ^���K�w㆔� bK���~sF.��_�!�˶�:����p���-c;��b��.�^�����pS%�\��I�3A*�{��}�'Y4 ���6Ü㭄?\�M��L�\@���;B�5���"}t5�6k��q����~(J;r����g�����<�"�ڊ΅��kq����¾"�y��:�do����D�x�U6�EA7�y:7� ��3��"k�q���K�����K-�"_��V�<�V���#��u�8���tR�
�
�S�³o1��@��W`����G���Z�K��v�� =2�g*vLN��Chbq� ����W�fJO/x+���]��K8�e:��sSz����[Q��� [���n`M�^Bӂ�q��U�f�ۛ�O%S�4a��i� �VaR۹��ܛ�4>X>�<'@a��z$�36��/Jՠ���N�UB�_,|{�@w��㽊q;՝�����a�A}T�y�������g\�od�i.��#0�w���^�eiZ%���X��\FL�@�����^�oW#t�&x���9��+���� 7��z����7����'ZϋA� �}ޕR�zg�+,A������O��� %���\��mE��o�����(r��������'��?k��B��]�F��9��Ƅeܝ�`�&-9�,[�)8��#�����(�[YC�7 X�����X�&����dVG��S��C;���ݱ�����JB��f;@=o8�wi�v(��K�d�h�N����Ryʊ�"���W�R貵��R��sN�Nw=� �S�bt��=�h�, �=qc��H�_b�QC��A�d�(��o�s�Fhs\��΁ ���n��G�s�������8s�����8��m\<�ņ�(1�[�}��_�
H�?�p:��W�"W7u�B)�t7�������0N�݁����h�j�B�(�Q�3�d�5�vf�W��Ee���j���Ei�TE�5�>K�!��*��о;�յM̊�y���Y�U�=*|�\)�^�_�+nwT���D�������ӎ���;�[��t�A�V��l�/�*�WL �
2����$�"�20]� ##�9����ث)�. �cJ�֚�e�L�w�:\��O�hx�Jֻ�`Y%}������^Ͽ�ވ�����P.e\�'L/���S(Ni��,>�|� �gOTv�����S 'W�\�����X�8n'����X����R=fV��t�3ʻ?�\=Шp�4��lR�*ȹ)p����˯X�n�=$����綒~ĵ�X�&���+�Z=�fw[ǎ����XB7�X"�Z�5,Xe��D5�uWF���8���Y��E��le�*%��j��B��_w�e�][x!����@�r�f�ӌ�K
�qk�:46> JYw�:Γq�����x?N�rY�h��-��DUm4�>�O�ej�<�ne����v���3zA|����fd���
.#L�> %� �w��`��D�wJ 9��2 %9���(�J���Kg��ٰD���v�ImŚ`<L\���(t�����P���l�Y.�_��(��ݤ��Bb��b\M:��xz����7[�qACtN|�y>����G˙~>��tÔ0kn�c�%tA܈*��enHAq��Qn�ר��7ѱb�ź����3嶴$�dL�T�Ѡ��b���P> ��_�\�.�������������C}�FoO���+�uP(�KQAh+�2��2�|�P�ehQ�d�;G�6��!I��⦐���*�������Kv`+�nt�C��C�#�h�ag�*i����_�cO�\�=eo�|vt�(��(�.����۽�ގ<�J�5��Jjt�2��Bn���t��TG���m8%:���L_���γR�,���ÿ���? �Ao��($x]��ȗ#���[��T�l��d���h�D=�,��ã���L�F�.U�+��s�3�m��u�X�������ާ��4?�͚z���X{�ϙ�dBȁ#��FP��p�<���<�ӨƑ����Ux#��rSM�~#`�N���}Hg�=9Bl���L��
��f�p,�yj��q���?Z��m�kߌsz�/�Y`)�E%��F�1��P�h�sW1?5��@��$��M=����)��p�zj(�bFì�,�Q��ٜ�`�����Z"�\
��K�p�vg�ߨ��\n�Z�=�S;�	�n�4?�<��'
ծCDz������A��$j�p��c�=�&(��(6����26�x�g�f�u�*�-!ȮE������^!��$*W+�6���ߘY Yg߻oRlB�r�`�lJ��J�T���@���F��USP�c�3����h��Ky����m��-oZ)�o��,��V���;wH�7������T�ިxdz�BѹI$;i���Q�_L�d2$4�Q�>!�ϧ+���:~��T$�E�b�F�m���lvqz�?9�V2����`��ůM ׅ�P�h�����~l�(�d���PlH����4x[an��%=�H��_�E#�Ĩ�|;������Ѧ�$ױA((4%J[w'���Kl�V�g!w*�U����DGD�	�d�y1j��ap�u��єè��2��+E�hA��X��k��gh���� D���A\����<�,w��#��}�t	`����-�
,O�̢��xġ(T��1�\"����=׏��<F�A��"�-��w���/�(�5�U�~".9H�q���o��Y��T���X3�38��`�o݃�T0�E��l��W�Y�@��y������_e�x!�=˨��Y�%0�Ố�����&�Gwe?��s�sb����4��\�������گ1#���y�h��}�:^�Ɩ��G�Զ�^��
�ۤ��h�Y� ���=H��3�t���QD'��-�Y�Ў���7p*�ٱTU:*"{.-~Ȳ�e�fylCD�؛p�p������K��Y���a"8�?��q�⹉Db�4pUoP�� �J_���'���z"h�\o�cA5md9��<�l˾pU�Zn9��
cyk&�C��8�9� ���E"*J\�%|>�0��HlmH�~(�p��!V�M97Žq)�4����N����g����~�Q��y*�ם �n�Ko���4�)�l�f�3��K�}���8��-�v��^��+��+~,)&��C�k:)D\,��������������qg�Ŷ��u����yj�����[C@�ة�(�l8�,����l�se����r~�nVWNE��xP�`z���8�"T�mI��^+��ߍ`�d'�4��zrK떱�L��ղ�\,~���]��h�h�؅��8�zK3]W���I��Z��f̫�[B�K��(�
v\����o2>���E֤"�L��훾�ַ�4&��T�ƁSX]E���9u�6��T#0��<v-��D�M����O�e���8D��V&$��.�Vm��$��d*�H�X�.��̀����3�^�qFiV�,��6���H.������0�֙U�0�N	S�XI|���>f���V���Ҿ�P�B ��0�}�)>�S�jDA����-��ͻ�y�A�N�E�6���ͥ�Ka�Td��8Ʌ�j����|v�݋��sk�W�Z�|!OW� c�]:�A���z)�,C= �V$Yl���9k?�*�&}c�#�[��z�>��[).�*=l��e����a��K�k�˧	d �C��$��?�ęE�I��A͛��
l���~;]o�˦�X�������fh[���}�px�� �EP+�|� u;X̜$��=cs]��#d�P��~�"�
 ��LdJ�q-�Λ�*���%�˷����P��Y�l�󣴊��^��Tk��S.Ű��<�D��Q����b��={�q�U����m�����ˊ:�n�F �(�zc�3i'��*c~k5]�y��oޭ���R���GY�!���t�r%ֶ'�<�vL�oQ�.7�獋e~�H��c��@2�\�u�}�Q8a	��z��;R�A�� �o�h��#��h#�eI�4��y�s:ꔌ�����9�ܴr����~�1����W��o���<{�3U d$ߋ���.�=������Eк8OA:J.���D%O�����"/��!?�A������(̐��V�Qp�0�@��
�;=_�#A�m��	{"�*V�3+��}�x�ք�����k�̗�)���:#�T݉oK�M�Oڧ)_ku�E�{<�U��G���*.���O\Wz8��?lrX)�f�1�/Iձe��,�6x��]ӊV*�Y��ݪ��S�!c� sB�O}8��2��p	��b=]%��Ϭ�D3�zfZ�0)_�vN��ԫ���NRt?!~Gay0XZ������$L;z"�h������]���0�O11����L~�M�U��d�a����-�A2���U�S/ǣ������CEɊ�����G�uح��R�$�}b>1	���|l_xzK:��O�x�]��J����HAE�`Lh���f�PF��)Ё����t�`t��D<���f��|���^��'z6�
�зU�t��qRk/�jM6���9աN"��"�&!h,��>5뮤1b��&2�̷ю����ؠ��:fo�j�����ރئb R��oN���y� �3�eS�ѝ:��y}#���` �G4���.9�������ԏ����Y���3�kˊJ�gLcH�W�P-L�ւ&��p��{�*�wQ�U���!I&�82���笩�g�yd2�W�0@{q��t���n�$��=�~Yێ�f����Hv	�fŰ8j뿕��4CCݐ2|I��m����H�U�
v<{��E��#X��y�)^�	����	�����%�N���űmw��L��*O�Р_�,�Br����0���>�2C	i�(u{f�K}�U�,�4�$�,M�Ǣ���0�7��
���|�Fŀ�71�G�>���DG�_���A��8԰�I!/d���)�O�]��D�ݤ��\��Sܲ���{U3l- [ֳ�?VG��Y:�7����<|膓;lJ9-K-���a ,L�~ w5�o��q�@���]�,(�J���	�r��*�(�Xw����E�gM�A;<��Q�˩�(a���!���`!�v�s�=�Ts���F�FrB��7�s�$y��tŤ�i;�UG������B|j��9@�Q
�S1��(��b^�p6�p@k�frז���5644%!�F��݅��B�&�L,����?2�:ӽ�4Al�L�5+�pf����m�򥪂����m����u=��;4�7�%G@Y
�!�E�X�t��ٙ�s�X�#���w�� C�$E,d�*h����>��C ?��(�����X��H�6��<���%Ј�	Y ��©Rt��&}||{E�0��@���wJ�߰B�F��c!Fi�<*mt������:������?��A�b�g��vNz@�Q!ќ9��mB��!+j�|-��PH��75tHֺC&��-=hCd� �y���$�̶��.�G+4�'�N����@����#o��p6�ʠ޼�%@Йy �0�$3|��gJ��
	$�BÇz��oj��]���@�Vg 6kP��	6���
*p���y{_}B	�9y�Ԥ*<o����rs4ub�M��}E�஺������e"j{oK�n��h;�8U���x�?�`�OH��іd�Gd3����W���FR��Μ��,i���Ui�,�v�O6��0c��rH���R�
Q�B�贆���4��%$m�/$�C������zz�/]�:��QJ/�#3�]a������Nį��r��B �1j�������p����ڢ-l���	׻T.��'��mɟ���X	�/�B���,��෹��3�׋U��^|=����Z�GE� ������&���A�u�-��
��d^Lc��&;}�E�oғ���i-a�z1���~5 z�Px�F����b���-=U.�sk�[��M=0`��u�ʽQ�y\<W�<V����^���lv.�t���,�G��/��bjј��W`r�6�G��NH��ilE���g.=�.�Q��#��2������d=p8����� ���F��`?V�v�z?�1�W'�j��J*S�aR�}Ԣ,Y��`�a"���ǣ�y�9���MwhӮj�9���D�	��>�#����.J;O"Hi����k�B��3�|�P��ۯ�ی2�ս(�Y;���҉}�L�'V��XB\�`[�*6��K�t^������ �����V������z��% �SC��V�t��^P)+!Ō7��\��<q��`g�l��c|3Vs�<��c���"n2Oψ��8\LL}$L��N�xE�0�oE��T�KŎc��C����5��'�oS��K!�8����T�yo�q�HOh�y� g���Q�6�����.
KN'`%hQ��#���Pa�B���cD�����u�Q㕞Z3�@��R��|V���n|��x� �����E�F��+ܷN��^���}�,���q%^�t��u�]��W����'Щ_ �*3�׾AϢ@�Z�G:��8����������9�g�K+ �ͺ��G��*@9��QX�iI_tC&�6�U�{�M�	��V���/���*�Wc�mq�5�6�sn�HP�A��[VO0�i����o ��G~��E���̕jH;;o�h��V��[E�S��`{?��$�hⳚJ�ɮ���c=Ec�`�����Y�Y5��#7�h��"/^��q��a�iy�B%"��ʟ�d��F�x��0�M�} ?��[����T� �a~�Wb�=�堢���Ǯ�2VyD������8Ve��2�f�e�'Y���[q2 ��\�B���sAE:svX��P	��/����BS9�!(d7Z:p�HA���nf��6?5�L��ԗp�67��]Ū/�����������#3s��e�B7"�
��v5|��W�)�<��s�����.�g�I��6]~<�����@Q�֟�Ai7�R��݂�N���g8S��nRs���Gr�D�E��A5�?��Ō`'[�Srv{�(�n�orm^��!�`ZA��4��Fc�V��ij$�:l��-�1�M]Z`푂�F.��!���y���N 1������,r���_��EL�ߎ�4�[������Ѧ�-�;��doGu��#�
5�����܁��*�Xb��S��$;��?/�b�{�Y��t����E��_sX��B�Z��T���ˆHSl�Tv���i����s1M��޾YL����W:B�%�]��$��ᕎ'j��`ʭʉ�*�5i8��o�>F6*��QV�a�f�Pۗ(�L���m{� ^
u���/��ϻ�9�T�i&��bC�br���Ɂ�E�.Z8W��[c*�.M��h��9}G��!��p�[,{~'�����@�mv�M��(ba!w�@���55�}�����y��/=�K}��R~u���_�N��cyC&ș�wf{<Ga�ߍ�f��h�m��L����4�̭L:���M7�0)�E���M��
�M��Ip�bi���<퇐%<��y�~2�7m�/�[����p��:f���-��0�=��� ��Ә��6�h@�`���ć77�a�Z~1}�iϜ�Z0=�d$�h�`��%����������ٝ�
1�jB"a�B�%B����y./`MpA�c�OP�F(���.���x��Vn϶�i��3�R�-���U0�yV0kSۣ�K�z����0x/{{�i�IA�t?��}3�0e�h�n�h��ns���b*�~=���%���%u$�� �K��<P�)"�t�2
����F��V�Vy��KV���Y�Im4�� �~y'���U*�e��e�*M־IL��	��ßcH؛n��4��]�����'(ID�􃽷� ?�����q�L�����5�P����n�X�K�>e���z/c�H��(i���Pk~N�X�)=��V `0�%���5�fX�Y~VB�L�Y�~�t����e�q���;��glJ�9s�h�����y!���]���J)��?!�o�&\E��!����&Xw8y���#Vrj#��ޫ���*����JI>~��"����0?JGH�èjX����Y�8ԛ��_��¿���,�k޼�fS4)�/j�f��6�+���]����c��o���q;l\����^$��'C�G,����8R
��d���T}�k�lG��w���
��rS�ُ�sb��CĬ�;C{��l���cc�IC��z�u�е��a��E�U^���1��B�Zh��7�+K^XHf�}�d8�֏�Z_$׌�#y��X���&�6h�Px���,����5L�Tt�W�q���R�����)�l��9g*U2HN��=B
����~Q0w)�:u��:��wd(˚��7�ǻe�x `�b�]�,�2\XXʘ0��u�v��P�f��6	���)�������@�w4���2�:F�^���9���d�*�jm��d�d�P�zr�#������3���W�.��I��j�;m{��+���������]iu��L�48��RQZ_�v`\_����l�ab�V��ɦ�2G�~��i���t���5Q�`^)��\�uQ�����S����1��T�7��@��#�]N�U��R���G#HB�J�6���\ug�4�#I]ZM�E,W,v[{vB��t��o'z�Z�"�qt�j7 g��P��Y�I��xT�������;�[%	�,�9�%b�+�q��$f��)�����x�=_&��[��^��I[�h	.����2������5��0C!|O��~�>�Kj+�h��'��F�ӭTH�8[iُ��0���j�4��[Q�ӟB�n�H��r����c|t����Bw�
J eg����,@��*}�~��7�eL�X��X��~�)җ#�FP���Q����<��:��O\E�6)���zh�����Y��V�����e ��T�O7���j�R��F�#�-W�ۓ	�J�x�~�gݢҹza%0邛m�W8)i&X3�{-o�.)�X�}2�h����j�y.)����vZ�I���6UJb��[v�G�OW���]5��}v3�#I��'��޽hӀ�<�46��Ub�� u��s���{{&��-�������g�6�@K
�	KW��dA��I���5X�����]M�4t�Lz_%�Ѽ���_WQ#P[ Ū/�1�j�=�rt���id%�TȦ/�%m�l�|�H�TP��BJ�}]aR�*�Tr�X��ͮ�<��^6P:��"")ʆ[�N=�~�)��"��U��?��~3?r��+�Z�e'�O�K���r�����Ka|Zj���S�a2BÙcː�2���%D���K�ð���:WM���ͮWۦ����3-�]�x(��g���}G��fJ����ȭ��a�Si�� �o�`O+rƬ��S���M�3�y 	$�7��cƾU���'D���fQE��T��`-dDIe��^���a2D�:؈|]�-Y*�bA�I�O>���zYNc-�J�E�%�Ex=�H����S7!�)��ݿ��}By��1�K����c�}�^y��<��$,��=3�ܦ�~W��@�x������|2gz��F>��ǚ�m��P���L��xܣ!]LuL�W��{��Ejs?5�
5F+��'�r�w��Pצ����/
�+"�^����뮑z��ub+���!�X��h�����`ݖdjN˷����X��-&�I5u���̪��W���.Ш�#�Gw��TO�3��]��Dsֲ]�z���Y	�e�s䣗���Ӊz��ۂ���5�Oj{*��/e�D�w�=��&����^��-�J�+o���>��������HDf��}����ўzS��A�'b:�>\\ь/m�0�,���^�~�Z�F�O�dnH +��C=�6�B�$��R�0��vˈ��o�{M�(��ѭ����T��_�+Y�Ma�(D����2NV��:5�P���+�!gS��`�,f�|y��Y�D���оI#>���l؍n��v�`�*5���f���T�5������ͯF�7F��b��i�;I ;���Oѐ�}rP�
�����x�������Ɨ���K����w�гO!���Xs;`�����#[�p��◞�-� E��M'�����ə1k���g�*ql#�c]g �����k?-�B2��
��s�<����[�~DrB�����C��2 j�iQF���O��qe�?��@��+��kf����!Ϛ8�#Me��^�Ó�jJ<s��3|�hH�n�3��t�Zi��<q�E(M��h߅�:�D8;^o�ŤL ����^]%�s�G��q�����P���ș����㌥� %���40�%?���O~F���)&Rm����Qqk��p:fk���MfƦ==��x�����>��Zc�VR�*�υ=��]�%�P��w�\�Ӏ4ӊ��ҝV�:Bª���H8Jc,�Y���:n�5��>���p/�}�
��6�=��ݐ��.w�����(���<&����ȫ�MzZ�ϥ�10`����0]?��j�$����YC��]Xd@C�k�[�@LɊ8Q��֟X�MQR(.�o���7{��ߍ��5���U�f屳��D�J�����W�0t9�1���|Jd,��	�-R��Kl��;x[�N�L{r�l�]������@V�'���u�����rUR�VS	�	 <b�`I���&��4R����9�}�MA��r�ks5DG��o����s���Մt不| ����:MҮc
�@F����}�����DxXR�g���O-�:�1Qg�_��PM*IZ�! ��P�ef�K���ڰī$1'��*[�S`�Eg$q3u���5��I�EUե�.����|t�ӣ-`�.*��1y�3���D%.���?��%��{(@GH��q𴮁�*�;V�\����Dq�����2�ᤡ�l^_����6'�W�|����Q����`!h�hp(#9�o4���.p��u�O�Cg��F����	~����;�W�"��v��8�<6]�	�7�}˿(��@h 4��˜�<�!TOnN{�}A����p���ǧ�����DE&SZ�[B���sz`
��}~p���]q�����2�׭L����a|����q�W�f��1F��`��-`���ff�M~L�۷Dpj?��^�r�����!���W?ٚ��ׂ	@��eC'Y���F�,�v��+<�֙�̵r���x^�~&T�
R��V̉��܁�t<��<���}�'�4�T�L=���&k�Yv%zv՛Q�ן�)�P���H�v�o~@�LN�ez/?��$ű�I%$
��\����q�g���i���+��X7گa�}K!���n>.4���rG���Y�G�F|+�b��I��-� ������-��纱˫�zЋ���ʹk�4�
kbf�p��m��Dn�����Y�oAL�o�_�#d2��Ͳ�}�aM�WGɹJ]*�TK��j�b�{�i���.�r��A$UZÂT��#V����s6�ۓ�p���Ͽ�|I�R�7F�󙃠��(|Z/�5��l�q�_�0�(��$�Urr�[�[�0���W�W.OGHl��e�b��4L6g�ǲ�@\e%����eΒs�-�G�~���4�v(�-l�����q9'�ό-$Q�)�� �.I��|�X�?��s��^�ׂW;֩�b�׈G-��ҦL�.�h�<?��]a|`�W��E�K�ɡ%�Q$�̱�V�9�;d���_\����v%�X�Q�V�߾���*f���,����TЂ\�i��+Q)-VD�P���^�Mw��
7
b�2vo?��欔���	�{�嵃��.������_�~���U�n˃�,���HIa�F;7���5���jj����`�jVRv��p�i��]�����Vo�oя��ig�sY�ժxw�Ad-�xz&a_�ߪ3�J��[t�tn,By܃R+.��?�{�H���[�u�6H7�@n���R.��9�K�h(~d��?��z��ڣ����� �b�J�dD���QK���޺Ѻ��5�0PD�L�F΂��`)�QU��)'�uHv�#A����C�q֗5����rx���-�腬����.q�}YI�:���Ս�-	C�FdH?���g���[IYV��z!0��K_�*F:4�]`~+'2��ۜ��EKix�B�U��t'.��aR��_�|�~c�S�����Y�,�� ������C�&�DxIy E���{���B���0txXx�Q8���E�P~!��`��'��_���g��2���|�Iq�@�sϯw>Jz]�ݗ�孾�T�6Ά|I���*(���:��lK-��K��!�$��L�_����6G{Uuw��cћޛ�;�Y����r-r��x3�k���e��c�Bf��|�a�_��G��c�a�����;F��I��$Y�@�����u)�z��I{�qKR�}�K���^�Isƹ�_��>�-+�;��7:�q����*��Ҩq�n�,ӿ9��r���/J�+�M�ϲP�e5�F7h��4�I����	2��D߮��˅���O��4������-���Y�C���A��w��{n���&������7���P�E�]R��&e>��	�y�GoZ{�T`�P�jL���+���K��ċ����Dgtǯ�U�ɕTQ����ɯL���Z�n��Mdv��E�<�*%Q��ynm���$�з����q��R]���0~��M)~"nn!_�v��v叮�*��9�������&5m�ߛL�z���~�"�>���ez���`��R�˽��_���Շ�
�m�P��s����Щ�S�|�	���QI�y��3���Nl���!3�ǝ<�
Q�����ѳ@D�!Sz��YT�Q��� @�"�m��
����(��l�I�4@N\������Y��yi&�=�� "P�3�t�����E��tDȿ�eđ��~�C��9&o�B�L����*X�X�ԴXY��ᳫOV�BD����^$��7_�Q��Y*<�t�t��	�B �@����~�ۄR�5�N��3y��� ��&�j��}�åty�鈅;y��TmU7}�QD{_� 
RݑE�i�w	�S��4�a#�m�X�&��c����,�Y�ů`������d\��u�'�b���2���A��جbQ�������B��Y�-n�kVD{Hw�j��ˤ`�O��[*$ %�m�*�I?�[t{�E�������9�h�<R�
�����_�֊8m�QT���"fcұ{!ydyqu�'W`:���iW�v��
V#�w�6�FΠ�%���V>�\^g@�QL��#�u^Y�H@47�g?����F��\6BC`�����0'��dkiv5��p�h�0��IcXf��gk���|��$�:K.����?�Y���蟃���UV�8y$ߋ�ݵ
)���7���R�I9L듷�ylğ��qVH��YD/=���\v����� LK}�1z�_�S��}o]��\B��s��Er�Fb���+1!
-�vb�J��EG(וC��W�+G���i�%WEp��c܀OT)��&H38o�Ὁ'�q�f}^#铰��+����;�*�_�U���ed�I�uZXP�Y{'�ج]�Ȭ���)�i	Ɣ����9Ǯ��~|j��d�	������(&�[S_�*?��^P� 
����PTF�A$$�t,&6�r2����7�Lk�`'(�7�%����� Z�|�g$u�O �S��pZ$�ڲ�6U���0cS�#���I�af��.����F�vL�G�NԈ[����j-C(�/�22s��T}���L�=���9�e���1 ;�8m���fU:�TZ���i�o�1�"t�����?3�D��Vכ�V>�8־��2��:�ql���9e^Due5az�H�W1��v�&g���U3C�^\O}oR^ږ�TBD�su�b!�F�ű<,Ǥhg��<s@ L����p����|s�:�#O�q�ۡ 0R���7J����1���u�t�6)϶:{�\�O�UvL����}�A�Xy�g�՛�i�U�|�U^�S4�e�Tu��R�o�៪��������5�"b
 4�R����ܡ�{~���Ս��˄3]o�Ϣ�	�[��)KC����P|[Qs�w@}d���h���Ĳ�{���B^Q���V�߄1~���h���i�`6��7�G� ��o7�=��V�!�!����sAbU��c"ʿ��nz�a-:k�W ~���$�~�T�a��Z�B�a�/��ںM�v%���A�&�l����A(3f�̭��R���{X����{�1FFI�Kq���޻����:�a�K".>D��M�A �a��Cx�2�ͩx�f_|�*���d�y�"�&F�+�r���0Sn�[��G��]X'j��?��,^�a����K�I�t&&�������nM�Fs�g�/�1���{�x؈��Z�p�T	��5U�,�F[�ӧ7�"�����s��-�x���3�����
$��5�Q���3d���c�f���i��7�VZ�Zy��y�`�:lع��xPB>�Zwh�r�*n�"�<����R�Y��d����Z�K�6
ɜ �����B�mSOuy�>��Ayu ����>K��[2+�c�������U"��o/֦�>2�� 8/�U�wg(Jy��,����Q������Fۄ���vn���W?��H�Ɇ!�ߙâ���r�|�����ʮ�)8�vS{��q*x	����df#t01�Ȓ��zXb<�[��睶�#>-s �H FN��Q)k�,�NH���IOo�ʾ�|� ��o�(p�N�{Tӕ.��m$��A��Q� nn�#]@�o
�-�(�A���� ]d.�@cH~����F6��ڍ"��zj��Y���������p9���V.r|�?-⚧�	
u�AKYA󷓸K��2�_�m����F��sq���d����bj�����wm~�ÖjQ��	`������^�W ��T;��{�Hs��vbH�F�b�;�m�}2eϢ]S����E����#�m4��q�3.o��7�~����hv]^�.U�J�K�=��!�K��#֢3��y�����`RN���\�A8�O�c0Ǫ���js%�kaL�y��Ѐ�9�4��ة��3<+!�_�j�,FXQ�h}��i��N��?N�t�*��K˺w��SδM���&���{O	���2�I`�	!ڱ�M�ɾCMy�/'>ٶ����%Ӡ}�P��~��in�<6�ݺb������[�
�����Y��|��Ӭ���L�2Ẩ ��\���ݬf�LEfT���`�m:�O]H�A\�{�%R���� 8�=taag���E`�Y��h���Q=���F��b���s���ҩ8�U�R}�g�(��C���&��ն}�L&Isj�Ehpc6 �GE�s���j��2B��_�����@A��XX&X��K�#Y�m;o UT�N(��<����Hu�/ �m�Ȇ%#��$�]�~%�*4-��^ۀs�F��`��h3ƒ��|�' ��*�(�m�C���W�6�[7A��i�XLs9vg����B��;�:�J�^���1c�ÜG��<���:����z��70k��?��W�b�o3���d%W�!XR;����,�"�"�s���D�6���o�-;/���������>.&'�����r�)��d�O�s1WG��~��7!;P�����.��[Џ��Ceg_�Ɍ7�I*&$��s�N�`۶�&A7aTv߬���?��1�n?x�{�t��?�F^���~�:���l��	;#�����i��fj����?�t`�S�Zy��z��=��鑠�d�〮�-��Ȧ��꿓1���$r��Vk�V&�����+f	��(c?�/�F������$�@�OnY����	��H{7N�V�B/Ds9���.�� �>˨��G4Yk[����gb���-�Oa��g�@�L�Ar�bM�Kٮ(]���G���R�ON������Ƙ��>0$�
^ �s���t$OhX�,���+�O�u�Fι7"�i��=t�F��˳�Zo|�#���s�x�u-���@�.����z�]��y!��.Wn�q�Ǭ�����`�v�F�ќ������2��7}�DZ� ��MAV:Yr1��,��Lo��g3���D���Q<�9qTp	*�7'��N���6[�2��H�h�'v�i���\J��"�?��j�$�����E;7w#$��GI K%u��}��17��F�;��SA�^�����Ḍ7|�h»�lK
��8�o:�Y�+�)��@�g��O�t��LI��_q��p�O(�Yڪ�_�Q��B�.J� `���0�Z_���훇ezG��u\J�z+���`5t�j�2@��_wKM�V1ݨt����|���_Z���Ć�2����9NK�1J�Eu^�5�H���H�CU-�zGqU1�RzY�j�G��>�>���z�$ئ�h���v^��d>�h̠Uk!�L'�(W�Y2�S�����$��ax��uz9�n����n̚Բ�C��Y�����N?�ZR@�v�q��u�J$�ڟ&�o�:��<� �̂�ƞ��B�)��A����h�S�P��>}T*p���ӧ�����Ĝ#���s�_X�\��	�u��зg���d��jM8��sl��47n	�lXa�_#�N�����
i��� ���~(\=�"�/�^X9p����R/��g��!\���&Sض�&xR��JY|KtҦ������c#B1彩chäu�HO	�Ad':�^�1R'�]�U\̲�� ���C-#0!�E~K�6�BF�|I��{���D<����аʂ�!;d:�L�.y�y�X�z�U���Yu�i#_a0�M�u^�ː�D����� B��v�L���4�:t<�U���3k�U��J��Nu�Rj��
�p��p��(w�*g��^~bJ�M1���W�*b��++��_ޝ��|7C_|ca%�Z+�A���D� <BФ���T��U�B�=e�u�A�?�Mհ��N���܉#7'|���][HՑgo�GQ҈�hw��\|��ò�R�/��a��%|������]�.A�:��'��<��:ʪ��G�*�c
��2�g��e�&�l����A(g=�ٱ^���ϴcs�r�l>�U��lt��U�Tjm}^�Ʃ�;v�R�5���_ȭ`�>x�C1�w!õR,�h齈�U����Q|�[O���:���6[_�"�]e����PLԽ�Sˀݘ���%��c���6Y*��Z�c����*]�Xۣ��]Ut��޸K�ugm3�z/>�_�۽fc�ά��W��`����)9�;��^�#ѦNK��Y�6�Xg7������W[� �?t$-�.�頞�ɨ5B5%MZ���hH��T7�9Q�6/��~���*�a�f���y��d��P����)r���W��i�e4�D����c��^��[ѻ�C�r�F��} ����ҡD�Kz+]z�
mT'��;\r���=> td�����?�Tٟ�V���@�>㫒.]��z1��v�R���/��������Z0c���	���tx�=�����x+uY6���7�X���p�������G��A���ٰn��&�E�^����;��'���56��*���=�ޕR�^NE�G��Y�s�"]��~=��U��AIƪcC��э`����('�W�۫�j��!RF��;�o��r�_�onU7��V��8|��p�Q'���;���P��r�V	�b�<0��s�j!����_��wt���6u�&�S��{F��zmP�o�׫�'Ld�5��:������<XĊ��wJD��h*����e*Wz�Fy��q˰����!�`��I�K��~ �7u���Tk^@�J"*���'�Pf��~�.Ke��2�£��<��o��h��=ح�*��=��c�.)t�@���6;�ɟ�Ϭ�x�ѻ��lA��v��٤㺲�=ep�~���Ӄs=���o���2s-:i�u��ˍPP"��a? ��*cw�̱;����/�Շ�O�aD}ѿ��z٦�K�&���;��g+��Sz��ж,����Rψ)pf7��Aӊ��>������z%L����h}�Đn4h@���٩N��<�^��@�0�񈹣I��Q�U�\���R8ʬ�6�#K��W~"2N����������?[1�֔�4�SZ�.I[C*���b�ē��KLe��Ճg*��h��P�z��jZd���,L5Ḱ��G,��?PѤ��ݡL-_hvQq�V�l�
M�e+C�}� z|/@�M�:3[�ßx�V��}�`����Z�{sBJ�R��!���
����]T�%fb�f���y؊��ʵ�9�AL���!i0dJ�^9�!��$Ha�'݂�����m&1Zt�zN�!���>��C��1����ޜÚ�iI��VH���FK�u��,��r��(W,!ͨn��N���V�#d_b5w�so[!ƾb3{U�ʍ�Uٹc%��X�2)2Ήg������96�d��n��Ѝk�M+yi�6�<	�a�0M�,�%M�Y�<�r���f��\�n���ķ̥��<`m4)����g&M���v>�L��\��ϥԾ�W�9�E��a��b�Y{������0
���D�vE=O�E׆-p��{�dRs����+���אk�g�V$��1s� ��(��jp�@V	8O�~-'mT�u∋3�gy>��ʛ��+G�Y��3�|�Y
G�:��]mP�/�D��؞s!s��&�����+~<�Ré�E��y�����p�A���:r�lǻ�@l�.M�����}1Q���zy �Q퐺��:u������_G:u���f��@���5��0-�Y�y<��O��J�I��#Z��h�W`p"Q��_���[��Y�`��w8�!$#�^p���?�HDB�=|�0�������9��hUq9��J�Ѯ��Cʶ*0���Hb���u�P[d�i��/a��=�\�f����_[	���"��`v� /҂�v��s��Iުׯ3����S���&�����}�F*嵌�����E[(���@�_6�fH�'��_��&�GH��W<����Aְ(Y�m|�*Ѩ�Lg����e��Ϥ10��<�={�¨H�r�Cy�{����N�g��.��C"���"2��C�E��4.��
���"^�3��q�����	��E����H�Yl�i�ѸR�e�\���Ɩ�ǵ ^�����$
 MY}�մ��##�v�g vѓ���HW��0Tjq�jz�D��ٚ�;��f��	��8�m�ɇ�١XJ{�SAX����\�=�A���׌��pu�� �Y:�^@����e�tp�K�Ŭ;i�}D�ٟ�R��*��O�y�ܥ~΅�8��ap�Z�K���u�%��UP����M��������9ԋ_��wۡ[�=^�d�S�̀��H\�8�-��������խ&?�΀%�n$�#�w���|�,���b�d��\ߍ�1���sP�D���a���:�_� I`�Ŕ���'�h�?���»V���V�4FMȬ&y��e��h4-�/I� z��=�_A�BV��H���և��n(��i������د���A��"]h0<��5'Z�W4�l�W���ś�	�(�	"����6B�ut�Yp1)��_<�=Ju��]F�u�E�]�1��M���*����)�Rވ�:<�}�h���B��?��]���+�Kٱ��d�Y��_`ǀ��6��-��u��&��>��-an+
)*�H�[δ�Μ�2HAi`��ʡ���B��˯�	i�q�0��=.�s.�Qȱ��:?x BF��I�]F���8]���yU�s�^��7��E:ng*
�-"��J��ε�C��������=0��8f� �q."{�<��G�-	|���H�����OX#��]���9�sr�!O2U�BA���Nc��������29d�I��{���b�}��F�̈_�:��I�{��m1+��-��{NPJ��8�3�h�����[c��㞣��-�0���j�x���o�T�qT��A�}ҰA3h�9��^��F)�Q1�42�D�����0�+�
X�����m�0>�\�ea]�D]�&�Ɔt�6ezr����_9����'!�dz����!rϨ7��y2%ӌ=X:������n�(�~�4�a��uP݇�m�����c���5Bk?��o�9�
�)h|*�MS��>n��9]|���( 8���odc����䭡2�U�U<*G���h�+=�ȎePezs_�uP�������;#�T�C��Q R�5��be<�����a�Y���.��e���2����mZ����K�j!YM�|�؉˼/��9Zx�(�Q����fi]�'��ʪ�苕������4tO(���8������k�0�(�@�op_�X&4Px��z��%�׻+F��IV��+.�F��#Ӓ<Sb��Ϧ�&o"�\��Db�m�17-~�z�b�t����Oz�;v��)큸����bl�9HOq���a�#8�h�qD�������8��׾;�{���T��%,�vI��/D��I�h
��C�����3�qn�0�nC%u~L��ʮr�U#>p��)I		v����g��B@>��&�:�j��S�O������T@� W7�����Ɗʬ'NwSY�*{fCM�e{�%�L	�4�i�M"�����{�ъ�ƅ��� r�x�/�ly$L��z����G C�T,�1�ly�HhΨ�A�UQ��X��[���3\���?��v[gew�3^	z����󝎪�e�K@b�+v�3�)��yCa�K�l�Ch�>;�|@�k��t�����Czg��_��O4���ϥ�e���!��׶jf�2Q��<��W-����|����$q8��f]��VP�gX.��V�X���	'=��r�  R���Bo�/���hp�~n��oIX�bN��0w��\�j���͸0��j8|!�a���r3�1�D��~c��U�k~aհ���X�S�8� W�*Q�{R�����ڡ�;,��hHCH���C�̏�\�Vي;�9L�}�tc���+�*	�+����'�}8�ѻ���@��8�y����}/W#�|�T���H
Q+��33�kX�͠��W��M/��Ŕ�R�6]�V��:���4��Hǽ��
��HCǀ�[ӯ�u�<?��lye�^�'W���e|j7�@:�*<��ik�k(gY�7���h�ϡ`�G��A@�hGv�w�y�ܧ��O�wcV?U����.eEL�
�5]�@�vH�?$zk/;H�'37�o���������mq�W�0N��x��:ň���Z���������^�ʀ%{��ZR�Q'7��ꑐ�P(�-@�5��wZ�u2 2��g+O�]�����L�	ra����Km̓�ī9�%c	o�fc���[������˴��U$�GY�����J5�ǬK��a��Q/r�܀���mF�3t�dq�����3t�7�����(�yk.Q�}>Gc(gXb_�S&)�<�t�~��ۥ�)��ּ����!��G�Tj��B.����f� ���%�l�7j�,<�ǘs��8�v��+1C	U�קJ�gvY���C%�[w0�Fb�������F��SD�_u��|nE6M����E�2��6u������ 
�j8�4P'(���?����&S��s�,z�����ƞ*��c]�-e��:�b�G#��;t�Ҥ*o|��;Ā4uZ����ǰcx]�+�b �`f:�vd����2b�Ox�V����0j3᝷���4��KMrQ��[kR�٘Me�J��\� 3/v�-�B
C�j><�����rF��T����Q�|�V�D�8�����:���&�ö2Z|�����a[ �q�� ���4�r�ƕ�Z�h+{c����g��{�:eWF�Ь��w�*�$�oE�ٟ5��C∋��"��w
��	��VPcB�Cr�K{�c��D]�Ϙ�S���[��sI$q3|��J�F��໖qI��Ӂ�=t0��`�,��بޤ���2k�c �ɱ���Hﻺj���4��[�(-;}���yV͊��6�;�J=Î�v�\����Q:J��K�ߣ
���Vn����%���{�$��22�Ө��t��z葾o��ٝO OmF���9�4 )��oxgr��`98J�����ad�1�?������}���Y�CE��	�