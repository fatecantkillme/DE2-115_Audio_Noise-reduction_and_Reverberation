��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<��h����Bo��}�F&|�!��5��'*�oܒ�8b��@�������O�ʌ��6,3p�Nd&ץ@�C`f޼&�����O����2Y84���?ŷ�D��RS������)����8�ά��e�VԪ%��,��5"%mG�+�sA������ԞMkԉ�EU�Z��:��e�$�k�@%��G���掿�N���_��~��2��'H��E����!�����cLfk_�|�n�<{AJ�*��?�:���[��j!���n�]v�ϼ*��k��0~�o��D���� d���)c��	�l�Ž+1��oD�7�g��Zp|�;�(e)z�ObLN�La��+a`�u�*��/�sO�1��%��c8J]q0�����q��S�i�b���{�Z̪�+�I$-��' ���Ce���!���-��,�g���f����%m˖ȋ߀���Ta��Z�;3�I�����i�_�ޘ!���y���z�f�����"�:��^m�v>J�8�=YXnu8.�����b4�'��E���Aռ�V���.�W���In����ds&NL��-w��_J�ᬊ�j<�ބ%�ِ��7�d�'�I�B�+����Ņ���$N������@�y��{TߍQ g��X����+��Lh-NR"�D�����M[�f
ѵd Y]8��������mӸ"��M��8'�b��ē�A����yd@�̍ё�Qo�����}�X�����C?�Dxyx��l(\I&j�/$������vOfl�q^�f����o��i�<�c�h��/�Vb���������"�!f�vb��Rv��eEfҌ�	i���w2n�ya�T���V3�X]@�W�d�Tݵ?r���D5�~���Q	a?�r�Pj}��;R/��3�((5���&�΂Mϱa��c̔S�` Z�����yx������?S��h��o�� �8+� ��E��U:�'$.2FJ�[�!ĕ ���u��rP޻c#���8/�ܓG�t�C�h�["��V�QK(`ע lЩ2�?��8RHBE<?�c0M��N?�ʫ��Z�,��*QP�����8����y,�����`N�G1@8��}	�,�a�'I��_u��]�i�?�P/�y��T���h�A13NL1%�\�"��S�RF#����͐>�7�x�/�����(�r�u��#����Zɱl��� %��x5}\k�T�Ѫ"���Z)R�QM�S�8s� ��N��<Ô�4���C����vɷzHID��n�=)�[Q"~����d`��}��a��iu#t�r��"k�>�ϊ�=��w��	K�pﷵK!�/��=2b���ml@�W��A�k+�b6����굄�3�3X�_��i�Ja��t�Ya��	ԽV*�_�\b%�}���0� #�X�EUew�c�ЯT��zs	'�9�\�O%����;�+����d&q�R"�I!9Vwx x�>WCX%�xᇡ�m�"5�aT�l���Dl[ ��Č9�T���{�6Iw��X��ኈ��� B�7K�)sc�Ԣ�`i�w֏�	��h����X(yw�]�������H��b�s3�W�,B=�o-�+&R��j
�_RMr�bn<̚9B�x葙��%ˆcL��xE桻�?G���&�(,��[���푱/�����Z�&�l劊�����WsU��K�'�~�h���#͍w�7 �Fsm��c���Ql�:��A�� ��0#���x1�qf� u�.�g�y�S�C9|C&U6�O�7.�ީ�Yp%�(��I&	�z,I �`=���@e�Wi�.{��%<���C �O
�$�m�y?
�n#B~s7���Ƶ�����D��+C0�`5!o�*�YR��
����\�y�	�}�@�g���X��O[Hd<��퉾j�i/5U�����Q2;�8���g�8�AM2lx����,+�o����,l�Iy�%��r���r<����,<��O��YeZ�F)\Ou���� J,�����U୥'B����dl�u�#h��^jqz[jCK{�*�!RG�0�؁,���ZK�h�%�>_��(�K���r�P{�{�(������Z\�މ(+YT���"d�lQzLܕ�Y��`�Pup^E���`�>r#D>���`�]�|�@)�n�&�_��X���~6Y��>�>��R�����R�Tj ��D��H�k{�ƚ�����TF�E	$�{7�5i�G�
��y*_��]���G��
���ﾴ��54=OW;nt������^#8K���O�~E����g�w1�kY�,�b	�L�?ɉ(XP��Y�	:EN��@"b\nuP.e@%QX��p�J��L�+3��S�l�5�-9/��U��a��@����6����ߋO���aHOxi�?O�wi7�έ��NN�1\)Q��h/h'�y�q�����n�jӬ8�0��r�����2oe��3��^u�u���e�����P�H$���H�_����x���d��������.oA��?�ԃL��Fx::�t���ftT��oY�Vޤ����np��JM�=bqn4ƚ���N%:s�1\t<���P��� ���{��WD�V����
�a�eDݓR�[^hSr��+�*������gG�b�j����E��G정�^G8&��;Je��� ҡ+�,�c�
������-c�V]�x}T�6v�w%�� x0-�����8�����v�*׆_��:��Y��/�>������V�O�㾤��L�, �FE+w�ș����Τ˛����@�D�kOD3"�KM~�]���f|$�نf/z�(�en�����>�EV�I:_mBE0���2�B�A����ҢozQ�,W��Q�v�į;H�k���I�tU�-���q�%~�Eb��U״�t�:^�V�͝�W���ۧy)�(\8f5륉����.A����z��ÌD���ϐ�G��������~�����/y@�y�����no��u ?Ş�V8�;�xq(�l���`8���(FCe�AR;x��6?<ށa̽���є5���1�'�'A���)�6cܒ��u�Gh���6�;x.|�b{�<�lLϳ�"ډ�׃������3M2s ���#� F[���HF�p�h);&�6��G����e���\��>�c�v�ۺ3j�����e\%uzjS<��V__�!km@��B��i�*�7�ߴ����Ը������b���G���a��,��5f�-4\ �:ȝ͌e�)Y�>�����O)�v����-6��fp��[��b�r�Ⱥ����]sr��t�ݞ�׃V�yr������m��2�ʔ-Zj�b|G���`R嘧�x-n�+���P\�bNd!T@��{������熔��&���k�!���LL�8��R��2m�ji��`V�<��O�8�L�ȢBN��PV��:<�K,P��J#���������G|��hZ�����i��ފ�P� ��+'��CF�S�u����a�<ݼ��!!�wˈ���J����u�"���9*�6w��.F�\.�:��"�2�?[:OkeȰ�K��_:�)k�H���N��gB�����Etsr��G�j�J�Q�:�΋��ڂ��u���0js��Q�2O����g4ѫ���哅)�����k�t�}�t�h�6�:�h�tlo�6�`|U�e��+��I�@$��tH/�~��T��Oah	5�c�Pd�IƑE�1�R�~��%�X}���{���f��~n!���=�EqC�`D�/qP7�ӵ����A.��>I���ʂ(�}��>-�Ч[�Q���|�d���ƢH�{�_�J�����7�Za����+1��傚�y��IG��l<hk�a9y�m�r�Om:i~N��z�RԂ�V	h������|üh�{@������7̒�%��#�{#�A�=���?�<�ƭy�R���땫O��#<c�Y����Z�+q�M�!������/��:^ǋPG�wQN��N�A4w����1WM�k�/�V*m�*��f�K9�&Rk�y����z0I���e����iT	�m�x���h�5Utt p���|�;Z#�-W8�s^G�s�7�[��ǝ����-U��Ô�L��R�������%�-�}w8d��L�
\�UJ������y�%W� ���)"��Oµ笋��q�oQ�K�Ba>WI�]sĆ�g�0�� A%F�\�lU$�D��03&�ϖ��M��!������8/6� ��/�4ᅽ�M��u�-x�[949��Rhy���ͷ�=�ݱ(/Hc�1�1X�\���X�@�о��R��M��+ꅧ(3lHS&4l��1Q�QK�Y�޲�>j��_�W��a#�<�b�P3��'��KIhHW`��K��"]E\�AI=ePK�|�Ph����(��ƅ��B ��Dl�-'6i7�2��8�=�`;XX*�o.cJ�m(-^6�.�D��	�·n�s5n���} ]�p�j4���	Syj�W��C�􆏁�?F��%��꥕��t�Sf���Ɋ��R:���.��1��1��u�<wy�ύ;��
 �2VꏮB�Ǔ� L B7so��;6F��X��0��ʦ@��t�5�x��9Ѩ��K[i�D+ A7pӷn&�;�V�}�*�8���Y&�O�����Y�K��
���l0�H*'"��� 97���P�f��ՠ����@=y�������BC\۹qqg%���e5���ɐ�0��
�~=5�|��0RA�.޸w0*����ݑ����[a�k}�H,�:wl4�U��������������Hމ��0��bE���Am�4���dR5:8�l��c�W�R�P���G�y�wa�w�m�3����̟W�_TؕW
(0�N����V�wG�\�M�j�����;p��Wa?���S%S���:$C��>�e���^��6�*Յa�I�+{�{`�C=C:6���p��e]�4LQM����X��c59��������̼m�|a����������smQ�f%�"�%�z
6� �AC}��.b��.�0K�!�e��f�� 	?�+!1�Q�T*~3x�Wb0��3���`��u������m���U�g�U8H�E���`����H����<�{�{7c�n{���60�}!)�~�>6ʤ�x������O�"� Ha$�C�*iy�Cç%S�}�FPc�U�D���/уy�~����ưEZ;�WD���;+��W��ʣF�h�Z�8.7_3�k��mݒ��@J�&�X�֚��^�+�Aק4�l~/�J :+��;7~Mcg9��;�A�,s��-� ���̬���%PS����;Z�9n~����h}��ye��'&(�R��*V^�ϋo�"�W!��ȶ�V��b�?�<�n�΢�J�Z: �i�S��jr�u��}���T��l��n�u����Ό��*$�%!lm�e}1_� %�<[x���eF��*e�D�
�@E4�")a��T�b��Om7�UA�t�f8 A��4��
#��ޒ�8\N��bյ��öY4��.{��~@�QO5e91� %�c�+��U�d���V=��Տ������n� �ţz^g*éC��V/���#�"���X�U��FP1�F��.?�.��_o���V��������Rq$F����^�e��X`�4�fd`�P�dUH�(�^����G���B��3ܬ��W5��]��3�Ma��}S:A~ �]��f(k?57��$)��o�u�weoa���E,��^,~��v��[~F��X�}leۖ�n�<
힇�9�wL�\0#F��;�Q�io"�/e�Ө��{���	�.2M�e��j�칐����ؕ6��L'���H�Iړ˗�+��u���{��������un���Fv;�*�v�*Sa�����`v������ �jK%��W,�W�WQ0���ęi�+aC�H^P)z�&�G�W /�	���쨌5��RI�03�.fq�[�{r{��D�KPÜ��!z���{G�'J89��'B jn���%P��L�ʺ�(�%�C�70u��k����	��}-�{�y���m4_0U���45$L��l����:I33�^'5P�\�q	��&�|���[�m_r �|th�#*6�るJ���.#H2tfS�QE}�/ZЏ���W��j�F����[��N,]o�s�PR�_�p��@�`-juB^j �六�$�]pX�8�9rW����T��Ϣ����c���`aڅO��B�yX��H%�G�M��Y�;t��I�^�L�j��V�5x;��dVA���%���d�;���(Ž�`��7��)8fc���_�6i�9�yd����s�V
g��ҁ��^g��᜵�5�-������u|�C�R�*��N+���s���	��Ex)����#?]�y��3 ����ҫ,����6��Ō=�8n�5Ţp_uyO*��4;R�k|�%����vs�3?cd��4��P,�t���r:-�����1f���c1׎��K�p�4�Nf�*7p��9]�뀥��R���{
7i�A�&;�X@|蕶�n``�-��<�2�)�- ����'y�|8ROZV#�!������M�n��3G��96F���1S|W���"�~m��]���Ɣ�[�\��_2�3'������ή���P��~��@7��]�NY ��q�ah�_�Y>E����]O�ǢR�������K�P��@��%o�o��q*k���t�ѡ�1 ���B{bYԄK*�ƟT��d���į��`|O�hg��� ���^]��D\~o��"7p��ͱ�8n]�^ c'Ӊe��xM[��Y��u;3��f�/<{��9Cu.�m)�cLZ@: � [�\�������<|11X5�B$�ڙ�d����
��$!�_�%��o���!(9d����}^j���a��<퀒�ŝ!�BI�V���F#U�s/��ZvyM����
��@k��P����3I~���7Dj=jkVǐ�L�H,2��χu�q���X�Yb.��}M���qZ��gQ��rISv� Q��Fa��|��b����Ts�� Y)[�nxHn�z)@� a�x�CTC�8 4�Z���l:��U/8ma{���*C�fӢU\BI��٘4��q��y%Z��h���Qh%����Z|a�먴)��4"����GG�h۩��ZF�Ode�A4<4�Q`Ň]����������J�$.
�1�0�䞠�D#N��g��#�}�3���i:��x�|6�f����h�)��ڔ�O�)?=2 ˢ'��˩�FH�Qc}/~�M����Q�qk��;�R��A��d����(�X��8���N��ċJ읖��(n/�^�T���2���W��N���d���0SЙ
	� ��e���?�s�&��o^��y�����B��Ni�6-rI�)���(;K��
#��}%"P'�H���W�w7Ꙇѱ�B�����=��C.�BȽ���;I�m�F8�Ǧv�"��Sp�i��l*�F��t�ٹ �CR|c 1}CM|���TD;q�Hmc��|g!�Q�|*C�=1{���/�Z(t�ߝou9��gK�`���$_�X�5q�yX��U�*#.�tq>�y��Eh7ir&���
S��	����}g�rT�f�Ky����],���꽕"��Uû�?N�A$�u�0y�� 9�����B��r6������u]>7'T��cȱ��GgiR8�i�[�t�ή���3�ezh�B���<.��/�¢Z�"
87�|���y'�j8�*�=��?�E�R0�����;�2T�Q�{��~W��'K��5~1N��'R-�r��f�����8��m�cJ�����ڿ�(KC*�h�����I:� Y|�׾%���tZܦ���t}l�`"�>�n��<������.�V�V
�t���W��j��}�?��2d�L&�52r;5IY���Ė�Y1j�ו�q�"��/��OS���4��)%�9�nk�V��ÿ�n_+!�W6�X�������-��>��/�J��T-GT���æ$�:k�cz������A�^�{�E�T�W���X�s�$xhu��`Q#���w3�l�閪�KS�j]> K�8�k�9�`5gJXL�a�Ҹ�)\Q�
 4R�R)ݚ,v7��NE��BY)]��0h���<c�����I|�!+�>Р����)B %�|/4Q|?^mŖ��Lq��~O'�4�I�c�OIM�Nː� c-�R� \����bu�ȱ�f�&�>�Z&=�.Mw��mr��P��Nq�o1����V��p����o��i�sEA Wc�%o�4M5dV��g�4�M�4u,�9�C!��Z@N�W�H�)`r�)_|
�S��� p��jǷu�����;���F���g �������7�|F-�/}&8�^39;�K�D6����F{���r; ŋ�ܑ�����m%�W�Ҍ� �n�|���V�o^R�G��3�}���>��#���}B�FiF�9g�#
���O�o�K�x�R71��������^���=$�\�!��m���G
��\�fc���H����t2�l	J�cQ���"�d��CҎEuŅ�]+���F�ψ�6�#t��lihS�A]3�a#b�Y62j4�!>=/�! <we�F����m����7��JB�f>ר0�!Z�����)u��J���S���q?ׄ ��L��_��躼͸���O2p��;�f�	�}��*�$�")�Z�[��m�Op��}e�x���Cc4Ԙ`ZŶ�)��^��x)O�'�U,i�2�����
��`C�	�;�T^5�&$��Wxi�f�6�G^Ѭa�v�:���9��~����M�=��$����}ag"����X�#S�օ(�صK]���=�W���X��C���Z8ѷ{�R�k����`��4πCjx:PRV¯�{�z�K搃ɕ��W93��z�7���&��L[(�sB���N$�o��)j!4a����
m9aW
k�?7�T�X\��Ko�G<�W2�.�
��;DX��xQ<K~(P���=	+�Pϼ���©���+tS���s�Dz+&[/Xc�Zk9�c�T)�jSUґ�����A�3��z?�a�#�CO�(�t��H��n�Ł(�W]x=�[O���3�ڡ�!���ƨ���S�Es3n�VJ�U��r�ֻ�]�{{0	$�lᔪ
G�v�j�],8�p��,�p�~��
�zƜ{���"�Z�U��z[����O�o�*u�1�C�����v��YY�͖QY'=�q���v�����7w�z[~*�
97N���Y�|/5x��"Ɯpߏ$zO�7�GgÄ���>o35�˿�2k��Ii�\�tEZCov{��P���=|�a'#�����k_J&�;L�kz���k���T�T��I�R��ȹ	� �:BcB�ev�(&"�+�C���Ra�å"\3Mx�®��Z�VY�� .O�YsPHQe��Lᙄӷz������N3YJ������Sx�	�ѳ��N���[7A"p�ۛ��?�l��D^�8E��䢗1�!P5�J����4U��+Ѳ����&�o���@�`�ﴜ�s#��	�?z��=��2y(��#>oW����eh�|4�4�V�<*��
1������ B*g���q�9:ұ+d�JF�� ��d��'�F�)T!}���
����z"h�a칈�y�L�_��A��1��T1���!�c�-NLF;c1��S���a�X�4k�)?�2B�ZV�Y�]=�|G*m�⚾���aY�*��~�CD�dK�/���Ұ����u�Z,?D����W�m�}�+UAn�r��3����{7��"	�h-*l���������uQJ��@�G�S�+۶d��.��~�Y�Y1s7r%/d��*1c�2,��(�9.��f���F^�Kԝ���De ���w��҇;�ܒ����d8������D�5�?]�+��Ka����v]����^�8��C����ɬ�(V���*�e��/�h�H�gZ��"�������9�����92�����8�G�.�15_��Pj�`�{�xꋘ�Tp�(vX��9g�i����u�F�ϓp*K"�t�g���
�(6���\EG�}%\���s�c������""Ύ�N!�Z���̿r �%�8z��\[�'W�-r��}�t�|F]�pP�U�0��iG���N��M&�EuF�/�HS��S��-N��W����P��b���eo�*�:�`y��@�-��.�_`������u6_ΜB���9�LQ(���"p��y�mnH��	ԑ�Gc�PѪZIh�o�Z`S���ڌ.t�E&e�� -`h�vv�y����3�f�m0���@/Zf,�
���^[p:�����o�y�Y8��h0k��ґ�PLJ�k�d���4�V�j�f����s��&V	��Id�{b:���}BQ55%�B�c�ܚ�R$ ���t�U?���)�t�u�{2}0!�t��(|p⓭�{���6&J�5��dQG	ȑ��q�[�,���/��\QL�)o����ءR�=}�9�3Nw|��� ���ݺ���m��n��f>�h�����b,a�9�������BC��&�g��,�v�/ܡl�r���+����Pt��G��)�yXb�����>� �V�SlC�5��l]�)<G	G��D��E�B@$z�,��@o�4�{��yR�t� @��U�V��f9Rq@��Z�ga�~Y݀���+x��P�BU���)��xl��0��ѯ�r�J��,>����(ԁF����4y���5s~Q�o��	jf��u��*��9��8'1��d�F)��%�w�c��ǿ������$�i���iZ� 7��H����7�%#��\�9�I�L_ٺ��1����6�>�����J�&����"�WdRC�Y_D�ˆ�4�r�)�!�fv[�I=#9�\߂�Ga���̭�Y�]}ǩRDTd��3N��4��-���K��E��&�@�1�	��������-?�G�![�P;J赂���/��ŗ-9X�c$X���$��r�$�%�����=L;t��|�ğm�J0mH(1"@�7�HG�w�FG"����Sڷ���>%?
�k��e���_�Y��@;���-ɤ��Xo[G&O�})s���@!,����}a[�EL�;�0��igV0k����g���$e�UX�9>��H��ά����x�J����l�_��oE a)a��YXIX$L��������C��2湆�|}�t��}��Z��|���D�H!���£�<��� �rc�������	�7t:�yt>��#lup��~)��V�(�ծ�B��4��� l�V��S'vR�����G��]Y݋GE�Z�C|C���u\3K*3���xX����F�"�k?��t��u��A�|N�|Nƾ��*��d�`���x&����\����K���
C(�#X�a�J�qS7�V�Mcz�v��J���5����_�_���T�d����N���>�&{��qlƳ+�N��v8�T��_kȚ>92�jBwrt�$�A���ax,Fi�H+M)R^{��v���zVB��5x� �L��C&�Q{��h�O��ňwø�Z}<��I,�h6�P�-'�{d�jb��ܺ��?���.�%T ��Qs/�=�ʿ�Ժ��VC[�<6ͥ0�����]5�'�Bu��� Sn��r�H�}z�KRr!�i�՜q��6���0-��:<L�^a�D�K�}^؄�g��(Lˋ���h��(n�kn.r�֨|�2\���؛�#���H�)�ѹ�0�sAzf�7�y�N2.7����~�����	V�*m�K[#���4���p�Y�z�0�e���N�>�$Au�G ca]ɯ����h�X|��4�4�y>��x�,��X���Ub��}��;������V�6ig���|n����/D�7��bOW6�G���E�1D��<4�\�p2�4l����I���J)�a�y��ƒ'����km6��bprV�pAg8jxVCo�#+Zd�I���1 .+N(�.��K�B�������^���������bѪߩ���Ev�o�X��tq�u����AUC��#�|1���f�A�q�kg�H���� D��Q(=�s�� 6�� 3-��W����[N��:F�^]�;%_���[�H:��'�6 �S|t�s�0Fs���)�2�
��.j٢.(&zv��4ij�߈Ws"�]�cx�b���a��k7z+@�\8�鞂�|�in>�]�j��h��}��W��M3��'�;]z�j#2
8��������wgS(�i��-��Ӎ1�i!�}��z)/iN3Z�4�;�ڥ�_��f�'��ԯ4����R����o�@N�(����ۀ}MY�V��1�@En:�n~~X�^�6��s��襼�k�kth�L�#;�t�D7�T���Oj����g�ԝB�g�|ãt����)�$֛>�TT%R�rV��L4�~
����=��0�����jg�l�*�N�_n2�O�w�,N���Cѡ���窯���h�uM��Y�m@Wz>,x7�Re00�?��7�Ќ$�-OM̎tX9�nAG�)S��j�^�Y?q���<Ȗ[]��QS�po?uؘٰ�Y�J5��G3ua���Ҙ��C�Ad�JT����C�\�^���ߴtT2dK¾=��%]d ��U�[w6��� w,!}��T�Y���� LԬ`�{���]��.<�wV�h���#c�C����?��|.����F���I[��x$�IJ��8 �M/�G�r��!�8����;��Ca�S� }���3y�UR�f��>�)��+��\��5��hBP��*z�?l� ���fcօ��j���<K�o͒.@ɋ5��M�b����485�
�̖\���-�hm����zw������\s�_	d�_0Y�K��I��l�3�a��d����/���E�Oު�ŕZ]껏�φ���ZB܆�y�����jiK�V���"^7r�Lhr.��UC�fm;�4���(����S���#v%2{5��C|p���Gq��r��gdG�T�p3{"V\�@�ήh��oԔ�$����>	�,zd�� ���7�]�g������y�]�Ii��qY0e�����lUS�=�{�Bq�d���s�u{�ja
���'�c�f�фu^y鱊�bX�h� �1�o��/l�,~ҔIpg�I���
��9w���F}!N���ͯaM����t���0*Y�I�����ˁ2������?��-�%
�7�`�~	�-ڜ�`�^Z���I���ِ]>�z��
�E��iRG��8��W�tmn�B������pܩ������Xl��ށ.n����F�6�WQ��k��9A��˸�tg���:?M��A�G�"�����2%g!���6�=��%=�z->t����i��6���8��(aP��[�![s��0Ѕ�?";�\���$Lg"A��b�/�E�[��&9>6��p췷w���濨j�7����h�K��zڱ��fN6* fp����
 �d�:�`�H%�AhU���C�VM��$���o�is���Hdsx���w��{u���6���PU��E�Z��$=l>��kΞw�3#�L�S�iF<|���@�28��t���]?�ՄE!�+�\��%��)��Dx�#H�sXK|D�tn����K�*��lR�l���r������ai��so �}h.?0��G������a0'���h����qD
�'*i�=�>d*����ÆZ�)���7��x�Ӭ4�~$	���KP_K�j?*��ŶY��7�#��Y
�[5Mҙ�����E;�Ԩ���4�ѧ��rzO�z���5�c�c�C`���]�n�� ]�J��>�0߸��CφV����1�hS�	>�o�d2�j�@��L
�<R�0_�����D�4�π�uS��c�uH�2�q��#�f��2�-�i[�Cs�%�sLG6�n�)r5��{�%�cW�і�fDܝ����k�,��P�z8U>5�h���F�Y}�r��I������l��)� ��9/"�ie����B>���v��#y�F*b)�6�,�-IJH�iA���O����^�����_	�/[�M3	��3	>�z[�u���<�����qlM��>J��vm��)�);F4�U���������լ��͖��w�5�d��[��}��Cx�{�.���ݸJ�q��%�����F%p��ڿ0�y5K�8�P��K�FK���]����n�L�#��t��.,y_��t�Q�k�<h���*h)]4r�[�`�G�o�n�|5�<DD���;�9�b�7N�����r�1٩5D����
�����mf�� wBi83�*��eQ���}����l� P���[UKU%�'5��pȓ����`cp�itʔ�|�=s�*����x-�}�]�]�ˊt��w� _��VyX�y8ѕ��1^|�+vȳg��d׏۝�C��|;D�G�E��0�b�B
g&SɫW2���?��Q�Yս?�Z�� ��\g[������m[��,|w�Z��z>��J�ˀ�V����+�</��������������(��o��ҟ{��UM.�f�`\�����t�_L�Oi���δ�,��� Á�� ��\\��.�vy̬5,|�]"P��J�^�����3G�0��e��պ��[2d9k�E)��>!��7���3A-Sޡk�h����  '�����ˢ�Ռe���5j6B᷍�M�E��P{$O6zA���HÆ����o�<y54����F`έ�\�0��C/k��f	��d�S�s����V�6k<�� ��|N�3��䆴�t����Pj�G���~��E�����3���H��+�McqG�_0���f�(Y�k�w�t����To�20�5=5Z��guj^�_��8Ĳxy�Z���}��S!���إ�r�#mi2����Z
�vhh[��.?Gy�,�5��@�χ�Y�f9���k#ۤI�Tʱ΍�d���uS�L_�Xp5������i,e�=�����^(��S_(��������H������f)��ӽ�ͥE��-#���{ �-br,[���ԛt��8�6O8z�vu���͙��}s)/��L㠢.�	��� ��&Ӎo��׺"���37��=G�G�`� z@�2>��(5T`�� �Ri\㓙ʘ�7Y��Ƕ���N���V���'P~�7����-�2WQH#��V0�8W�'XyӁ���$����n�b�_)pG��T�m0m�5�c�\[T�o-�(�9�l�@�l��5A�1�bQy��	pI~���CT폽�����D�s��kH�ob�����஼�L�Ly�.`����	���W��!�n�'�̍Ғ�B��nr���~'	X�����-Y���7���o��5�;�(;.���(S6$|p$,�i΄�"Zpgs�f�OU��؝ �n�߀g	1�{=��w�`�@hg��O*��תb�WO��H��\bU�g��S�e_Ļ�:��F��֬�
:�AV�O��Rt�ҟ����W�ň���(���� V�#�a5)';j�L����I���0�
�r��٦��q�7�>���)�F��.�Wc�=?sv�o��OIuG^�kг���괬"�7��]���ej1g*�c�wpV�W�*v���$}^8�V'GОJ���1K
�OD��KR�[+��Vߙ��7�vζ?
ǣBf��{z�_a�j�!�-��U�����ҡ����L`���J#�}b绸�7�� L�cj�L��]Gu/���sP�g�Ʊ�L;��RQ�j���{�DK���� {���$�*Cg�\]�p�-���S��p����� ���K���2Y�B}�V�<R����Ez��:����5�l,���\�F������8WN�����]$��N,�����C=C��`ꜯ���iFP`�oRa�̀Ot�5rFL��N���Є.6��-P�q��T!`t<E�Wl��X!$��ґ>�.*M�A&q~���/���m��X'����22]l�����mJ�����F�F ���t�\��4�<����M_�/!Z��xUʁ���Oi�KA��e4.P��. )JYS^���6��ם���GǢĴ0����;]1�<�W��)�db΄���;g����u6pL!ξ%��<[K�9���DZ3�\X+��mf�է7��?�O$����#�H�I�*�����g���K����J^��Us4HU^|��ք�-�3�b���l q����t�K��X��Q�sݺ7+�>�T�A�6҇�&ve��
1��v��6"�hT���ѧ�N�ņep�1^���P;�;ϐ�ꈆ�3�)d���np�Vy/��~��&��O}�	��t�m"���Q��WS��T-IW(�,�U�e�C)ޝ�%�p�
m!k��-nm�!A�6�Bc!���������Ðxh�G�i�y�L�c ��%ҏ�0Fq���e� �MZ _�H�!7�YVY�8x��ʵ8+�U}K����ƅ�c%z�d�6��ٵl�4�t��X�p�Ü���
ɟ���&O;�Bd�BAk�d�b����Q>�oT��@��~��q� >�����蓖��8�;Uhy�L?f�<8+�F�J;'k8���Z�}7^ CD�@ل
�2�\Di�UՔ>�w{���<i����Y�;L�u����\�K�4�u?� _���ŋ�)�E	��]a'2�s�p�y+��e�Ќ
���Z]��<�!]`]v��s���g9��*H������N�I~����x�uV8�R�O)��&ڗ&�dW�Q�!�W*����.?���;��V��IZ�^T��4��W�>�Y=	���aDt/���/-"�Ba�#�*m`�cE|����
,�%�\s���Z��=������;�A���">J0�j3��b��C�6�Z����/�`n������'OS���iP�i ���	��睃3]<yeH���B�+�l��"�B�
��bB��:�L��t'�qI���N��9G�E������^R���^�E�W�2|"UK�+߁z�`���A5T-"���ݕ�r'���;���J;�չ��Uj�o�����/!P����2V�rBFAf�]�A�^sڀ���T�+xL�8n�C���ǨOxp$g6|V��4o���^����4�����ɒl��������`��j�p�  K�Y����_��݃�ʔ�08��xp�.(Q�c[�J�4b����1)�_t+�pn� K���+��]�wO_O�<A�ʳ�D�R<gz�7�����#����O
k���[�1�P�(�ְ}n�T�ݼ�1�yU���&�eC��BG�U��݅�dF�2�54� l!W�z�	�"�)���8�Ar����:x�;-�9�ۇTZQ���1��>�~�r/c��ɂPM��[N�{����A-!��$1� �%qt�؝��)φѥ��ͅ��2�B
�� ;&���ˁ(�'���I��5�;�I%^Õ�,�F�j���d
�5�W�Yj.�� �]V����}��0/"�N==7��1�7>p`��������,�]�Q�?������0�DBH�x�"P��/Q)ѽ:���^N�.*/�����sf"��bh���?��|���|�g&�x$a�t����Bd�$��騼mj]�L�u��Z��R~4�ZkH��_�����Wd�*�3F�k9�ؒ.�Eti���e�P�A�Ǒb��� �t��'ڱ�r��3Y��^3��u�k��o?q�z:��q?lG��r���'֩�15|U�3&�$Qк�����/�!�Z�\h�%�����:%gm��Щ�UXq�jSMA�!(?PL�G*��1�/������E+�u�)��e�}k���&���e46.�z�Ģ"h�F�� ���]�#�;�@�Fo��3-)i ��l\�Q�,)[d[�q������ ���Q����<�n��J�m3��ͯ�-��;Ti7v��;~qF�\�_c}P��j{�{��a�kyWp.�����x��+:G2�;T)e�������K���- ����=3��ȩk�X?|
-�aB¤%嚫��gv��Y||f?!�y��H3�2��G��1{��1��lZ���'�\�R=�#V�ǣ��7��Vw� ~Qj�%q��/����2�^zjǹ�]h��-v�j8�Ľ���G��/6�)W	<��K<���16��6�	k�aB�V8�={P+lЬ�;�Br�l��ޏ ����r��_�BV�� � Ĵ�G��[�mA][j�L4�R㮅j!���ꁠ)A+.�^+ �������%��c1��.nSj�	`�q���E��shȎ���4?GZs��z<�a���(^[`S Dm��F�1�w!���L	3!�1 v;�]�q))���[{2c��L6�6�\�+N�vS��� ����H�������^��
����6'����I1�T�J�=ۡi��e�E`�^�5��L,o�h�D���g�Z�<9\�������DT)��S�>��V�����UKH��4�{���j��Ql��:M�`�59(�N��f�3�.�5p����K���-��_�N�q�ϥ)����wm�wtw�Ʀ�v��{���b\?�Ck�CYM{p��X<\�6�K�����L�!'GH�u��5��]������B9RJ�㻢�C����8�����6C�K�]�j�N��(2U$bO�'���O�����[�V�%`C� ���G[�<*%�Q�JE��ڡh��g�;�ȣ'$��`����d��}�󞡫��-�߻/4���ذ@���XY�|���[�|��wŤWhv�^�i�\�:�]M���T3��{���d����w�M�w�I� %R�&#UnAϽ#GT}������c��#���zϐ?�CgpX�}�4'�q*����ă�5�W�ȍq�bH,���%B�ᙿݶK�.��I�<>�w`�n���!��Y䇈��7���N���H�#���"�+K��Ӄ�)v��<z����m��Y����!�����;�E?�D���#�#M�@K�{���d�T!CZx�+�!��f�n&tБAlB1�]rP�❲oy!1�|�p,�r�� �7kT}X�
K�+�W�YŚ��R $w��)����uny��"2�a���4p�;5��\<�`�C��8o���O� �����bvaOn�D�Y��h͹LӺ���3��d`� xE�Ń���ް� � bϪ��o��#�*�D)/k\��H��а��\H�ܑ	lC�bٹ��*y��\��ߎ�:�1�(0��f^#_�WmU[��iU!;�zq�\2^MY����R���D�ϮQ�+s:Su�}�O�������|=<5VlS$R�f:&396⪦�U���['�7e=���A�6�Ih�i�&��L�6A��j2�u	�L��^�*�E �nMa�Z&Z�ƴsj'�O���üN�
�:	E�5Mn��54�l�֠���%�'�/��X��K���|���m�?7����������Jh�+y.��j_+�Fn��z�ʴ�Y�@���t!؝�6&�O���o��%�tf|���p._�P�٩L�M�(��|,侃 y�2���̺QZ6P02M(�F�%�;-�����zc3�:���a�&�%Xp#<�����E�;�Ŕ|��܁W?�fa�'n���ޫ^?IW�D�ּa�ٳ7��rZ
6���3��A�*��iO���U^W'\�|�خ�6}�w���7MU�P.�zt����}`��{���͠�����9<*Q�y���,V���Պⷀ�fu�Uxwݴ�
��݅��~8gku?��dK�	[���5��?������W�K�l��dR�'�������֜B�5k+� v���*����l'��Zm����=�(ɽ=m߳!=8�рş���.�>x�\��l\�Gθ�a��:n��m�(�{�o簴ȭ�kF8R����|v�a�M|�ݲ S^���+C��v�!?�(��l~nm�?��&Ҕ
�=X1f�$T=��r~Q�w�x�3�ies�}!&����=6
�T���n/e�N�����.�O���hI�/�y��"��,��5_��k�)�TR;g|�#~�����)컕�-h� �p���Ԅ*��._Q�����\~��z�O�ہ���H�w j�$����ټP<Dߨs��X�'2��[�x^�����Q��K�]��[������{��Ƶ���9 �hgb����p�e����| �Y`?����R�����B��|g��[��(�x�3�s۵�:��/r.�a���RT�T���1�g��A����:g ]P-�����5�hU��Eu%��`c����|��O31����_g�<�����.�JS���2n�o�d\�o��mZ����C�cÃ���eJՌ
����SSQQV�޾�n,�C�����w��C���V����-(g��KT���ҏo�A!�\����;�fɟ#Y5�v�I� �F�P_��Ǳ�A������W����$
bqf~P?߆}.#���ܣ(BɼVD�lʺJ����|%�����C�@_����N&��?�wH���)�og�V�o�J�)s"2B�h�����W�1��&�����#]	�z�uG�U�yv��z|̤a�`ѰX�#9C��1�U
M?wv��}U|�%��.)s��>a�*����k�9�_�d��g��
���t@�sl҄;�]�Dٗ�tL�6Sp	<�)��Q�����9��I��)W�[j0|���I��2��8���\�����6�̉U1�-�-8��s�r����]+���j&�	��YPlF���sy���y�����J:���Q�$���c�F�T�薦U�ۜ6vs��b�U�򟑔Qd�X.()�����8��gM?S�(���k;r}Q6�i�`�'����;�T�Ϯ��i�׻�0\z�t����/ȑX�
{��J���}��*j�U}�-)�#�G召��I�������x ~��).�&�0w�)����]ΐɌ������a�?w�<��Y�H��1Q�d֒�� qp����W̌{�D(nAt�K��~H�D׽={��j ��0]Kj���h��E��4$���0l�;T���a���PWȘT��%��D�Û�q[�Z���,�{�M��9��$-��~~+�-�}�����~;�-��$�-�=��g��Z�e��0+�#	i�+�0�9�Ty�rk��ӕ�@E�p�=�P�}!(`�Ǜ�d7�z�r��"2]]=&�ۇ����Y��cQ�"}��'g���$�D�uᷭ(
�2И���ہӽ�7�F��K���Y"���1����d̤����f�.�܄þ�u`���7���N��27s����lUwu8�R���7� �Jzu�h-X��"5�˧��6����~���HG薆شr��h�Q��T?��ܲ>��l =��~	DY���d*��j����Ǡ�����u@u��y�%�!'aF_�9i�oO���Ć�x(�G�ɂ�xY���ͯ�Y����)�H�L	��<�BY�&��q�XH��GǬ��	�gy�v������ҍӮ4E~1@6y�`��YL�T"Q��P_u�����ጽ^����f��+�cX�aOC���LdP7����-`U<�)�j����Y�ФT�Uɠ[�}����	�pM�Rg��{�����x�)^~�*�w�4D�h������'(�#�A�����N�v�S���9<���9�2#N�	v2¶BQ�|�էBg����6�'�*�)Zz�ra���"$�[���G[�;���k�bߓ�X�]�Y�z���y��d�'�$v�>�'<�QQHFF&C5���~�#���5]R��Z�
�_{�A=%��x��v�7G`�z�S���#Q1�����������J�"Ab�bB�Q1�����{H���G6��}��P���c�G�ZoՆj�)�<�r���:�]C��M���$HiT�Bp�E�4�sl�ﲰ��~�<�W�	�* �w��Ӛ�ըF@���0Fw�`S����Q�O0���}��9���ߓ�Uƣ��L��w�����?���J�y��4}/��Q�����ئiR�W��m��2N��c��)z/�����Z����S�pɧ�L0�n~��}�</��	:�(-����`yr��6�[ ]�`-FY>�{�%�Ƥ$����(�s��d푍S��}Af��W' ��gG���O�N�[I2����8���,ԏ0�Ks=��r�(��]5���b1O�S4�!��͈�X�J+P�@4A8F��|>�HW㕟?��CIV0���O�7�ڴ���ݜP��-�zWk�c)v�bԱ(�J�~K�	�A�*�򧁼$���|=骀J�XIN�gٰ��l�.��aƒ�y��4'J����4n�k5�
��sd
� �����'�A{n\��� �'s�Q���u�(��CO��G�P��;)s�֤`�q�&x�1�E�a�;u��Њ�县��$ta��UG<���XlZ| ��|uV��el�|yUs'�3�MB��䩏���'��,�{�\oqӘY��.�ɥ�vs��=����m��_�v��|�Z�Ef�ú�T���Ⱦ��̡f�H�����{
荒�PH*1�i ����\�!��LB�T,Z�fi�V�+�W�އ>�i2V7�v���Ƨݣ0)���3U��}E��r|8c�_�:�X��3N�
Ю��r�U�E8����35�DlZ��F�A�TZ��iع�9�o�5fu���=& �(1��>b���!&m�\z��PФ����+�1ؐ�P��y��N���y�V�O���)f�e��u��;� �|z�%�I��#����G ��>]5��+��e���}��La������(7?�ά_�# �5=��2��s�ss`��������.:=8�����#z�Y��Ϩ>��à��^EP[��=-Pl}�!|�oQ���>s/�uWCY�<�H�/��s�_�=`Ӽ��I�/P�e� ��Z�f����A������"�]bR#Sş
��ꌀ�P�s;�xB�*�<;FT�+?e���I�pE�c��}_n�����s:�6�!`j�dBOk=Š��H1��?����;��i;�.(��73_�'w�t�4 (�O�ɘ[�!�9M��$L@$�O_�m/��U^�v�8�������Q+�3�Q$>����{A���9r5�2|�E �bW��4E�L��3:��a�j�J<���thCyK����3족�ڌBJ��l�(�Z�
qU�̢'~�ϐI~�柒���q�Ċ➨[<r�J��l3������G��T�Ћ��t·tߕ���1.����k){W7^	��|�`F%������n��/�Ƈ/�y�?JH
y���,���`i�]��C��L��z�P����/�"Z��m6�ѾQ&4�šWgv�~A�r<�2]F���l�.�G��/Nt�lh���X+��$p�2����M><�P���%V��-��Rn�НY��6��0%��n�k4 �����Z��-k���H;뻧=V�iV����	p��~G�8f����������o #?�?���I	엁)|�I[a��z�s{���6���+�����׈~q���R�ʬӾ/�ߋ���Y�'O�Xhw��ta���:�nz��f£�ui�wO[z���;q��C�l~�_��XOwݨ^Hj*�G��Ke��>��rS���q��W�Z\Y�&iZ9^���3\J�t«$զ~\�p�K��}Ξ�:��MF�-۲g���g�ؔ��!���kgoO�SLK���˥�	'r�����vzXV$X0������F��"�0@Z�/ͷ���Q�]#	���ix@$�m8d�fɜ�i�o���Br�XM��
��%�q�tq�2�����-R&�ڥ����'U{�$��;E�6���Py��Bs�Z�Iۇ���ų�w��c�B�R��n�K�~���$� p�'G�XSSsgh R1t.�1u���LuB�E�zc��
����YQx�����Y�5�^'>zf���C/�vz;ʈF6�63� (�6s&��ll��<n�/�~���pnZ70ɏ���3�~ތ�~�O.`O�Te`	��Daoƀp�mqH�X�mP?*�j/�@�ϣ���{�lh��I8 霎='Ú��th�o�F�ۢ����:�!��7!�ʸ�?��r����~n͚�]͋۰���X;=i������;�H�a�v��x솞 �*�n���}rm�c���yԵ/�rMO�7�:𩚔���G�D�\�T��ڵ�F�����rj=�۷����߇���FB���@C���ONt3��'�� V�n1r�_��sB.�Bh�[��<x|SH��/��1$QX�΁�� ��awUs�5�l⽵����7�i�fCOr���&`S!k!p�v�p���|r�.Z��ϊ�E-ۮm��� �=P`����c�ʪr���]���:��|�dnr|`��b�)|�A�@Т��Bq����.�Vt� �8�su��HSb��W���Ku�b?��g�1֡>����#�wF��:�=�j�������4Ыt�)q� ���
�٪=�%C���cK`�,�S�8NXYG�U�p��avK���{K[*P��������%���t���N�=8���t�ބO�E�s!�[n��ꫮ�l]�S���T��}ah�����z+���LoM�>�O�� kw��LY�̚��in���v��V@^x��o��;%�1�N�98��!���5ʰ_�L�6Baݗf����Sc
|�����uӊ�����0�Db��2	�E�R��D���~#ͩ�)�'��"JP%RG���L#2�~>������@yìz'�S�ȩz�WsI�7��0A���/M�ѐ"�_W�TL�3��K�+��gmZ ���<�a_�cPG|��\��W�`ق��ԋB��G�baK�T)�pv!	4�4|��Q^�1��5HG8�����P4,L��v93���e0  �<��6��U��SQ杺�!~jԜ8�.qP�[(�]f����(f����&���[�T�Ǵ2������-s�+�I����1;�<h��/u�R�Dj�s6�l7�t\�P#�2g����P�_4-���4�a���M���¿�[�r<H�B2PAm>8����zJ��:D͋c���>ndݔn������^��oh e��٩�6�K�W�d�Ofĸ.��y	��P��*V*�*e��X��=�?X!�\^.'��Lϻ�2sޯ�7��B�0���=P�/�^�����+�A�*ʹ��dÊ>��G"�'I�c)���4i�eai�(�k'B.�8�Rd;i}\:�����ν,G4䥱`\(�>�H�ځ�	�t�uJR��`��$�E��(^�M�/�~"\L&��v]���љו�xN|��(롇�X�B`O�%��I�Rܚ{i}0��#,�\C� f���^$�9�dL�ϝ����4c5[X�
�g�Q��=*Y�y[I&u�Uؠu����5�%��ɜ������T�T��� A?*\=H��"=��Q� �ŕ_I�>xo��9�&��Q�tݺƒ�9���uު�O+4n2,kE�0'������0R5��z���`�� �k����7WR��G+����Ry * F{�q[��������aj��V��u�	�(>EV�ݵ��{mh�)a��x�`�:��(ù��&)S��(�ɱ��$/h�w&��qe�+V����W{Q6X��}�qe�ʀ|'�G*���2���fW�^ �� �_�&ъ��Y���n+�jX����*�k�b�G;���B��!�$76�k�7v�QO����%�E����>3��f�7�p���,H��t[^<R?���>1J��@��8�/)�@��sۀ�"Qz��쪦�^^���e��e1�jW����{ �j _�O�ڌ��p�{t�`�5�֍sv��B���c�/o��%�[�B*|h'���+N�����BF<]�<�mR%�Jċ��.5V���K8�Oc�1��Td����4���F�rV❂�����i���7^nh����X�ne���y�f���<�M U,(yj��\�|^�I��%漰��-�Q���2�Y*�Kj)�1ꈘ�K�6eJ�'GBC�F���R�>�f���ָL��X�ق������B�
�|�	%�Bt
A�f'�wg�V�( 	��꛽��rr��GN�9�f{)�W����k�c�dV��8����*��s�k,��zu*��}���$Y���T��I'^�z/�U�����3�U ͞`�t-&���R��<���LQ�ۖsoQj#IH�U�19�/�]R})��CB]e�2�(#ʇ�.�ӄ�SR�#Xy��a�F�f(��Nы�w&���IE�	F�KuJ��gjؓ!��c��&��V*���fA�ή��觙���E��֞�j��������(c7����&`�!�—e��ՀCS��j4��}��"�kĄra�(�����9z<z�<�H����k�γ(����C���mGKIq�.Lw��ei�v�A�P�l�3�!c�4�w�)6+�:���6�e�Y�U����ej���g��U��.J���V�	��_�"ӿ|J�A�n1?�Ϳh1U!u�eC��n!�E�aE���2뉏������R�H��Eघ�+�*����ho�s�+�K�9���m��׌��b��be�BGZ���9����߾&i�t����ɬ`����Kiŕ������&�w����Z�S%� 6�Ƅ���C�<[]x/ch�W���"���l���=}a�mQpؒ��WP��T t,�.Z:�58��������!�����'�uу�=4�k� @��E ��zI��?n�2�����+mq�3*���1ˉ��lJ�� ��5�OŤ�w��S5����"k��T�|�4@Ǭ1O̲{&��3��9Ƚ�ˑ�;�z�p�Ղ`eē��2�CzLT�  i	�{k�͍i��-�I 0N$9C�/�n�*㿙�TW�)3�h��3埊s�����b0%K���{���at�o;�M�P�z�6r��� F�"�؍g�W�Ϟ�#��wcsaG\���D��D�K�T�s "9�0Gp���z�j%�i#̐���Dj�J����l��L�t
��,�a4��D�L�e�BVu��xi�`���l�49ҁNs5�U�=���Fn�e�U����(�[�ò�,�6g��E`[�"mښo�ߍ8���ͪ��z�=�%p��gvw��&��(���������f�jk���\� �%�q�=G�>2������b���AsMU�Ƞr��VX�]��^�~P���V��W�㳼/	�/ɤJ�� ��^�i�o�}�R�{�Z��2F6*�U��r��N�UWK���x��LCR�=�`��!�1�q4�\R�ZF�u��H(j��X�wO�N�0,�=�S�[�O
�4��!S� �A�V���"
�:�ʇ���q�(��,��*6'bM��� �&CI�z�>��_��<�Q:Cw�b'ZVA�^�"3�e���J|B\
#�L	��~�TgD���b�h#�X�:��^����C��91���� DOy	�#K�.!��\���x�����T��>�q�ͳ��k�'���ja�@2˞�n#�	�t��v��� �ugP�[4Ih�<�sٳ�i|�N!p	0���� U����Z;w��"��!����L6y��Sr,
��<�+��$?�]�����qH�p��������;䩳��W�V�y���!�=�� ��Q�A�U22Ԑ�rY����8}�B�LxVb�EIՃ�H��2�w{����	�7�9�>�9�O�j��%Ϸ�2�~=����pLal�?���>�0��e?|	��/���y��	�a�4�3ˊ.�a~��s�n�4̌��!o.����<F��H��ש�ݕ&7r@Y��Ǟ��툵V���g#�����\+/��@��8���K�(���.���hhi�_;����
oU[�
a.A�u��fK�6���
�[��&4Vmilԋ/��= �.dߕse�Y��,����U�������2��%�uUdg�~: 2kG�S���4��l��OaU/��~�	�rp�iȟ&�z�P����%���QbE~��ƕd3��o}`����x=�o�u�Z��[s�w�h=�-�%�g�:��"�"W羐@�Z cO�7g�Dm|t'��.���
�p_��M���a}�����|��э��r��;Ĉ]9���R�@�d�b� nO�E��R��WJ��6)p�Z4k�
P���~W�v]0��	J�fV�e��>�zy���Y;� �)֞�d%߫,�W��qK%h�:�dݾ����#o�n!gc�wB7Y�������El�p��s^�B5L��h�R��^���\�%�/�_W�g�6$]S��k�D@ޒ�/��Y�e( .s]�����}��v-gN��v"�F�"���?E�I�-�5R��u�"u�d��tk<�}��n�	mgnA�����4D*u�d"����?�!���3�	f���#���`�+��o�����4S�/��"`M�b�t�b�]�EK��o�y��og��7����bˋZW��n
~�Z���	��ĎVf�<�~���麨!�u��Õ�V����d���9�<�����*	��`ϋW�G�x�f�8�/�E�;�̄�۰�ړ��c&l,����Fe��б��x�����ԛ#?}��7yf[2C�Cf�mJLs٭\=>83�_��`���t���+�i/��o��bZ(b�7Bp�� �D
�9�L�9�n��k�A��rR��n](�z%ҭ�uu�<�+b�l3�\�8���ng0��m������`$�oq���_��n]ۥ�54n��vo<�J���Kj�";�ݣq����^[󮎀II�P�4��X��� u�
�X|��З~p�e�X��&*^
�RI�[�Rci��:�q���,����Kz��jcC�i�ڐ�r9_�D06��p(�H�(��ґ�Br+1��]1ѹ;���{���pN�©�+�����?������TSW
�?��5��@}���#�������%2��P8n�� JQ?�\��-nR��G�n	�'�\G�XkP�����:B�n�ⶠ~�
ib/120C�糚�R��q�%�7��|������aqCx(��A�4�a=�A��<�N%D`Hs�ğk�Old��R�,�{:�7���m���>��%���y�"Ȳ��E�\�D�:�o���j�#�[`�n�^�Y�:,�v��B��,����I (�-����wc�\�SDC橚nT�^D�/�ԖV}})�4v`����^�Q9#�X����d������D��j�����T���<�Gi^#�Y�zo������wwͤ�a��㋰�Fd�>m��Y*��h��<�F)��) pH�ز�aU��Ŵ@����T.<�s��D�����m�eg{,!�"^1��`���<��B��������~.l��[��IIC��>�ಳ��OPw Ft"�%�B?`����'��Q=`BZ�(��c�~�K���"b�Z�BUu�8�cf��zjY��{�m^�櫣���Xsf��z����ۚn2p��M��}l�<C�� >:�X��I��,�s��g��M�AŢ� ����դ2k�7�1��V�3od�&�x����({��3�wİ���#���]n�Z�Ů�B�Q���c�2���`f!y��S\�0�]4����J*t@ Sz� �i��L��%�h�e��W4@�+��#��|^��ʿC�Z����=J"��a�d+�ȵun�9�:Xɖ���pf�4��[�4S^q<W���l8��L�D8r�����v��Q����vX�"���}QF����q��-����d������f���Q��(t������̽�0kB/��IK5$�C�ٚ�kq��Ue���:	k{$��4��1�j:��<��8I%<[�h|)�M�+b�I�\���B�r�����M��c����w0�;H�1~��e��4��{��$'0��v���)g�����+F��s2O�[b��.��~��V�	�
-����J�m�~j��S( +��?�Y�#�)�g�F�vIlvUh����vT�gh:	���z�s7ե-<�������#�%s���w��)|���Ah�|�̤*Y�m�N>?P��{�mcl��5�%�]=8�bq��*�y�(�b剚��8a��rs6���x"���o�� �;%��!uUX��P�Ŏ���햷S���4�sy���-�!����`����[ ��R���Rv0��1�x�$g��ډ��FI3�'��^�����3Q��6<�\�g�1��̒Xs��պh�.�kW����I���M���#oh�"�69�WOQx�`�p�?������G�MY}P���>6_�7���ܫ��lY[�{�?��H����~I�>��C�I�rW�;lx��P�U�q4B�w-F�q���Z[-�(KH��zP�0'��S���k�������]'4�*�]ڏ&�'��$6,C1�R��@D&� &)�ϡz�������(�Fy�sT�o�ߦ'�z�@MvzB��_�f�Y��PgN�ﱭD� ���w�5)b�����4�6�ԉj.��'��^��B#,�q�S!0��p�3q8��Zrg3����ru2`ޏ(�X�1 ��~e���~4��g�*Mƾ'�,����fn�x=�||&j�M��V��Ί�sݑA)���&!��O��1:���y��cdՆfR��-QJ:b$�MK5Xs�%Z�"Q�~T��7��Hw��xˇ��'7r�b�����#�S���d�N{*h;DP��fi��To��9����
�-�|��{�/�ڽ�W9�g#�����$'������}�y~F��ǰ!��2��\����E0!)���Xp���j�,Z��pq��ׁ�>3�K����Tn!i�C2�q,C��߉=�����S�8�����!�Z1S���R2.t�c@HVCƆ�B��!P.����tg5�[����^�a��yӥ3��Vm"��0��Ο���kf����4��:��gan��M� M]-Whj8=x���sC�S��'�:<ww.b��.��T�D7����$=R��`Mc��(V/v����Į�,�0@������/uڟ)Oɗ�ImG�#'����\џ㤂 ��f�W��L�ƼVTɻ��rVz7�W�b�ڴ��ET
�7ډף(-�u�J{S�S�����]�n�23Z����"�zݴ�h���F7�*��!��X�
[�b=2����]꯶�v�]�R�mnR�!��~��GI�'0�G�]�i�q:F�+���\l5M�x�?_����!�$�R�x��c金����E��L�
��{%��I����ix^O>]u���t�Kl�u��OX�T�pT��:e���_���p+Yһ��ѷa�P��p��u%Kj �x[4�a���Y�C��z��d��x'��
��f�@q�w-�1�VU)��]��/b8�t���K�[g�P�N`occ���śT�<WG�I��v���ǻ�?�V�NGJ���K���Q*�M�z�˚䙗���tu��N*,��P���w�}�����+��=޿щ��Rۗ=LдV�YYn\��Yrs
�Y���q�ix5@�H���Fq�h���7�3aL�,��u3�5�?��eE�tn&�q�0fݾk��񊎟��t��P�J�{]�/z���;-�r�4�$R�^]]�ɯ���M�2נ��#1;��ިGKg��������-���u(�L槊B�.���tHs;�2����5
��
:[:(P�]�؊	,W���ā�"zA��ݏ8;40��A�B�D@ &�E�c-r@�#|��4M�*\L��9����RD��Xկlv�f�Ѥ\�p�]Gř>��R������'�t���ǐM�p�P���&���a�>�m�)�q
i(��h�J)P�ݢ�5V4�-�栁��˨T��� ,����������n){=%N	=�_�|w��<�^O����[�Q5���ȈE&���2U�^�S�`���`��x�k���\��?�!�C��)�O|���L����Y�l��d���#����p�m��B�㟈v�k+����S�8��
��ݖ��t��.}O�R�Ax��T<��vB� �C]�� ��8�kyiF	��ޡz3��S��V�>�ޥ�� 	�v�"Q�aS�p7�z6wF:m���eZB�s+ (O��#��a�Ƀ�]�$;�CZP|R*J1J����v-�/Z�4g���R%.V.yHqv�vΘ���c�SYVe��:�ߏ�|��Xl$M߿G!��g���F��&��G )�}�W{�9Fo/�V�˓>�'t�%��޳PK7�4�e^���0�,rȌ@R\�����g�'Z"���h�z�kˑ	�#$QC�/Q��W\��
�t���`��ğ�m�<�\�~;�5j����`'c�t�
0�U��Tj�������* �,�\c걑��
��D���;rNb`zqx�� �\�զ�;��lI����'$��ɨf52�9�z����  ?��oqL�bw�R}���_�29N����u�L�Of� $�PLg^�ź����{�.��U_�u�S�	8��g�jB/¨.���p�-�Q���Gz�K����|J}��b�g�����:#S!fƞK1"���$��nvi�JZ�l�� Y@1 �P�z��M�%i���["S���z�磴��d�Ӟx�靶�6�5��H��B6��9h�@1!4����F���������alI��pޞ{��	F4�?vE��2I�:��@B!�A��ߗ"�����z�x�@Z{u��Fӡ��˳���G�.Sl�i՛v!�����@���bWMˍ�;���Ҷ+?F��k�&���1$�D�و�27ўޥ�lR~\�9��<U"��H&�Xe9ӝRf��9Ƽ�q�z;�'s�mL���A�n�����kξ� ��������ׄ�+>Y	����F'��/!z���@�*����D�VDf�t��p�h���o��=nl��-%�+�+R�i~`�<�f�`�}��iB��E�I�Q;����`�2CR��ˍTc`9�CМ��m9�5�3o����-ҳ�K/㻴\�`����<h�R2�S���u"L�	�Y�m�.�;�Dd^4%��Q&ĕ-o(�#�c	�.�������e�u���ֲ4���mص90;�{~��w���n�X�Wv����	���4�ўD�}�"�����n�C���0>#l�kM�J�/�������(��XTFoK(6/'��)�xr_o���5+���x&�CT��w�3�tDj[�!������樓���
s>Ձd�Y䲗퀞��nqXG�g�,�j"�p�ŴP�ԓ�N��r��"����ȝ\ar8XƎozhukS�[HG"v����_�rk������t�P���P�v���U�M${+��u�~���\&�L���ī�ш7a� dAr�,��4�A^��S��gF�@se���?���h\�;���Mt�e�H�K�-�U����f\���18����z�,���-
3�I�������4�貫��F`�9و�5T�B��=�����q�(5v�M,-\���S�����x��JPɋY�B�H�9޶�!�-K��03:��W#J��YV�Og�IpK~�� ��*2@~�Ѓ��v�K��7e ��0w$JvP��k���=j��������t�c�H�j��@�d�i��;��l�b:��%4:&�/#g����S�u˵*�qHe�s����4���x��N+����߆\1x��v�c�d��HȮ.��޲퀛�=LP.[�O"޳�R2�%r�ן��s��������#�G�ӻ���1�GҌ1嶢_����U0���ǳT�E����>D���[b��>�M4�|Xݲ t�`R	��F�	��꘴A��^�4W���Y�&�f_J�39��w7�&�^��3͑�e���洁�ҟ�z�R�ೄ}��-�X�HM��x�A���Z/�	_��s��h9<��7�M7�=�]u���]*���>�BպJ�hs3rG��g��gTK��^�		��1F���0_?ċw�=.��h�299�^�V��h�ueX�w�̔eS�Z�%�ҥ�Slq�H�j�D"��|�������@�r�3��&`��*ݽX��]@4x0M�H@�oэM૘��m##���G�w��0���d�SȾT�D�#1CqJ��ϫ~di��[k�7 v����:��Ys-m8�������c�n�X1�c8��U�U҅cP�N�5��8�{����ĩ��$)�2�P?�n���M�:�^gЪs���F,4cg͈��K}(��� ��J�mf���č$����f�Q'n��"��?���|j�ͱ�t�؜�S 8R�P��f��������7(�u3l����A7��$Z]��o�H�o��Fk~���N�:�o�7�+v��e��`�/
Ȍ�����T{�_�+�$t��3M��=Z8��,���G!��w^��׀��|��
*?������d�$N�������F�s��+%w]�_���g�A��{jZ4��v���_�j��=�kkx�K�H%�\�&|�C�ro�L�+�|���/.�@�<<�Xq�ιlr��͸���ğ��w���j]��pLQ�5��,s��G�TE��,c�?S4��y6�Yp}�2S�PI�O(F,)��]х)ob����i�]�����#�x�Lǭ����{��� ��4`<�2R�����n�E�A�r��ҽ6K(Ï��U%��q=��Wy݁��>(X�����J��0��C��?,�t�}�Da�<�=����ċ�f<���R����RUfU���(m+�����#HCy,�*PL�y�a�Q���=:��To�&�k�[��Xv^C>�%k�w�����(�l�4gi4���'��vx�c��2�3�ж�c�� 8k�ߌ������R��<�5л�5�{td���T���k&L���S��;dT����䏞�t���I1���YkA�Bk渹�!�N�$�ߺl|*��F��6v�؝��Iw{o���+��M�cMA^X�T�'׷�L#���G%F�^�C�'�`��A���A�p�I ��+[7܇RE�Z�"͚�N�e'�df������سvu*�Վ��qh�]e������ dMW\�}#�:����glV5ة����B\p;��������a���uH�uk;NL��k6Z��^��+WD^:�ϫn���C���_�u�Q��'	�+3)�(������'~뭦��"]���9���y:�O��G<���/�L�BsR�3y���F����%�\T��ODeW?��Dl��7&R��vs9|b���6qy>���n��@]J	*�.J7�_e*hz�«8����q?�m	v>jf���"t����L�
q�4�_Nؔ�Wϰv&z�y&ʾ1���翊���TB:~V9�X�'������!O�T5?�h�|W9����/^�ҹ�.�D�0�p$ׯ�J���Ѫ�s$��Clt�'w*�>Q|�m#����Au�;�}��Ns}������+z�,�S�Q���d�����i���*�1I���0��̋<����p��q�
�fm�/T6[�m��������|ov��U��C%4v�b����0�)���m�GR�P�϶}�GB��6����E���?�ڔ����O;�p��R���J��ϭ^i�D�}��V�E-�P����O/~����Q,HړH°��F*Ȭ�/��M�y���Ѵ��X�r1?�&�,��( �W� (%A���c�*'@0E��C���(2�!��oڔ8q��W��i�Vu��Vu���CA�r���;�=NH���y:�6@in�%n��B?XqP������BgO~S:��![?9�����1q�-�s/����V��� �[t�I�[z��Y��� ���R=�$���T�tV��K�j'kX�Te���I۩��2�>*la9����N�M���'�7;E R{A5��Rx�U���-ζ�7z$W��B�v��ϟΫ�O�w�<����7�q��Ɖ���!C6�>s��`Ρ̠7���D9��9@�Qf�lkƵ$*8$����Q���kFw*�Ip\Q�gb<� �L�rd�n&��DP$r���e�Z/�+�i{ʲ��1��L �6�]�;�(x	U��Ŋ�J^a�]-h�� �����e���������+�U.�cd���Y�d<�o˥T��*��5���mcײk1Z��B�-k���\u$>��,0����Uè�O�h��u���_3�4�z+7~�q��~{'\���9���n��~�
s5׮�S�z3�t/Bܟܧ��,+���wK^x>P��7�*�P�{��[Q�����غ�F�Ҝ�',5De�:���;���S#}�~���������<�2Oe�SF/LST�w/ٖv)x��y+2"�2���5 ��"��h"��O>X@���| �o�]��!P�,'��A�2l'�=���Zq��rf�K�/����Z2��LÖghC�}��F���h�ޔ��9�����J
��npUs:5q�I���Wb���R�L`�a7%�C���uJ�q^��\����8�\uz��sf�EG�UK�rx���|%O��+�cQV�p&_|�A�k,��M˗������(2t�u�_>�5a�3�h�O�;�/���8f�'`�)ܦ�iY�#�dQp�řV6�:�y��!p�P��R�.����;�4�}��ȇ"���X�)L{ 1)�}��td�RJ�t�9�|f_6�D�d�<w$z�Rםx��a�����Uv�j���Ď���Y���!{���s?�]3���ɜ� �qk��/�� �p��C[� �'M[���V���Ӥ$�F��F�v7X�V�ٮ\�>QN�"�N���-�Ljxx��,-;v_\D���j��(�$	9*Y�&��a9FR���ɓ��ג��8���d]Ŷ�k/>]�t �Q:��K�O^����������Pj1��ϐE��D�p�y$r�uѳ-M<?�!��ƁV�77�ʃ�l]��-�n��1�eI��k��̕���-��9:��x�|�t��ҹ�M�1��-^@��Em>dN2��>��Na�e桠IT�!vԌ_}{p��$�$q&_(d��de?�U�<����8V �Nd�9u2'[���Z���r
��jyð	�u��
�:k�i���2q�T��7��9����^N�'e��zg�՜�FC�S���MTQ�x*����ՖLS�?61SicսTqx�,�ܒ�}%���A��ﾓ|���%O�6�T���br��A��a\���� ?����Q^ڿ�ak�ތ�t�z��N{,�_>u��wE�lMl$�N����m&��+�e��Lo�¦�/��Њ��76��Տ`A���ζ���4�&Tޱ��K>�ϗ�o�7I3 ��?�m�>�	�u�(��ɫi#i�� Kg\���a��{�D:P.�҂E�G��U:���må�o!/b�K8A7?:U_�?Xw��WM�YQ��&i֡3+�
qMtgA20��$�$	ә�DJk690J�ܳ��=۵�ߓ�
r�@|��z-�>��}�@�h�8S��n�GE�1 iQ���
΅�_'�s�O6@���n7ΗL��4!��r���0*^QFʪ�AF܊��,!��
ۀ���n���C{ .W 1kϛX�� ^2��]mBv���ߩq��+�ke���2AB$DU�+ހ9j˲2*�C�TDj�0 �-���"7��"�b�����r�o	�tM5��b��K��Z3�A�-a=>�V���}���<Qi��;�D�������*��+��e�:>�ӄmT�:	U8�z��z��om�O�lI��t�1��Ȅ� ������dטi���PQpE:����Kj�O�2��G�Ř(���n[����J�v�D�H�T�c�/0ۺ�������SL����P�%�$%A�M�NchG�V)�M��&x`qO^��E|]�SM|�l|@���Ѽ�L��n���̹���v��*	��@��#�;��T+�6P�c���%�\��L��|yaTd�\> ���r��-ȩy}U���L8�x����`�w�)�Ͳ5��!![,��Z��/;��}k�Ǿ���eq�+ /]��������j��Y��Ù�3����- Yi����E84�B �琜Ur(�ͷ�v"Qo�<���/8��T'8ٶK�cV׮s�2Ά���)Kcu�r�򁗻ӭ���M�B��l�S��fڄ��7�?�?\9��s��U"-{�w7���5oP:�I���ϢlD\ݱ���]�L�K4�9���nk�`���EH����_�3, �c�ZI\Jx1�r��r�{M`�S��]�
o�/H �o)�e�ޯZ��N"�?Ђ��?�[isّ����r�1X�T�A{��^wX�d�DW�<`$��G��>�P�������yv���GU!�q�l���p��<(ߪ�~8B��Bo�QW�sk���pkP	@����s�Rzae�@A����/i���*~6�,�W�M�ﶓ�i�_���K4
��5`����$e����~����n�!"�s�u]7���H{YŞ0C�k��m�3ј�p<�L0�@S.�&�-{�S��$C:�F� ��	���Ǽ��25�^{ݽ���I��������̧����� <��r�/0�M�1*�и�r���D�՚�8짦P;<9(Q��@�����}_��<"�!�L��D��<2o~�*�ct��W�k��7��Ѫ� C�mJyK*˴���eȞp����'k�6*-�����D�=�~�=Q�$��<5w��>��I�I�rE������0J�K�:'[?�B��0A�Jf�z\�!�K�hI�/w��>���:�l�k��&�`2�5������->i���5�	��� ����L���n�g��L�!;g�o�v���2h�
���u���P�G�?�>���2�����<��W�N�	{��w�i:�1Y��0G�-(��O�)��2m�؃�&/�ڑݠ&z� ����:e��A1A��0)�����TW��vi����0?8|
Frـ!�u���Eֳ{o)\�`c� ��A5�y�,Ջ��dbl��aI�kAȡrd�G���I,u�ȭe�b<wÇ�zm9N'��q=v�:Ə�=>���f��EC�6nSJ���l��(*
�Jl��	�މ2U�Y8�����h�۹�87��u�|?��j`�=C.W/f���+�\{�P���#"�9��L���F�� A��>sl,~c�
�-H�}�& ]͛��?=V��g�����C(�6�Ҍ���](�hB�t�)����o.����{��B�ǜ)�fN��N�OA�a6.D�B^A�"j��b����_�z���O�:6/���<Ƌ�`�I]�69�$s�����B��G����X-k���t�.]�%�a%���5)�KPH��ɠ;NHX-d�� ����0�R��j�J�h�b$Gm��Ǭ�}���$??���!֋A�t�%k0����o8��Yj{��N+�F�B/"��5~��R�I2t#f�/����A����H��Xh8����O�">g'n\d��ó�OP��� �?g�]������x�uȾm݈�tr+�ľ �|���}䇢�E�|�՗�8TsM��Aآ�L��ռr�¨.  (�����'��<{���I 즘�n�5�
%�Y*����z�%���m���>�ĩ�>Pg����wK�	�i������o� Um"�Ga3�|О���X6r0d6�]k!�ʾ��Xv�@V�h����\��тDs��V�{KxC������Q}��={��%�}�6���z섋��V�����ꗊw��?��v���(��a}-K�ǔ!��\͹zJ�HI�^�Gw�Э.$��BgR.|�P]�����(Ȅ�E���!M��
��'|4�<g�t#�_[�0�ڟ�Y��V{�g��}`�l_�LW�����U%tOm��4<?�"y��^)�	!��,{j���R�LF�_rg�~h�Lq�X����)��K����?�7�?G��