��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<E��D1�a� �:w��I�ukJ؉��Q�*�)m���h�����g5A� ��;�P"�n���{�4�J��[����9���<
c�;�Í	��G%-:9y`˞\9�|��I|܈�0�)�j��*u��w��y�����\�=�
����Rͩ�<��*V�oX^��y����� ̦����:��������F&p����^:� �<n=̓K#�k�1�}OVt��sU�Ks��.s�Z�AkQ��� ��E�#� #m *�3o皔�O?N!̇�ys�s��X͕X�pK�J��7�������py�UA+��r��y�e�[�>
���>�W'�><T���Yx���5͓�
���!���tw�� ��1p�C:�a��
�jY� <��!����C�+C�S4�D~%���9���� ]ZJw~�Ѳ�}�@�/�yd���22�����/Hj昖gװG���e���!���XFF�L��E�Ғg��F8-@]"tR�!�Ӟ�� �@����=w�O��W��zWg�F����@k˳7�3>r��x,1l�����)i@���:z��5�)�g�W�hM�C5�R~Xu_��焑U�������V�t��`�-.�0@��.�b�S�k���fί��i�=wV��X��I�y쑚���'�GL���C��(o�ǋs�D�+#����u�o����W*�&���{�z�'�����c�;�����@p��$�7d��,@O�[��o
��Z���[��><E7E����"�JAq�ONŪn�k��d\�9:�tr��jR�������z����#.�����ʐ�)+A�p��&*�iG��� �b��kNS�&�m\Ǫ
ꪤ �o5z�4��$1/5 �Z�)4�E������,�/��fNZ�rW�"��F��i�~PC����ʸ� �^?��z���M��m�튩�k�@�����pC+�Rc�_r�k ��nu�Y�Ǌ����=��e���À��L��Q�C�cHrh#��FYD���tX�&��U���:����a
��.t�8�ap9��p !��-RH�~^M�ևkL>wa�����C)�5��&<�j��`&pĹE���b3�&�,8���Hl����&��&��%�C:L�&��=���o�ԗb�ρ�.�;)^�gt��~ő3��z�d�OZ�]{nَSR��$t�  q#�0 �*Z/���I���%��)q3}URy�>�>��X�#�N��&M�o�+E�h��Z)�z[�7{G�2��e�L̮�pqV�!7��!q����&��VD��Т�n�a�[Sl��P?�GB�8���-s�5wF+'&��)P�)�83TsK�/�]�i��h5�n�`M��H,�h��9ɋ<��2��zHZو��4����dw�]/M�c�N�-#�3!U7��f��f
���=����αW
�e�YPb�	][\ͬZ ֨4Ny�C��'1d�?|��O�.�N�a�a�6M��&M�u�
ڮ��8m��#��'��]]��կ�i ��/D���E�!y�[�ϫ���m�P=��z��+.{1	lq>
Dc���-��ϭ0y���@J�7�ʋ`�8V����'�پ$Ef���*x�1� �Hs���cE�� Y�d�(�A=��]�q;I�`鸬9��t�����n��PE�W"-R�0��6��뀝�Q~�S��Ao7���4�~���� 倉,���e�˖��3�>���)^a>	�����l%��2v��U��ul:@���hT�f"}P%���b��z�{�Mef兜2���ʵo*n~�w�q��U�G%�9��gPZ��'�����~%�Y�<��	7:F
�y<j�����6j�T2����A��<y<�l���"����/{���#���f��ׁ}��2�y��Yu=f����l��Ci!��KG;�<G�K��f�*��c�ݚc��!���&���|-/F�����1a7�?i�(����]��w@l���w��7���'���{_A��F�V��}�[�/ZZ���0[�k�O��
*��dt${R%��g߮�-�/L�)�P��Ki�.��f���2��u�M� ���0C�~����r�}ںۥ����kR��֨���lX��BATp�뚠r��A-܍czֶl&�
�2�)��rd����ȑ�0�_"~2�7\�9����l9ZDk^ww����x�����y�CL��s��ؖ����҉�Td�̐��M����p�a��};�q��ET��G�r�a�&9j(午U�O��<i�u��}8l0�ڇ�^�nz��0��8���l�/�#�'1�����z,�_.Kh-�+��T[����=���N⛘;�C�ژA�����1B� ���Y}�N��_XxЂ�ǹN3�=�"k@�D�� �\�&��u�O�-����r��x<�9 ���SE3���(A�w��4���SG˞���k��Xm�E=��U�m�U˿	�H2ǜ����c0l~��(^(��$�lLe���N<Iޖ��m"�S�[*�y��V���u��XwL���	�Q̾�\%�:��\i��B[���jߞ[�_w0Jd�B�]�'�q�MI��8풋YP��c'{�K3{�wU��J�~I�틫����O0������↴�K�UJ¦l�q|!���kW)�!� �y�2��*���<�n� m�M�V�Y�&]�S��[�oovO��|��{����Jiג�l}�(�c�pSUE���1;��f� ��}	�M�g1� �.'{�m�o�o� ��'F�*���ϵe�����l��ѩ��%xź앳�o {�Ά�:��y���H�U�z�J�и��Շ�*�&'�;]>8�e��n�-�������
 �!�q�Ώ���M�g]�˼�ͥ���-;��5�}��8�5A7"�c���,���|RA[��eҙ�G�V�r�a�b�����BقV��<�� �.�/0�2+݇]�}�>bю�LP�]�^_#P����Ǌ�R=�\$��7��f��z��_+�TGR��xXW��ϲq2��y�р�&V�	�$����'2$�`���>�&�ԇ���"��fyX�8��E8@��Z�ӧ�H�E�� h���z����|����U��2r��LZ��}�̒I3$<�8��\trϝ�UiW�A�_��������s<�u{0���f|ja�_qo�H�sڼl��5>[�Oy�a=*?T[�����~�����ŧ��A#x�,v%Z���(+A��`�hg�_��9�*�D�6�����1(���/����t9Q���} ���ɞ�Nn؍=ÑQ�����i< 9l��펿�;w%�u@��U\,����=���Q^�Y=�����ٶk�]uD�j� �"Cx@������
���>1�X���av̡F/=NUd<�	ﳞ�q�$$�q�+%+�����֦-�b{�=4��86hu���� ޥ�����e��K��N���ip���I
#�3m�Z��vK�A���X!�l�ک�r��*d�((�E;��LO�0S`��%J���J���gH�$�7�o��G݁�M�Ə)da/	;�;=O�B��I��;�T���/��q|j��l��ɧf����+f`�u4γN�k��Ε���̡���z�����vl'&?BU������e�`� 5*�����`��kfK�]N�P!�<����>/���s?����g��5U?S[ ��2�`��ȱU����u������É=ϻ�g����Po-S��cCa�}���a�f8]�g��c�K
�)oLd�ɷ�$����N'^~� ���7�q'�b�d���XZώ�f𛮀z��FTk�1���|`�'4q��M ���j˔�4#�_A0C/��@�)"h\�3��X����޵(�(�tc������p�Й�l쳢�[�..D��d2'���O i�T�}t,X3xh���9q�5��1�b"�O9RV��s;��(���}�[�b�X�.�r�*�,��5/���L�l�­��q��`!�+e»=��$��s�'�>U�����u��qgòM�_�܃nd�/_��JS��k���s;i��� ��G�F���X`�u�����~�o�nPM0a|�d��`H�^ǂFT��+^������#�w��2H>�,�@�]�0���z��Ŕ�օ�b�ev�R�����{�o�n��O�4 u�O�Q�j��ы���u\��/d)01v̻a��K�H��z{�phS����!K~�F�]d���g`�i�r~���#����>����5�9̓j�ʹ����? ���)\�9������6H�"2�����M|���.72�S�O��[���{䳺@��1����E!�J��|�i���+��pd>����-�t����K�x��\}�o�vQ�Z�s�/?�O����u{�/w0	�
x!^���R���U�L泌�s���pw� �P��z�Z٨K�#-6~��҂Ҿ�u�q@yAZ](A׀�C;%gN��\�؈��~����<.J�N�H�k6����x��Gk�K�Usb���b���ᆜ9�/��>��W,ن��JXd���z�a�q6�IՅ�U�ή}�f>y,�Ǎ.��C:��fR����lBcCT�`��g�s���ouM�����x�
��*(�|g޴�oR�x�|�uӁ�$?U�#d�c1��U��9z��n`7p�SQ'=��v"iJE�i���0f*y�	t'�Ӝ�Ѐ��pft������͛6d�*��x�vr��j5��o�E�ɛE-7��,��\�Q�ĺY~���-@����U*ZK�xEw��B�J��"�f�v����#7�;���S��E�y�УĻ{%��ە���z2�<��]e��������+g��C̆{��za�Þ��䰚�?��п�*���2�"��/Uɵ���\���L��χ���.B-��f1�J��!�-�U���,`�SA�n�(�L }a���$Q�҇M��k3�cg������D��IQ�E��Pd��RXG��E�Yv��j�H�;g�$�|6�L{#�<	��͒v̂��o�8�,㿯�;٭x������x����7�-��r�gWf��3�Y��7(n�����ZGLj#~	���@H{<ŽA�K�>��~\��4*����4-}zh��Bd����E�@� ���KWd��+i��4y���3������$IN����T5^�A���J�2�"D4/���z����u����,npT-���h�$%��~�(�]/�c�_v�p�G&����l7��ݜ�U�c���ʫE��5+C�u��4��Q�R�M�5�_/OH���e��z���SU��|m����U��?2��6�c<3K��t[�`c �j**(��e>jݗ��wh@���������m�#��gN)
�AU߈^S\Mۓ�	J�[�L�|�.9��l�b��y�6�=gyxif��=v�^�l����s�-����j���)dњxi�R>�E<��N�c�_�Ig��znCU6j-��nl��@I��Q�whi��󁻵S�ჲ{��~��L.Pһ��]��3�H�F�W��O�޵�!�ao�{�`G8W85kV��<�h���q+C:o����!�ztuc�Ȥ����ȝ�k��tCM��	Բ�;)�Ymߢhy?��-�^����������^������֕� �[4��$A�ʳF�ck�U�f[~��L��ԠÄکnI����ޡ�G�)�"���59fm���&U�@��s�	;]���"DhE����?9�R�E��fN�\���� ��YE�
|= UK�嫢�->cC�X�$��1P�<�{[al(x�d�sn��$��ٷņ����a���آ�Kۂa��v�Bs�N�c��*���Ǖѕ�Z�Icp?�QFs��'���o^�RjaK^���&�W�h�8#0x�/�$C�[��nG@V��0� ���AX]V�T�,�֦����		<��D�s}^��qN�/t�^*�7���VN�itSS_èz�cF��� ]4i�O�+�t�fls1��u��|�Arڮ[��aJN ���?�z�P3l�:��0�`qS�KҰῲ��̫Ý�UO�Y���.��V� �7��۪�!���F���ؕ-���=/|��y���^R�D���]�`��`(�-N;�ؖm�.�y
َw�`_��b�9�h��d:o{����a�m����@	߳�G�Դ�T��+?����c(Aڕ<�l�'�5��2ON6+�����LP�?�UoZo1�&D��.���,@R� ��:����7�Y�x�� ���ż�`�/yn$�}f�Z��0+��ܝF.�t��/���S��V�@��"���G0�[)`�����6k��إ�d�r�+(���\������(g�������Be��$iL]wj�}&��kmt�2.�ه՜Ԏ}����q�p���"ތ�yzY��=mJ��~�㦵��<B��(a�o*�E>U|� ���qB^��"�p�42����k*sا�9\�W�"�X�W-�_���h�?�7>1"]�r��7UG�~e�y�� 7B;G���K��&.�]�](:��d\C��Z`,��Ǒ�j�S�B����jw�4`eu��k��c8���n�C��_��gKSJ G|�T�;3����
��K=��Uc<��ڼ��U@��^|v�,���=�,m8������j���F��-��vl\HF���$�bt�wk���(�4�_2��V��"4y��1���ITX���ǟxZ�fb��[FI��Y�~q\x8 Z�]"�@����17��U/�bM
�\�UY���f��NhJ���2Oq�����M])�t#kՇ73��qH�V�
�:т�KHqA����d��ZB�/�rh�>��`VG�<�f�P��]�ɭ�|\�M~��|!���c�ND\��u�� �C�&��+h6$֕�a�U��Oj�/k*��D�������6���!��;rn�(�P�w]ʓM����+T��N�#�Jb�\Q���6�iiE�O)a��2V�Q���8:GҌ�(  ����$�����fD9mo��J�:t��zϯ�K��w1�s���V<�R �����5�A��=��V-ziX1d;ڱ�{�cʅ�� �Snl�C�F�1��t�Ҙ�]�8����_mu]uLw�5=���G(���#i�	���ʮ���� ��u|{nЋ�/����{F ������9���v���X[/���E�x�X������FA�8��\L�D�!3y�\��V���v`FB�{��A)�;J��6��oZ¿('�C�X�*��Y�+�AW^F����BF8��4��8�X��i����8u���tR��m�r4C�s~�����i¤f���4�l���%Om����v�3�*��.�P2�D�; j�Mі��7]�0��~ei9ZȲWaB㵍��_�Y3X��4��fV��E�
8s	p/M��o��5�!��M3XR�Ï���(����_(&�m�9�'��Vt}�T��0�;BԿ�Z���Yjb���]��cՁ���l����B�P5R�@���͎{`�.{ԑ�bc�}��#��/�
�r�y�L+�|�UE`���~{�0�q��S�)1�V�ˤ��9-�*݀Qa������BB��%¸��o�L�t����P\�o֎?Q����H����3<�·��f�b8v��j�"i<DOpdr��耣(���*ICt���
���X�qԜ�k|$?�9����¢�".h�̵?��j�Ƽ���/gb������R�I��^I�^�Nkp�_7:aŧ[r;㻝xS�j��9~Ԕ9inny$B�������cV8�N7wQ��w>9k=�53�G�z�%�҈�����\� =b�pB�2���WU��m��P������i	��J>$v
Y����y����	<$ �����^�a(�[�&2{������A֌:[�T[�����k��I��ⷕ6!z�;��a�0}�x�:�xe||A�i*�\	�+��>�cifS>�ڸ�l��]�$C�'H'_9AB�6��E��m%��Q����~�0�+�?�Qn�\ӌ�ܙi�b���Θ�2C&|�B��(IRn�D���t��D��ג6��K�u�`i(�"p��C�/UX�E�ի.mS�;��
��W[mZ��lFdҳJ�KT �6�rW�渱y?y�;Tx�?�
\n��v��,j������7��·v��9�G؇�@]מ?�s��=��T>�nY�ބ"ߍ�*'9�_e(㙂 O	�g�&����0y~׽i���(�译N�
��_F��G�@,�c�qݤ�?{R���3�+�H���V�ÛY�0�y��'^�]	P���q[c"I�d�k�J\�#���M��~M~��L�҆���W��K~I�p�/�J���C �(������j�X�vHzH�6�,�[C�U�t>6n;]�%�ڴ��[�/{͘:��e
��.^��1�(=��-�9�Hs�#�Y������%���+>�"M��R�e��.�WL����Oo���nqEh��Sgn}��Sm�b�����.�vD��=(����T/}8�^�y�h!|M�SBD��� /�J�JBt��'Θ�[�[����%7����˨���hq/���l�R�{.X,���5�g�b�U��k>��#��3���p�@[�i�"?�|��4��=<{��U�GY�]UËuS7={&Cl���	E!�w��T'�M1�S�m9LO�����h�ag�kw}�9�!�ɔY&��E2��?�_�OQ�h�/T�f��r���d�i������Z����)�9�oI��!@䇊���F��k�4t%���.S�ɴQU�����[��菧4v�<~½2N/�� ��V~�h*z���D� Ej��%���jży������b]�C���S�V�ꉕ��k�caz"nP�xlA��мr8.d�)�~����]p^?�E���[oic�0��<�W���8'Wko���Q��pK�ȓҴ�9�;��G��ls�eM��[W�C��OBn����K���D�d"�lR�=h�@�Q����A�ɍ�m�5�'�(�h�':&�G!!���řT���X�u�e@CԵ�R5�����c�)��i1���!	`� �"��ټ;�̢a@~-�����	I8$��ƚ�����:���(>�a�c��F8Gnf��jM�����_o���4Dt��g�~N�y%��{:f
AeƮ#���.�Yל	�ϑ����[�u���庰qe�#��(��*mΈ���4�C�=��׭n�Y�x�����<a@��>ض��\�9�pΏ4�R�\f���;8d���	X�<�"���
�n�kN`��ï!!4��~g#�p]cP�@!6����#��e��48V!�#WާM~zϛ5;&�S�| ��J؅&�Xk�L���#6S������֊|$�p��������c�ls8eD�C�]am�]���/=�Y5]�.r�#QPz��F����W��0�i�/<�.�on�"��1��}�z��ζ�G`[��𪙧��A>mI�����ÿ���5�?�v�
���ޔ5>vgtp�_�d�V�,�6%� �z�0�Ҏ&���`��sy��&�L�2c3M��E�9��-?$ӏ}�
�'�GB-��/k�-��-xٛF<�^�nh�e���n�ueāF��"��*׀���,�}�(7[qɅ��Zb[����Qh��yg���)��w׭���x^��;T:|�w� �2�L}�gP�Z�w�0w�y&ו��DC��J\e~�U UH���%C܁{ot�}��r��3�z���m)sH*b{Kat�� l��mzm�z�Z޸;3�a?L�(>	��Z<#&�,'�G��8�;���^�9"7�3O�����R�Et�E]���2����;N��
:0<����@3c���ΘÅ� \-`��2�;5�L�Ǖ�F%R`r6s���M����;��])�|�Zzi!J0�aú�+� ��2����%�|�;b2Y�6�M;�]IQ�}��,տ��aSA�#���g걁!r3Oi�G�6�8j��v	�o�r@.A����,8���#{}�m�(����e��7����f_��X�uNLr�]SF��>ʐ�v.����<�%8{�3
%��R�Teh7�^�!��p͜s�`���a��!��8w�16I���
�3)������@��sN��>΢=ll$r~��98���J�x���!��0%�}�AD�\����ownb1t��ɬ "D��J�#ǧ������@u*<�H�Å*@�.
��L6Mc��:�"GО�)~C�>g��Շ��h��4�P���ܑ'd~��[�V��kKa�d�T���X?��ުEf;�RsD�T��gr�5�MH�<&a��^G޿��-cЦ���tCΛ<�,�QCCi�ˆ���_h�P�>���0�KV���մ��`�~)kZn��A����Rlq���V_9E=ː��2N_]B��BH��� ^j�&(N�8��5ۢ��JU�L�
`t��$�ި��lș����� �lU�e�b�Z&W�ܮ�l�$\μX�"k�`rx)���ϻC-[IYy�u�d>�;�i*�g�
�7E�� �)���`��i�(~����q(�a���Z�-r��l;T�Vv�5���6�����	ؼӬF����d�u��1-k����[q���2( �:{�S'kHT�ᦜ�*-��0��������t���W+H<e�q����7c��9��m��nl���Jf������?���i	������5��b���5�n�m��S�KB�;�e]��O���6q=�f<��c
i�"�b�X�-� ��{���>��}g.n���(>ý��"������/<�2�;��w�7��U�I�;~�B��C��3�_���X�6�{\n+�O.����ɸ����XI� ��L�10C.���S(���eiv��d��9���]V��Ks�����[PE�Ywkl��9����q%�w�R.��<Y(�P�@�ٝ�.�M�qOa^�Un��l�k��N���F�t�l��=`9�sbtN���^Hq�ߙ�tV4��=Y%Wp�~��$
�֝�흼�G�Dw���#��Y�����'cx� �Y�;`�frbBn��8-�U�X7t�|~�~���݉�LN�0c͸S/��<��V	�i���,u��
�p�ʫ �l�yQsu*_ w`q,@wc�`uS_|�a5A�h�w��!t���ݏ3�)�������C�w�%� 'đm�i�8�S��0}5��RG4�\dL���%���Ik���B�L�Z�$����8>O�-q�Z�'�s�"G@�o�s����<>���ЅYv�F�έ�~����H��{&�UdHSQ+�1*!+xK���f��J�sV*SQ��}��w ��)� �W�/��Z㣝'�\��f��D��Y�u�G�BJ	�pPK�vr=��~U��[3"���h�$���MsٵHp˳���&`Y�E�W���Z,x.��w"*��)�d�i9�ͯt��=�5�����ػ3������buy�'-�b;^����Њ��Fo��Z��>X�7bw����I�OQ�i�꿙�rg*��^O-��KlOV���'ƾ�<0���KZC��.hR�����j²Jx=T�"~s]b�b�L�a�-�o����C_�b&V�3�Sl�@ ��d)	X
�(���)���v��Q����h��Q��u0�WI�;����,�Ma��w�t���]9�Z��v��GL8Kv�ƀj]�31[�
'�[{Àn1��a��1��_�`ؽ��o�H2�U������$%lHo( m�<��K���G �����1�TT�*!�w��Tp��r-&��S['�F�`>��w/�)���
sw��|���dp�\��ZZZ�[@<��F/(��J���[�i���]K�*3E0��A"~,�}!0
j~�[L_���TeՊ��6vDEt:d!�h"��<W�W�!�Y�X���9��������}J[�v��bq4A��r��')>_��xW6������cI�t�o*��x��i�������O�����t�m\DC �n��,ݘ���uug�A�:/�af��6��>9��顓���aLG� �l��t�3�c��030��u	�В iz"+�a~ �V���3��:��y��%3�H�V�����(�5]Jz�Q�'θ�uKN�����T�zn�(k���c�0!�4��$�~ۙ3x�c�D�cVnPd�͖�S�8�xWM��48dN���4=g
�5�M��s"�G�S�8w�B��__\ߦ�\i��싡:`��?�����y	Wy�<��a����Ƌ����X�"!��1��[״��}z��,�,�Հ6ZR��~���羃 Y�� ɛ񅎽k� �D�-J�]�[��X�л�=����y��-�(3�TOXP��Ё��@��S�1�mNZ�ƍh�-��r�+�����G�6��Ә����j��\�{��mZ�.��C���uOE��WL�и�EԊ����=ř�䠥$4N�	��ޅ��Ӟm�� �=zA������(�w�7�t�h�fב>���f�0����!f�X}�UE��p1k���h��)��X�����"���a�
tJx��֥�������7����˼|��=�#i�>rF� V�.��+�fXY�����M�|��g��נQU.�p�Z�|��)u�75��?���8W�)���C0�x�Ҿ��q�s�IR��NQ�0��@����x�� ���^�������7��/���/�Re^��a�bg��;��6�J=?�L�q�!7��q��K"��K���u��̹�Yz���r�S�V4P����#������g�?At��&;�;˻�k��e�H�P9zGe��X�}v-l��A�a)��Ӻ(]�:PD@��!Rr�M%y$�4�7�9L�k7���r��Y��X�*� �J��q"��u��3�Q1[4��h��0�!���H�]�F�c=z�wM2�l�j�x����u[\��-��*�YQG47�bن��\���Nڈ6a߷=Qrו7�'�ԕ1M!jX����ЮtSH��2Z��T��?x�a+���$0�U�z�`Pq����ucAwYcߜ�ܙ�n�{�Sp�G�� Z�L��ܞ�Z�~��"��f�`��o=��LxY:qϕ�n��=����(�W�����w�>�?J�L����̍0����������jѧ׬�m��GXp��mmP�&�=�������ke4�z\�!��JB��ȓ��ު���߁LF%�(8 S'F�%V:����Җ�i����*����Mp8��"���9��Acn~�Q�MX�>C�F�7��G|�����Q�r�W����ige�w��ߵ�p�]����Bᛤ�#�m�/�5�e+�}e��Qd#��oMq�cc��+aNW����ϝ�������0� �}��x�]�e_4�3%���>f$��v�SIB��d�i�͂J��y�ͣI,I�W���7�]�dYY��l6A"=Y��T���x��r�t����{�=���AY`û+�"�?�`|n���������(���%�L�s.����yf�Z�
�P��\,��@��� ᰾��� ţ?��F��bd5	�7���)�1��-UE�1��;��ӫ#22rjd���'��)L��VMn9�`�q��%e�Ĕ��5]�@��+��}%��jR,�p�E�5�x�Z٣���z��,X�Kx��>����=l�5M;���GDs$���;�}=�-��IV^ǜ�yI8K��:�ֳQ����?�^���� ����x�Z�)/yvPH�G�M��U��T��d�	80G��2��(Д�=�a|���U�- ^���y�έ��}���}mP�K���<����~~o�=B�$o�O�R��~��ݧ>(�,G�?<�:f���T� ��Zр���\
%Z�l|F��Kvc���-�3��=�'f*���j"m�6��@Y���	lQ�������m
ۅ1:��R5>I����ńj��P��-0�d��kPQ��6��UEv�m��bc�i ��"���ːQH�Sz���%��j;�"��U�q��>D�y�̭a���K�xr=SqZ0<_��qc�z���!>�s1�`"3�ɻm�m��H9ЙVu�9������S��&��:D�(����Oz{�.�mSv�����I^�у�1J|����������G��w�'��x�5�SPJ���̯�b'O�_�y>"�Y,��"��?��{r�6�@ ��kd���i+�T!���f$A��#�5��곷-{w�Oc�)�|�zQr� ݢG���FfK*�h�݀�|��?~]�S˴3ZD��͂�)�^��^k �h��'zS`��s��s����$�^�PZ�T�S��f� �c������c���@�cY�g�A������9�N��7�W�;�`Q�k�Q�X����M��x˃�|�Q`�������ұ��K��|��ǫ��Tz+`t�{qE1W�����p��b�4����+�x�6!KYu��9�I�R=��o��)��wnwuzmK��� j?v�9��:5I�Ǹ(��▊�E�O���)�#֯ґW;�R5��X�����Mm6LMg���k>1I���
Nv��mz�Z>�ׯ#�R���O����~��d���I
�vOfuuxr��T3Y�m��FyQ=�IR4&��}��#$hR�ߒo�|NɥX�I��=��E�L@+D�WH��sr�(Ӵr@bSO7�RO�ᙅ�R��L�F[��-Fv ��3�ž�V�2�=�A��ƒ遒��I����I�}bE�:����L�d)�?Y�0�W�����>#�+�%W�frj�w6���� wC	$�L�����?�N�U��E�ڦ? �.㭹k�;�^H�ȃ [kq)�~V>'�� �iG��,�4i�J���P���P7�R�z�řQ	��y�Q);�4]Zd�Z���Ϋ����̧H�e�4����5�+�Asp�����n�7*�A+_8C`�xk�czэPs�u����m��~a �w/ac��R������ć����Z��[�J��c�^���<^�KI\,S��l_�МU?�����>c��<�ֳ��9��r�9�Ŗ���{:Vo���EJ�L+�	Ҕ�H9������z�%�����|&i���]\�6��e�d��-*d�s�GH���c��O˕Y	�I��§+M�#��D��|C��,���B
I��L/8�$���`����V�0N�C蓆���G!:�H��r�������'�F�WM�TKl��^`��%̻e�QZfބǻ:M�E���~B4����,����~g6�o��=����f�˨7q�j��u��z����,k/����Ŀ���d�q����i�m� o}�����z���n6m�,�h��T%����N�z���m�;��	)�I�q�H�2J���r\��	<�}q��%e�o�Pdw��e�����#$�����'���@�ٔ�o��r�S���Xjx���e�˩4�VԿ�(�[�Ӓq;��%���Pp���xG�wT#U�HU��5��V�8�۶�k؁��mbs���AKC���O�Cd�eW*ջ�I&�YH���6��L����F�3zF[�W���'6JW�	��7E�~s��AĂ�����Դ�:����~��򤲚�G���� �
�DO�	g�2.�.P�R7�M	���Y�x�e�HfϿ~�W��0jdsu�}� Z�s)J:�ѰU���,Pe�����+��Pvq�m���Ʊ3��S�0[�H��s.5�U�c�_O.#��N�ROj�+K��æ8��m��u�-ֺ}��Ը�o.�{Ơ6���T�X	T�a���?ćۺ���ι�bO�ͶT���'p��p���d�(V���۱u��3���9�6��C��qE��
.����φ]���9f̐I��+a�����V;E,�sP�jg@�Ƿ[$,�I�NS8�O���x�ܩ"����'�ڔ������5�#@�,��<��dc�vO�:�[�?�k}�q-���0ѯv$a;�\�{�Rs"�C�Y�� t��+P���W�Z�f����_�� �&����R,��n4X[�7Й�zqF�M��M�����󑠘U�n���l�+���_�C�&?q�c�"(`¥���ř�Mp(� �~�u���k�N��.P�����b9	�Rb� ���ۍ+����+�ԑ|M��$t�B��"�����vO���#F8O>T����"��l��3X�Zj�� `�8�$�;�_�<8��t4rb�� ��*���y1��'�%�慨��Eh� J�V��1*<��柯���o��J�j]�Kl��Ժ�Pߵo��>��B��Ճ���̑�ԏrB��zC2l��o5���t���P�>�_peeX�A���X��a��f$��뀆tZ�p}]�+q%�0��=5d��8S�d�DdO�K����UV.$A#$��Rq��z�x���ϝK��9,FEuHς���du�o�����,);	�.8��]�h��	��Cp�V���U���m���}��v�&���J%�z����_k�_�G��3�P��4�5ɞ��sl2��ݶ�n�g�l���5kb��,=_`���az&8��֑z\�'Y�xA�����p�����%C'e��ɳ�D�F� ��&��
��,H7( ��.�Bw(��]��E�訐�������\�3�_��T��qG�AE
���5���]��NFr�0H`f�����h>�b�_�|^��d�^H����!t�B�́ӛx�d���� ��V��s �z�0�YZ�#�9��d�`�@l�2M`H���^��V� pn`�;0�ܾ��
W+�&�$^Rῶ���vnZ��v�u���:��O��.P?����^Vh2g���xK�a]�2}��􂴭����[\j &�`�R��^�/�9i�'z�����}��Ya�;��HfxDs|g�|.�� }���=ˌ��aZ��`����Cz4GK�r�O��tu��SOy����B�����\���Q�k6z��s�8�|��������d�)_��3!m���rBЃg�xH�l���4�4f��Q�q�i��t�K���+}��b��6Z�M�#/E�O�t��ed�k��ð�޲'(������7�vZ�iP�����׻a3�ל��B���^���К�?������m�V �4��UW4�� s�}�[X�
�3]��D����qQN콆Ν v�E��C�X�{(wZ��lq\�W��sA�U�u#o��=#}�͐+�Ò��k��L��No��ѵ\�ѣ��r2-��*d�b���6�����N�^F����)�7�8=����F��Lȿ��tti!��ݴ�������{)�;B��ב�\R@	2��w�n�P����o*�d�=����_kw���0���5zb0���"H�E����uk0�OL�of��ԋ��^v\�h�c$�^[i[ ��mxWu)������s������YVr�(g �{O��z�l�/����Ĝ�����H�3\��\��7��@����ɓf�t�Гt��j>.-�>o&
NTץ�4AY
��+2_��z��r�z�EZs.��6��2�[����Lð�2�3��ˆ��^i��/р��%2��p�m�˟�ԛo���) ��0��T6j��&�d�Q��;�"�e��	�c#�.�{
��]�5���*����O�o$�i=)�`g�|c���SXz}4�|\[t�܉��-f)N}f?1V$�����$��,�W^�1��W���;�F�	�2�V1�k���lR��||����9>�n���vu���_:��~��n@��a��;������d.�P1¾[��\j��K�B��M2���G(�0�P>�̭��R�3g����}�Xi�
;#�o�$�E�`Yz��B�1�h�]�%���/���{w��y�ї�C|���'_�P��U[0y�,:Ԯß��l��61���6�ٞ����o=8i@���:����Ԡ���T���S�>֪QFLʱ�	�2c�qǙ����`����
��Q�亻Xf����;�>�vy���f�28i�JS�#�kt����1r����i���=�T�("(�h�1��	S�L6��r?�CHX���M=�� �|x����GJ�$�����t?/���x�Q���^Ɠ�yYB2U�my�&�"�p�j���"1�
��G��`3�>A�+"Bsn����V�&�XY�Y:�N���z�+�p� YX��!�R�%^�F1��ۯ[��Ȓ︀r|f��v�󭇚X����wH�Ԏ{?�g{�++��w�	���_��q����O�[��������!��c����al!�{֩u�����U��k��ecQ�9)MR���g�eN����Hx�5��]�N ���~5�DpE@�,xg{�`R���4�Q;�8Z�w����
�]n�����O����d�1L�9)̠�Y���;�Yr�^�B��c�T�"�׬�~������'VH�P������)GZ$��}*|H��wA�g�)22�T��b��r�{�2�ef�Zc	%�p�!��4�W����Q�?5�����F"�$n`�c�'����_�!V��,O)�{]��w3R� ��9B�_@$�>�΃���z2oR&�pT�Z���,�H�4���F�E�����9,���#�O"<x�$F��.����		�P>7K���}��i�#�������\��"��[SjE4�����)^)��*��	�*��r��_��O� L���ny���V�����@�_R�"�r���\����C�貹���Rȑm�|�|M�!�D_J����t�]�+�2��u�Q�\fߓ,qow����!!�c%��]��B�2%i�x�لzp���zA�	[��ě�R�7ƙ�'�;�׮OG����6s�lfMq�X���Q��n�_epv����T�3�f���+v��5^��¿*1���n��lw�l,��,��Ü�D����t�z\}6xK��Z��(�u=�T?���d>� 96��v�8���N�=ۼq�织ʣ|�cN!�w�3#�m���J�̈́���3x/� fk�ه%|*鞔�1���.I/9�r���H��ۓ�\^��QB�cݕ���M�Ҡ�`^��P��X�z߇-&�����TP|�8)->kAs�,R�ܮ�u�{Ԃ�?�=#DR�YH�R	�t���U	�����KU��[̔��D�p��R����u�����.�oq�����j���.侇\���^=|�o�����8Hy�(:�I�.��ʏٸ��a-���Ht�)4j�������z�ʸS����3��O~\��P����*�M�k"�D���]�/��g�0�l�����%sAҼ�Hy_�R
��=J��gyv6父�)A>Q�]�^D�����p2'�`�wƩ��I;ah�<��^�n�:	���S �j�H3�F��,��A%�d{���y�׳��{~֨>|ƸjЫ<];v�B'K��_;y'n#[G�&�ͥ$��)��~�:��O��pC�Q4�x��x%��3|�:5���/�f_4��k|���T�2�$c�k�\��fP�}_�}�(X���\�����~��(5q��,��)�J4oe2�q��߮��sz(�p��X�9<��R*��.�� U�(p"�Fid:3*�	�|ʍ�谙�Ρ/&t�>U����,~Ә�:�I�� ��j�q:c�h��W���͛9�y��u����>?��PV,W���,�����x�N��@����
䅘��d�zh��$Ut�Op�e��ATS)��E\죬�ȣ�����qBT���n���}��k���$)#b�%!��fC�n�v���2g�  K�q��F��!�/(fi�����\�M�g���n������>!����Y��/�ǐ���s0�+a��օӏ&�2l�v?���$Lp1Ձ3t��s=��7�J.)g0�4�`&����^_�|I`Z�@����n`�AYx^��J&;bT���,�~�	ɐ.����_�}̦��.�Y�� ik�~�*?m�ާ;�˥�{��ڸ����ѺBN���߻�%�����e���lN�������u�A\�4���9����!;���dcG-#e�SJ��E̗�~9�^�i���_J�g<���2<鍒���R4�JW�Ɍnư��"�e�P����
��'��So�<�T�as��[��^���ߊB^��i(��&�J�nQ��{���	�C5H��;�@}uf�K���y˳���:pՂ�d�w�tU���kmo�w���M��?�a��Z����	Y�����S�Y{3��.e�B�,J�[��v&�i�GxC��%�@�+�P������3Z���+��"0I�_����Q\�y��ypOgH-m�S�"��ݸ�7r+����+7@�b�'ѿݻC�A�4 �8����.�ð��	%S��0x������P��nV~�^.q����a���(��h�5�uĨ�+��.�;&�jF���VB����0+"��i�2nM�l%�ޑ|��y���I��p��3=u��� ��� �fe����������l������$�j�xC%F���4P"iq��G1���z�mgTs9�󺉯�P�m�l��π�NH(�ǲ�s���l���+�,㚶�D��jq�s1 �I��-s[F�-g!�q����h�BO�D���B��IX��)�I�ر*��<O�ƛ��O���BsS�\�c'}kh�9����I޲�.�Gع�������Z��J�b��rH�n��ZT�\�r�F�kr���7��m��� ��P�U/�����']��[E�� �����0ֺOy<�V��8r��L	x�s�;�m���8e� ����h�\&b�o�#{Tw��zl�m�X�>5'���0�
�s��$ ����h[�r�)08.��fo�Y|���|�!�l�d8jd�z�6`�"�7�>���7t~� �c'Q����_/vR�'�vO�]�$��ċz� ����}s@OA.{J�9V}x�;��j�fg�h2&c��SS'�}�.�6�̫k{�Ay���yL(~�K�g���V�mLY��_?I�R�27
�*9��G������&b�a���|�SbYix�l��c��L4��|F�4��Eڌb_O�+���Y%cַ�N�JtG��؉��9,34z�]ɉ_?��D%��dpy��ѻQE�6'9O�O�Ӥ<<���nB@#�	/�,�`��G�����~n6�v����y
:�Ō������z����m-7\��4 r�0�Ŋ9=\+�%���f4���M�w�	�cE�ʮ���)���#��.�3h�A�r���,,K��2AЪBG_v��kScH"�ׂ'б�Zٞ��
Y�<��ŗ芆��(�BU��M
pZ�՟������X�%��a�VKf8��D��E��*k��v��7,�?���z#�1�g�h4���Ixl��0�g/Y��[ n�Ċ�Y�Bv�B��+���Jo�������m<��>A7,`���sMʔ�-���/N�gQ�X�#�H��S`f3]f�rH�ُ��B������R�D ��nT������^����92�\4��F57�!���q�zS?�S;�n���%��֜:�X���ZI��ϳ��fm�[���j��x��%1�ԑKy0���Dg}EjK�I��6Ҵ>t��C=��hJ�P�W�$�*n���Ӥ>��P9I��sM�E����7�X|.������KNP��x�4iMj�5F��%R��R7<&Z0�pʈ� ���;o���;mf��NK���>.DB_H�&.�s�z��~F˹�ѕ�\.�ɹ/���S��7,0Ѯ��U:~� d�$���%�t��%(�չ۾��v&����F7�z��F���	� �`���s)[�a�NC(>F��;� ������!r��jJ�b{ԗ ǀ�1�_3�L����G��U���	��qE/�����K��ot��)�4y]�!��}�&�t����U�����"��Wd�,���5�H[5K���O�#��D��B���]�;>�	�'�vz��)�"0
0Aٽ�~֦�ɋ`"Ig��<�3O[���r� �حY��?�q��njѲk_ܪ���~��_��ҚJ#x�5�#���*�����u*]W���T�/�`�zȥ��{���&%�:����Z��(�I����ҭz��b�윰�&^�*�'��1	��lN�ĀF&&��MXY8W5�$�eby�"��KA�y vU*��m5iE�1|���5��k�n���� �e�*(��u�8�����k���7g:��d�)�m�?X.�E&JR����:4?e���;����N������їAKS@03��*䡾.t�ڤn�8(w�Z�pKa��?*+�W�r)>5���:���u@��������B����_�(�����*D�(a��B��#���骣
bs�N��I���E��&�Ȝx 'W�kSQ�#��շ>/h�"�杖�?`����^�ŧq��¢|Ү�.;P8O��<K��&�W�h���e��)����Q��@n@��_�A����,�D�ƞ��Į�lM�7�������%yt���߹ĉ�0,�*��uC͡�/_���"��g�k�������cT��<�dJ�:�^���aE�� /�x�s�����wf�`�c��5
l9�=��B�zకH���ؒ��G<����}�';j�4��%N8.?���x����-�&X�N:��~�d�$��IV#O]O�N�	ll�r����iܫ�g�n}�O��3�7#�&���k(� ���~t�����Kqu��C?�KG\ʤЈ��p�N�EJ��(�`������moe��8>@�j�y������&
e�A\9,,~ߐ%��O����4�@&��o��"�n&�� ä���\��e�$�Kj~�7��B�\.�e�s�jD_Ss�*�)K�f�	��j�7	�m��}b0o`h!x�}R}xz�����5���U!04���!�&y�I9�P����S/�ȋ&,��=�XYt�]�]���qCo)�kI1,�{k�����#DQ��-܃N�C��7k�.��߸kG��H�՞P*�c��R�3Ƈb��`N]�ux�:_��u�c0Vɫ����`��f%��&  ���U�C����`�Fsҫ�(��|>��m6|]@��M)����ʹ��A������u��J?Y��m��b��W�^�޷�a�����R~*��g���)<��0n�J@@��{�3N˒<�Zv�\8�Ĕ�-x��z��2���=4�����Cj@�t�8(Q����#ݵA�5��j ԕ$^�����(�p��뤷����H�mH�+k�����鉴i��I�1�X���<�����s��_���H���H�F�!v��{�|Ũkm���6��2�px232�a����5y���������'�;�����7�t�C��@b��1E^����[�e���O3��~��.hw	v|�y���� �3T6#� ��mW����<��ajw���z�?��~n�H�#���U�{��+�����T���e��f&��31��{s���J10�P'FW&N�P��.?PXH<:܄�yĚz537��ʍ�jH1n�L�����S���q���K63�2������F�]�~`�*I�w���Bj�P�+�@i��}���zן�l���Cd�L��&����@H��):����E¤�ɯc��ރ���I��gMho0-n����CE��D��&A��5eO����r�P�yw� �f;t�jųQd�}H4�+�W�!H�(oƍc�oiu����C#�%h�t�Gd�?A���@����$?��)v6*J��XE-$؞ŗ�k��_��/�P�K�,X�BYa{��ņWli�ݴ��{>�b��P0��O���Py
�4E��!d�_�T���|�E��d�����
�<
�'�4mM�3���
[2?[t����^ZBpӷ-W�*��8�)A]L�m������V0����B����25e���6}�-ϋ����!q#dت�8�]Ć�VM�ow[ׯ���KT�1ph��z��(�[5U�ՠ��]�S�f�t��6(߹$���a�;F|�՟]����ΆB��aJ\�$������}�4G.T[��Ȳ���
�2��K��;i���w���\�M�2ߗ؋�vo#>.�I9{��N�35a؊x�,e���G8*�ë��([��0�#($7�4�{?��(b���m����U=�ܫ������x��L��8��}H�?+^�G���W�g[񇁍��B7�x���\Q#t��lp����" ~��@�EO؜�Si���㯆ő&�&Y�s|���s-:��I��@ �oF?Ȋ퐺G	)�Vf(a��Ϳ�	��L	EF�.f	�x�=>�0�\!���Y�7���/�m��t2�i��I�$ww[2�j<���l��T��s����7��ԟ���M���%r�bY�iʀO];���Xؔ޴�'��@� �2�NÎ�Y[u9Z'��ܐ�q�B"�L��&��LQ���|�����u�kP6�b�1�#��e��VUk-׀\֓`�(L��ZF`���a�麂�f��-h����fk���[x����3�������%'	 �[a�큵[n$?~���Y���;y+�B[��_��y���PXK�r0���{��*��3��JX.�<��;2*�����_{e|���9U�î -���:{�������1����fECS�����͌`�z�ߌ����{^{������H �^o2��������^����|�W0�M�jߖ#��
K�Hٍ:�3�Y�~�x1T"�w����*���j���q�r��XH��Aâ�uS�4<�]7s���g�Pe*ħ�t4��N\ ������|s�J��V��<{w-hf����&mT@=H�qT�1��t����$$D������"~#�*V�~���m�x�/^�&+U��`3�f7=�ko�����'R<I�0<�b�\���2}7Z�Dd������aT�c�z/�܋���RT�̜W��t��>X5f����c΢�Pf�i�f8�W.���C�Bq ���4۝�lJ&�r��T{�=���q�ϢQ��g��K�q��-0E�Pl�Wi�?��>n+�BL��*�Ok+@�!U���=�V��K�31��\ϚI\"�$�x��t����S<LM�.���c�'�6�8'@�cq}�U���e��Ǚ40��59_8��O�e�l.�q&K�i�tp�m�j��� ���Hז��e`��J'��mtଲ��2�'� �ّ	�K�96]L~��b	�`uf��u�LePhե�\��-����^���t�[����ADZ������d�{�^�L�A)!�r/���
�e��D8,d�P��bM��D��wqH��y� ��Ɲ�rN�����F睖A��=���c)�b-(o�;+�j��=ܮ{��Ϝ�z{`�و�͛UVna��|��3'����x��]����x��$��A.�[��?M��#��h�J\	��AHƍ��F���� �g�0v�������	�h��I�����D[Ǵ{$��x�Q}*+�T%M՚0QeU�l���:�w�uU<ؖK�B%�^�R��e&؄)�_M�~?���t������q<`�ҒPe�*���y�@��x����q�i�����y C�Q�s+>��Y�m��K��C�?�n���dtB$������N���M�6�ه�	��V����a��ԳEb1����6[T+�	6��R�t��ʑWJ¸��G?�����A!Ԛ��5�S/J���D�0�Y�.���-��h;.K�6o9X���"��{&e����Y��+�B#x	^�&񼿱ݦ��]��� [��P�M'���u0n���A���ѫ�}ճ�"�Gٝ׏�eƌ6�B%ܾ:�)ϟ,e�lP���x�TN*׹��r	 "�=V�n:q9�)b����#y�Tj�{�L�I,��b׀i�^�����u�׬+���&ս���`����7�E� ���a ���B�Vy��3!D6{y�F�-f���O��{��c+su��HA�S�C�V2ƣ��î7/uP��.v� C��6�U�:��ԣ�l��F�Ԓ��A0�l ��OwnT2
�-����*�+9�hф.�&�3�~{�Y/�����_l�>�<R!�^8\��z�6p�/��������n@�=A�r���¨W��G^.��c�}�mO>�|#ghI`%M?e[A�c��I�R��r��P���8��M}��7��l|hzz��l��=bҲ��4������"�q��=�����F1�n���_[Mr n��P�h�c$Z������p�{�Q��̶��G����0M5j`��w�QM67؀�'�\}�K�~=��D�n����W��~tf]�Oy��\��_��o��5a�e�U5P_ �,�����J⍏��o z��Y��4�qN��
�P�,Ѻ[͙x��������Z$�qX3+�9\	Bw�s�������f���5x�I���?��|ܨ��G��g���B�T7E�Uޤڊ�L����׻�r|��>�i�&��OsDIF�(�yQ�Hfs���V9QӢ����w��y�����|u��"�?>b�e9Dk�}�z�p˚V���}����Dd�x1|�2����rG����_tB2�~-瓟^%��%_$�;�by��#E�6kg��?m�� 0v���OS`yeV��|y$�1��Rz�-�M����4=�p5��)Uw��Y(�;�~q���؅;���X��b���۠ˤ���RkΓRq�_K�RÆ^e�c]+G�i���\�RX�IH�+?=�-e=����"�"F{��x;�#�r=��zٮ�ǾW�(��p4��m�y���Q�A�!I�d7˻۽�+�_쿱�m��}Թ��)��/��1��mBi����#`]|���U�Q?����L<���Q�;Tء`���+p�@�[���~�[#xE�@�PR�j�E;Eq���;��-\u 3~����~�E��u����/�381mPfAV�aF�Ry|�maي.�S�����/��5}��0,��Z���0�LC%��X����5�ث�to�����Q+�I�F�fj�?{ţ��O��#C|_��i���u��P����&�d��)������!!�7���P1!��g�s�������4��	��0��Ԛl��@`+-�E���E���/���n�z��4|Vf�g�Q��0X��f���1�n��CCEKJ}�O�����Pu��8R�ZJ��N�۱�T;QZ{�՘叵�y�/��t�[���J��N����$��rn���S��>�PӦA�i������-�C�/�k��*�\%$X���*��Hv���EbB
�Z�UE/w�_��2��#έ�ў�^��O��S�)�7�y�D��_[%�J���|�-`��� ��*@Ia�(���bǻ� �}�T>�gɕ\�j!T���/���/K"��r.?��GB[c��w�^���n_�^�?��w����׋h�v=�JX8d�SH|����o��?�dh�^Ա�;o��"���M��?�83�K:�%�F|tb@&&d�C�'�QTAA�i �K��>I"B���fpcXb���#pE��^+��A���o3�O&e�m3�����Ϥg��)`�4���?%ZG}�.o��n�l&�`긊�v% �3,Q����B�VL���,y7�"�sG�ȍ�+�s/6�L�M�*�DK�(�n (����-�9����C
<zB<倫�8@(��aE��~a�<;�;#!Q�KÁ������b���qs#M�߀�2�l�liK]�DiY�/��I���_�L+F��{��yL^�D!@]�o�ACN������hw�j��U�	��l��Xū������i��F���M�%_�lu�"��\�>o\��~�fi�3r^u�C�Uݩ7��P�����Q)����cf�>v�O�)ᮮ҉RC���<�I����MF�E�������C�=6D=����d`)"x�:��L�ȉ*�1i�+��m��\�B�.gp�_����ǅP!��������އ���3kjMZ�Oܸ�Y1��/�W�/�ԝ���q2���:3�y1k��	`���8��а�RgH�=��p1�-�y�vݐ��� �Ym��(�p��|g\5�V�ѺT5����hN���5�Cr�C���ϛ��,�!0j�`@N�-�N�Czy;spw|�C�z��orw�A�eC:Z�*�����+�"��,���Y	V�8v��γ���tc��(��x��t2��7;���LW��!4"���>ًx������n�q��M�al��'��y�Z�5EH���"j�=*`�� ����},ݺ�f�S�=���IL��)�<��c�niU+~ �Ҕ�ODO:�o(C9�>h+v?�W��z��6"��!��x���\
�0Ϲ� ���n��R��n)��O�B75g�;�?3\�N�z�F�PBk�߇N�ַ,uw���bt��Bk���z�çkRCx�O*
X(�⑱D����>a_�4]G8'�<\x����:-�'�� $�z1�\����	A$��1j�DK>g�����!�f1q�/�m�}��=�7b��ݍ���󘛵"&+`x�K_k*�e�%!�i�&T�;�'���D�P؎�:"���5rI��_�TW5<Y�lT� ��o�@}�2���c*���[��֌��Xڇ�I"d��q|��g0莗�W��g(:�^D}�V��6bTR��`q�Ǹ�F�:r��*s���u�F#g*{���jش����ҳ��:�n�?GM���Q���'���|os&3��e��D����Bݖ�i�e 9.� [�ae ���J�)y���l,��{�z��X|��k�f����-8H=BSJ猡&,�7Š�ۻ��|ڲ�����������L��Yw��Iv��\Ċ"����{���ڊa9�˶Nq�Lj��^2 x0�&I����'���0��y_A��q�N��^ӥl�ʸ-��ǊK�:А���̢���V�a��j��,&~�0`����ʤ�{����@�O�h1���o�u��r�"��ufҸy8X��d��C����V����;���T�^�Ң�m�[8�}[�zk�*�A�y,q^F_ 1�$(1� 
b׃4�/l������{�|YuV<�+hd�A�~��D���?B�;�MNҜQ��[�stAp�uRصVy*��y��6u��>����Y�����Y���{�s'S�P���f3;�9Eh}�ڝ?��b�t5��c���JV��t(!ɘ��}�X�C,ݭ��q��_V��O�-�fW�b�-KN�Y׏#S��w��ק�Q�?������D#�6���؈^���zަȨG�\�u�[�$��'(F��)I�!����1RE�o83�7Y�M��F2r��D̞C���:��E<���z������J�|u�1��#%�c�?�-�sY����U�~���7�?܋��\揘����1��_�BA��t9�?�b8/��N�>��ʢq�mމ��Bw�\�<9�]H��.B}
_�f�ߦ]�s6����C��n��.�6 GV�a!3��O���y����z�Fr �J�Ce���\ʒ��R�I�A������8p/��kP�9�.߽v����I�gѧ�'�O�^�gG�kw��I!�j�:"������%3hIB[�&H�ۨ�$��mO�l�'�!IΙ�xj�U�3��������Q�t�C2�=U1'D�h�s]T��̇�vxe.0�%[��,�7�s�)�)%�4�Hj�?���R����������cc��璚M�c�Y�_<ӏ�o�/?|���7�� _���yI�7�X��v��	�_d:���=G\��c�US��4�r�4���$Y�7�:�qՋ���E7�D�M�ĥu�D @��&��V)t����t��	m ��4�,fZI�[ԧ@�J�U>���3����xi �+���n�������u�MӜ��\�o}�t
�(}L��EH�m��i���a�<��N��&��"��m��yrs,+����ө��I����"5b���x;�I�)�s�r�ۇx���i~)��#�=��p?E��ye���s�܇���=͵�/{�װ��O��%2T~�������hY`nV��!y�ДwYyث�X�v���@��Q��B}n�ٍ�&���'OЌ����\kH�j �b�����(�\r�3HlΫ_C^���>�4^�!ilm�U 0���0��e��5x�m!��9�fYZ�kC���O&WhA��b~��e�^ߧ��<��}5	�+J��fԪ�bI<��f'�v{ł��Q�X&�m�|�2���RZz(���v�˸��gÉ���F���^��i#��mNY�cP�[=z�:TAW.w1�t�bAu��??-�g��~�2g�Ƶ!Qb vf^곕�X����%~t]�p��R[�Z_�>w
(%*uT�G��؛�p���/eE�.��eEJ	�5����&�F�������V�Q��!���G�a!���3�!�����v�B\Q9�y�c�rO��s�d�τ��%�%�����2��PWspj��[*��!��U�|�!P�~x~��^���Jٚ�=QJj8��6�fɰ���4���6i��'�uƫ�?K��r��QЎf�n���b��i��&�W~��U�%0o�����鰛؂!�z�C���k���ɔ:j8�w;�K� [9lF�|��/�y�k \�=ZN��ȼG9��&�"=xo+MdI \�Z���#έ��Ȧ����d�ҳ o����Fn���_#�	>Z�V@r�u��\�7�F�y�9nC��b<1ۧD�;�g5P{rF���>/�D	���Ou�&����H�ŔF?��?v�h�ՙF&��˾Mr�@D�ŉH��\�ϯ��-��4J��_�y:�H[����)�-v���v�h�|��&���� d���Ts.	T��B�* �Z��8�Vߓp׀Zޢũ�yG��bڄ����<y|��a���Gl!ƺ��3͍CrӍ��/r�l8՟��@A��l*p�?u2O����mt�r���������%�P�AKm�M�ߤt-'	�s��R_�u����?�+ai�;��<��{�+fM��H�ߝ)a�Q�-r=%�H*��-���9���} �c��R�cp:�����g���xbUy�jG`T�S!M��ɧ���h{t�֤UV�C&@J/��O���i�$�fh���+A��:��&ȻաJ�/e}.*fw-�Y�h�'dDr��/���b"e䡮��ԧ�Is_Jg�r{ B���cj]����Vh��I����F���p5
�����͓�6��
��&p��_R�I]��4�ĽG`��\�G�6������k��s�FW�_26�%�r�����B���v-a���a:�"�Me2I��X������zvL��\��������@�����4'v��H��$�~�����%
�2�?�;��Ok�A�;�4f����[K��I7~��`�����&�I݃�-��9/#�n�:˨�S�Ź[IN�$�`'�k���f�⃽�;�"l����J��F�J_H�0����ٹ��^ʃ�iie�\]!�$Ȓ@9A�<"Ii���V����M�6���5�,���l۟\�k���?&u�ق�Wyu<q����EՖ/;��;A�7|g�1�Ao�$�R�{�4�!}]K.���f>��gT��Ԡ�� C���>�[Y�=��i����ߋ��DV��)0�u>�U��^~jr�����d\���c���vl��F�]����X5�$�����e�c�����߅���4�Y�ad�c��3I��K�˜l�:���1�
~�Ǧh��N��e)W��ʱ|�M^�(5yh�մh����X�����@�N�N�ΌUE���J��v��r�:{`H�5=0�5�S���ֆ4�:@*��ǃ�~�����O(Y��Y��ݰ�z?N{�m�t�(��xr���&���ŝ��$P�; ������r���٫e+�r�<�_ܾ D&�}&�N��#T�:�»5�,���H����S���j�����#������yg.��eb��.���׎!�!�2
ߋ�d�U�Y!�j��*�-���y\���c��2�iZ�؈k<�K��*�%<�۸��Q/{l�����T�h���j+�.4'>�u�JV�_�4)�ipgͬ��� ��2���4I������~H����5�}������H|��)��S�U�-Q'-�T �2��ܘx��G�?�Y곛�^���:��0}�^�N�!���lB~��	��h�Z#�"\�"�s���/��0z��Qu�m/�RT��O�����n��`gƪ���|/�!�n���q��c�jB�8$W���Bj�,!e�8��ؐ#`�*��e��C���_{��(P��:�|����ϝߵ �� @�(���|�wr�r�{쒬d=Dj��1:JR�$���Ф^}�����8����aOі����Rji�u�YT����
����0�Ɯ��ɛnfn��K�Jb�4��=�r�I�hA��3z��������� @'A\�G�g#�zt-=
�ښ��Д_���a��c0[R]�6�|�K��J�';���)�]�-Y�q������]z_m�wџ�<�.���p�߄2���6�~���0`^�OJ������V�=^e5%��$��	�)�h���ݍ�"��ق�@�*��"I?Q&�<��O�l����|ik�Can�& �4��XU,�U���H�~����5�=���@6���<*tt�K�\
;p�g{z��P#Dbh�#K;-?�d7�`S����y.wd\$-ZIDIC�^ U�E
S�ɇ�V�$+�?g���lAOӚ"+�Wx�n"f0m�5w�J��G��􋍢�&���{�%Ž���b�����n��T��!S��±�X���J~k�z"(O�u�-_�j�9�!��c��ٕ=Su����P��M�H�ev�? �> �NO��R�cB������-�=����sk+�x��(g;���;�i,�EH�o����Ly����3�LA�oṠ�\�K��u F��� 9}��C(��w� �·�ʷ���o���?*���'�a����ݮj��2� �:�9y�تGqNn���9�Q�w����㌙%��)z,�����5��1���&#� ����A:ÕWJh��Vu5��������a�F���+.�����v}�3%�hE�LZ���`����U��Q�����a��ؾ��xf�(-�`f|dڡ�!7�m���Fm�d��v%���="�>��?F+'�4Y�=��ۘto��5���A�<��r^�����&����Sg�`wVA%߃ݘ�y�w���O�/W�Y�	&�q��"1b�/����C��Ҙ��C�A���(P�7�d��9���c���V�����*�b�q%�n6�J#F���)wsً��U�%��*LQpT����E���y�JЩ"�ZY��=��i~lCHB��i�oxx1e&�󓐉��k�`�Bn��Ҽ�p�+��IC��JN�Dé��z,2l���������:�/���&ΨR���|a�WOGWyv���Oذ]\��"��j=0x�Ax�RC`yB�e>s��ᆷ�xm��)�e@�E=8W%~�N�kl�l׭{�cO(�1k��TW5����pJг�%�;@5�	G,2��*�K��sO�ڕ���M$�m���W�'�_�+�#��?<��p�~����a[If���L���dy�%/oI�ۤt�H�%8��ƅ��UA{l�n���o�-e��
��5`&:��a���ΰjxo|�	1���6Y2KmG}�[�^;��w��O'�If�A�	
 (�F����U���K��,�_;����4��A���d���υB��26�n���/w�\��uc�Yu>جWճ�h�1:��w}c�[[`���˙񝪬Q��x���m۔�U��im�	m���f`:NB�oU��d�i,[�1����\6W��F�������!
�+��gǌ���k&䔬5t�~�v��w'5:��({v���D4�_�C\�l=Տ<r�E�3�z{-S���7�W�/�p� SsyPx䔣��N�]�[��vhd�Bx� �A_����dX�D�������_� ��&��P�S��?�%r��Lށ3qʞFrr���E���.�:������I������Gm�Q,��)����沈��\��<�x�}ǋ&@h��0��/�y�M��g�;�{��#�d��eF����i��6wx�-�=5|خ�M
?���G.��rLO���������Ng|Z������\��/�0���i��gЕ�Y�Z�<u��=u|c�>k]Peܧ��8�K��F�v�a�0�V��Ӣ�ŢK�&��7$wD�wI;���`4d;�A���2)|�Q�D@���1Te�������_��3��*�s�4VS�"�bF|��������lV�������IF��D"6�i�5j�4=@��=#M��涿���k�-�Ãʝ �d0�������j�׷yn`��k���a��[����� �y�nj��R�*i�܃�L(�-�^E��5,��?�J6X�۵�KT�ߘo�V��u�	R�E,��s�3�Vܖ�D��yM��)ߤ��OV��q���x��E��c�������i�Q���blE-^jD����M{|�����[�=�v�#�����tc���!�2��n�����8��}?�ed��~;�湭ɮ �����S8�U`У�w�v�:��HY�4x�6��꣮8�A�ՙQO���O���������q���y��r��m���9y�e$%cҳMEі�G��,�\����3�WZ����"j��0�$b���0y�Z�W⎇��7ع�p��-߿�f�u+R0 ��49&Qg!x�������()g�߸>��:h�W�/o�@��|�i����v&��K���R�d�\̄\����d�	v1SC�(�=��%@�+���bM%ӋK�NqS;��<:�l-�3�FJ(��n����Oo�7�dw����f)**�'{��ab
T07�7ɵ'�������Nr�(�q�~|X�k��Vm�AxW ��_j��p�;7(>W�fg�I�R�3?5�A�p@������4�N;���̋�#c�썰��@
�ઋ1�ꂉ��Yɸ����A$<$䥬K�;���}��`��_(8���Ӳ/��+���r4�	b��p����
i-��^��*����'�;]�֝%��d|� �p5z{r���P'���IZu���''�mIv�rT����e ���2�˿cW�iVOr	a��.PЁ�|�#p�4��J"��#7'FʏK���C�^_#��jP/E�4�@�50�3�H���j퓾g�J��'˲^JF�*V1Awǿ_YS{H�` (_gdX� ���զ@�KZT�Q�;�Y�vA6���r��оB��w��Q6,�?e3�6���U���m?��9r�O�{Z�qc��P�����N}��x�g��sQ·�e���jśI���X�#w�¼�h�$���G,�ί0�'�X�������Ѩ7��@:"]��P|�r��;���{���/z�Х\�J�2��bTЋ�N��	��
B��Vlw�'����w�ɞ�H���E������%���_ach�������p���/˺$�;�K���۾�v�ƥ�">��Z�%�l�9�$��v@@�����l Ļo��������hM�;�.۩�_
!�V�p��^��8;�����5�}��282���0nC�0��6U�Uf� 0z��2��1gt�#"�.E��0�]��W0���Žˍ���$� eer����O�-���P��0��YG�����K[�FsJ˝�yXT���`T���(�"2I��ufks�Q���e�P*?�����!��Z�6��5�)`���ӑ:B�C¥��� ���m��~5l�urG��ɯ�481'�^]����=_6����"�9���b.��
'>�2C}]ON���0�n2�N;��~���'h&}�'b�m���v� ܗы�Ų�n�f��(D��]�qL:R��DS��Z�sd$����Ѭ��ğ���W�X�(��g�Yd�%�D����ڟg�;>��!�;��F2�؋��ߖ>X,V]3v�˲g��>
:%����%���Ex�V�F>rm����`���/������>G[�,��jmf<��x�֛a$���҃2Д�+�Z��ɲ�"�5�~׳�Hp������\�Ē|..p�T2
��1��"�1����:I�^'tW��N�9�rIN��_��V;Ǘئ_T������&�/�G��(9/����>Φ!�a��.�Q��eu��rGL
���}���\F蚶~��KK��ӎ88(ND	�����J����5X�,&ɂ�|?X5�Y�H;E��{�(�ӂ,����H��B���cҗ�o,>�Jk�<ru����{������K�E����k�r㧀�uy<��/�<&q�p�s'W���RPWJ��Y遮-X�֣�i��d̏08J6����4
��(�����Լ?��������l�6{x0:�/�r,Xy:��S|D25��|
cA�#O��(Αc��U�/M��Ǥ�;kTw�2R}<�\�I�"'��9�*	l�$�ØC'N�,�p� �fw�M���4�8��@	y�&��1�Kz�T�A��A�}�!������E������[�5QM�uEa`�K����$*�����I����jbX�dI�L�xZ�66�/��N3ϭ�+H|K�� 04V"��s�d������v��h��5���w�V���\f����,�wJ��;9����^��Fcq7��������z��YK���^�i��)��C��%��+}�vIxDM���d��Y�#8�d~>߈z��-c׾�+�dDf	�N��P�,^�����f��h��4�1�Q	����n��f5��O(琨+�z9������i*��'Hg�=�u|�BA�a�5[K2�P�	���}3���t�V��J�I6A�1R�R��1��cY�Nk�鎲�@G=��՜/H��"Rh���-� ��1*�!'0�g�Rq9H��Qk��E��P���#5�S��5�:��d���+�RR�:���65��m�Ձ�e����Ʌ� =D�1��}ȥ������y��[� v���&�܍D$S�E�e���I��d���>]��tفF���^�+D�+O��R��`�3�j�d��Ue]5f��
������-v߶l�B8Y�s��RJ{UMD�Wd��GQ,t�2��_H�wX��O#��D�OI��� y���J�xZ��W6U	��c챭�5�xw�F�v�"��z�ꋪ�P�{o��"3SA[+NF��*ݙ����6�y����ގ�/�>1n'fU��Ը�Z��3ڙ��9�X��F�@fs<i-# �R�����˛!��?�͌�hzz$Y�CDEirV5��
豋(�[vc��{������@�'H�h�-�IFd�A�JΠ��R/�CG(��-~ʮ(�,Ä��N�G����-I�dW�ef����Q@�s��@`��o�V۟�!�g��F?����h�����F���f����%$,]�;û'z3�6%�|�C ������2��v��2~/��ܤv/4��]ƴmma�4YA��@�}q��'pXs����6��� ?\��<V�G�@ɹ���c�W����c�j�� ��2�� 2>��s��or�sVv�*dU�|�x}M�LƂ�m��h��I�n��f%��.��)�M�!g�S���:��T����'|eyc�Xq����KՇ�Z��iI��Ҿy+�D0�c�i�G��Q�4�*�mTa��Qcea8YNph������燇���C��j)_��Rt�_�<�RFTW�|�}�&��%�]&� z֮�2�d��GLn�u�,��/��:��V����5���X;�7o�L�hb�z)����I�t*E��_ZR�z��a'yaE��� ��|����ق�
��^0����l�j#������~˄��fl}��n�����#��o���\���^;���>�W��m���IXq8аɏ�cXN�3#�I��[:��� ��xFL��0�}/�>4!w]� NNک�T�.��ds��.&X��l���KS�R������M�5?����KI̬"��B�>EO5laW����廍�[����<��׻;��F'���Q%�{��f
�P��&�P��73�(�(�%@�Nw\���C�"�#����s����"O֩�cOl��0^��k��xE��x���a��\��8������H� ���AQ$���Ip�k��s"��|�GV��g�ƕ��N�a=FK�KũI�Z�;��#fZ�C�bW��X?�x/Bv.�;n��,\I�أs��g�.��.}0��v.����̬�&����'-E������U���Y�����%��(w@?�����v5�?����0L2d�=�H���d:8S��
���\�YL�����ࠕ�����`+���L{��y!&�LU�(D^�?��r������yf�&���:����iI<��A�UdG���M���bT=K=�u���y�u�uq������}i܉��qjH��6[*`���9l���}����i �^�U	!3���F�<��/!*�p��b*��_߀�R�ӱ�遌bđ�R���C�}�q��/�^ݕ��ځ	�&$k�u���#�G�6�����)��}~���]iů��K���vk��JA_+�R�)YS��o����s	5�Qc%�+T��{s2k�a��{��
H�(�ܸ����>�y�����]B���	,۬0�{
#�<n��h(�f�JyrVq�zk1����<I���>���ɽo�#�m@�&�$�Ws�(�iL�aew�<[]�K�i�PQL,-���k��eE;jX'�S�TǇ�!�t�U��)K @[b��/n�;<~����u��x�l�!x�#���)S�+�������V��6�z�����XQ��<��e��G3�c2H�L^�<$�3",Q��ϭ��W��Z҆�_��˷]\�;����L�g}�����r�~�	)��`��m�H��U�%�R����5-�
tfȏIU��ʟ@R�ǆ1\\Ӿ�Q1Iչ���3P-u�Y��D�|���K�N򄻷�,�f���i��s�|�aӿu�xpd���"��YΗ����v�a(Vp�f��u�7F��b�'��ƙ�uP�i�˿�o��/Z�����q�gF�'N���ff��Q'`��yY�ܔF��o��C�9�������3�S�CC����s�%_��;~(�K�d�����.�v�p����!
j��^7�dպ��YU�ӴgGR��W@p���.�a>0�l��E�p��uţ��q�ݻ�dVF�G���o��y��~.�����V;�૨F]�І��<��I��o�X���>]��3�ʄ��F��|d+,���W�Њ���f��Y*fn!v {��C����|�*�~F�,g�<��OQ[��f�
��*_�߹��m�J�N�J��Ʒ�)�Ҋ�����n[���09[�����fZ��M��u�oW=/{�>�)d��ߙ��ΨcN��QdJ��?~(�a�jFu�ZCaAx�_f���N�и���+V8G�����[��7��g���G˫`����\�6a�0J=G.��Z��`�b���^�xa�>_D)�[:Ն�����=�C�cqq��Ѱ_
j���֑�9���=����i���(0�] �x䥒�)[_�f�Rӽ�|�D��W�1��U�rS%g����H`z'� �7:N�!��ٵ���^�"�8h�h20����/�&�7�^W�3�a����%���=_��Cڿ_7��H�L{0�����{}�3Vs1��]�]��*z���$�ђje��ah*��U���'+w_�M��v�tbPKXǰ��S˷��YN���3���22|�G��]9�F5��1����;&��l=�
� ���`���`݁��F�aT��C.�6����g��C�EC!�,d�6P(g�	��#���d;Y��܋�m����{�J�%y�t�Os�]�s��֓Kq�R�-8���R�y��v��#[�B2��8�\���� ����[s)���P�aw�p����Z	)��DJ�˵|�5��D��	������z\Hr�u] ��Ϯp�#-��YLwB`"r�5<���"z�'?�U%b<���1iK!��p��ڑQ5��$�~�:܏N��rA n %�S�Tū��fV�wE�-]�#!v������}y2���+�0�{�uAؼ7t���s���J�)�>���lh�Rz�1t��O׋;>,�מ�Q�-df��5�yS824@��s�Ht.¡�ȼQ�O�`�Ǉ��>��R_W^�6:��{�	��H�6�,��5��=xCW\����N[���O�H�/8����J{����/�U�KӇq&]Q-Zl|e5Σ*W@��b�] �0^u�������"ak]��Y�"���S�h��d��s%[��-e���g�KCC�>vIN�L_�c��������(5��E�{4kp�� �@<�G��l$���6U�b�D��L^��Z=�Rz,gY����}I��Z^�o���Y����m��!P�H����I-Ö�c���Mw#�Q4/������v}?�Tȏ�;��C_�3 ���ɴp4��{�/��'w#�ξь ��.[|-l��2�/�	a��)1�я�/9���J�i��y<I#M����u���wS�PN�>�2�˗ ���u��4�����p%�:ЩcSxYɟ}&!% n�Q�v���Vĸ�k��T/�2̄*�(uo_Ē���c�D���.;ٔ>�� ſ;ڥ�G��}�qʣIM�Z[�}�>⌫�݊�b�{�Hr��,[p���GY~E,2c]�S��|S6:�@��=P��χę,�gi�xM��f�G������3�\%%P�7���݀ipB؉`��#+��Bl�V�3��čg���������bx����1?�èγ�eE��ah�
�+��?_jq`�}��%�t�I�"94̚��B��E��r��a�^��b�&���%ύ����3	���_A��胙n�2���Z����^�ڹ=w��H!�"U����>\7�wF�a����I_z?$ri���u��]���
�%���`\�b���"6�za��&�ބ(c2���F���%������Ʈ	G�_�����?�d)z:���;�#�ň��G�]�L�a7s0��:Lvb#�a����sI�����"&�vD����ǯ�>���U@*���?�G����է��65�>�5ֽf��u;�$���P�e����~>.�X�J���t^o<��o�i^8Ȑ!w�c�)QgC|�Sa�>�U�G�SF�f��`l\�U�DoH ޲f�CP��Հ-�8K�����q��+�'+l�����3��(x��S	jmН�P�Rt�}mK7h���H�u���pe$HMdYJ�����Q �P0vQ�7�x3iS���/!����%hw�:h��¿�B�r|�ˆ�ڭ�ŭ�e�}
=^⴮Q:�l�ۜSR���h�¹�r�Zzƒ�+~i� �VCe2.-a�s��Y__�)���o�S[t:�hW|,vc�ۓ�yŨM��z\�s�+��Z�O(���<� ��4./J�_���=��4�us}X8M����Nq�͊��6��wr�� j(�.z�o�X���_=�P~��a��z�k������K�B	=FM�o�Ћ�1����@,n"�#19�@3�����t���a?���̤���7��@U�QF7�ѽ6wsWXm6����|�ģGA���Đ�?>?E���,N)�_�v�ds���W��2M �(Ձ
Ƹ1�<��A��3�S��(͞RY��8)<K+��<�\�z�gT%�č�<�`+����O�zf�l�}��Ug���8O}eĊ��l�X�>� ^b���>B���cA������T7N�}j�����&�h又R��o���{�C���C�w�}��6�?�#Q�5Կ��4���a��e��_���ݤ%������'<��#��o�l���E����Fm� �����1~h�������M:s7�qc�]s[�B��p�<��*-�t��ON´�� ��,��T�F�ve��}��0B������1N�8�;z�/��isj�5��{�Y�m/)����pL
U�Ke�Pc�)URF�~&/��cZ��-01I]VdC�B(2^�?@��ݮ>�ƲԻ��I��r��*E��$xL娶&��� s�^�Q�S�y���w���ݳ�鈸�d�^^�IM^)g���\�y�	[d˅�8��5�Fn8����]�*щ��1���v:��w+�Q��='�w��Hn8� �.*WH V���	q��a��Ue���j��8�VG�`Ji³i7୾_&��x�V�9q}������Uha�˝��]�)���z�ɰ.t��,��d�eI�hn��ǰ�*�inD2�5��'��_Z>��M;,%��`@�su�n�mě"﹔ώ���-IO���8�E�0����@gђ��s�gH�d�
1���~�:$�gW[�/Y��gT=�6��_�W�� ?HZ��ڲ7����_��Ig�Ͻ=��j�%��>�?�_�C����k/�n'�w�P�KmR0,�ҳE��;�p�9mٖ�u8�)膗SZ��V~��H埥@@5��������Gx�A|�n��ksm�qT�Wrg[��j�s��n�9��J`W�q)v@d�2_g�Bt�dp�/�)r�GO��ޠ�-�/]Zܗ�j�<i�f���}}G!J ����M�[��u:��qhuT͉����>�o�M��*�=�H��R3N��)�a�C�JVne�سE�@U�C�q�U���RD�2*cgu�cD�g����w6���>9	g�FxC��Pi�Qd���u��;UNf	�-fݻ��l����%(j�VN�1�:v8��	����tw[�4��M�Ǽɥ�֐I�Ϭ���]4vf��a�jGGy���v�(��B�Q6�RY<t�"Q�X��3+N:J��y�\+��އ�22XkBד3v�74<^���/�X$	�.(R���0[jŷ����t-	�}���g��Xu��B@p
���Pr�����89��#i��C�H<\��4�T�v���R�j��!&}���X�W`sb�_�{[�R���|"����7���B����w��1���ݐ�(]����s���w���I;9䩥>�'��-������TB��|�n"ڴ�@�f���ӂ�
#� ˼�6wt�Z�O6/N�T~�ݵE�.��kҴ��!�VO�]�7���a�]��%��\ˇn����5���|�z�ЎaZ�D�[�� �[x?�U���7q#Q���{�"�s�3YE����y�Pڐ����'�T�P+���������Ô�Մ�?������)���6�_e�ݛ/[�'f!�Ǩ�7��a�1������	����HD�C��+�K�����4݊.2�0U�?>��1f~N?
3�FPFe���0���#��ez�y�R�jSf	��h�*B{�8��Nj�@�I�"�y��u�F�c�ꅽ�X+���>�e��(�r�������~���N�dk	�Sm�P;�r����"�!�c��2fI|��Q#紈(R󂖭�k�\��o��Or���h��7����.{���]wš�V��n�bC2�Л�O>Y�??��d�*?�`7�?;q���_�6����K[���/"�_cdV�a�a�>��~����=[��6�gWPi=�$&�hgnM��q��F��d~���g~�JLgEz 6Kۀ˙�� �|�Dl�\�J�����(ݔx;� Iq��%�7�7��$����(IՃmJ�3�����)�'�5Ʊ��IA��� F�����ɝ�y�'L��vA����*�Ʃ}X],��p�w�Q�j醕�m�i�
�q��F<�I,Mʝp<���E���dWӺN2*�yTf��_!j�5[`n���C��>3���MX���v�nxr��S��\�|�����I@��G ���Jδ�#�ev��=���A뱿HU�M\j��E�gy�Bc�2*n�*��5d�q��<!W�C��l��mu(7-����jR8�8F��$WӷX�q��O:�P�:\��KE�~�� NބE���ܑ�͓�Y �h����t�.k7'��\Ҙo(�8��<��Z�-θ���%��+{��Z�&���[-�7���[���Q���^Oګ�����|�����mÂ���1��[70����s�����:�Y�sw�X.��� 55�dQ��&�'�[< "��� !�$�0߲��bՠv���S�t{X�
�U��o�N@�¶������~$Fݿ-�~}BQ��<��=0�����t��@���R����fA�u0�HiNq,:�5)j1����_�R'r�Ec�޹�� Ļ-Ű
6Mm�U�l)0+�h}���
��܏w��Q�/�Bj��v�[��9�k�Dm�9B?5x6}��U	D˟^*б���X�E���l��S����	�_���S�;�d��w�7�i�Տ������F�ճCɄ!���s�Y�Y��E��h��nʼs��D� Y��&~h5}�
����^6NO����v����s���?�W��nf��V!4��L���.�'��U(����X��H/n`R�	�v�z6��kO� J��O]���e|H�l!'�VzeR`(�n<ӦE~@_�.A%y+��6�_��[���PZ�)1K��f�sI4:�B���Gٟ4�:zF��; ����K�rTDnX�g���*���&�r�V��ql�@��o��E*x�ݦyc��ݟ�(�_�7K=!����x���������d�#��M�"5�Cd�S{��Ґ�|�����-jW ���r7E��(�1�Z�U�cu+���v�vpu��.0�S՘�n���p5ff��G��c k��W��&�GT� ��^��� �iۨW@���[b�~�-�W�x��8:̑l���උp������.('t&�Zc��t��'�r/!���O�7_{GT��	e�:��ޟ��4D"�/#g# �.�������kA_�mS��sF��Ӷ�ZњFF
1\��3ԘZ�6v@1gw�N�`t��[>��?ްr8��|�Xō��uy�f6}�������xFaVw������S��T6���boW"?�ޕ3�\h1ƴ�H��L�`F����`� K�� �!��e������|�@���	`��-����	�4���6g�~�PB� ��j�\j8h$~����� \�̆6�학��n���}�^�5�.�t@��ր�\{̔�P��X�/���]}w�Ij�V�.N����\�Z'jj�w���3ѩl���t����^]���G��Y�3ՙ����2y��V��J�S���+z�vg�C�2Gu�L7.���8GDy�ě��h��St1[=������ԌO���$���`!* d�W3A?I���2z�wLW#'�ҷ_���#{�&:�e�\9'P�l�d��(�<�RĜ��<%g� �)��R�{8���������Y��~w������ȱ�|hڑ���H����e�T�����~��~K��z�S�����ϻ-n���OW��Q�I�{����@��UF��M-)TV���z���N]�f�{�zRu��2�]_��M�- �̆�n�bP7�5�kB�>��͙Q�-�i�%)�d�BHS�6�r{�)�
�9ccC- Q=y�sk��N���aA�9ڷ�0l��� C�t%����zu/�ˬ�y~k�V%�gw�@t��2k�M{��}�1Z��=U0t��ʆ��
�{�;�'6"&��em��	2�p6�Q.�S1�r* ��N@p�_��u��V�w`��ʷsE��Ӑ�K	��ZN���1�o�n7��4��P��>4��-��Z�>��]���Aju�AjB�ֳ�����@ �jL)�.qp�x־h��.3�Q��W�B�j�ե�S��<�n|�ݼ[��<Y��z��8"�w{�g�'Ēo�#c�.䕐KK�w�EB=�82>�Y\� 4?��@š-��i��
�c����[��,v��V����|QL?r�P����\O�@��6���@�p���e�|������w��m������N)�s�[�HM,���_���T����O]�
&�ꌥ�iS�S�x�*��Vr���F�b�Cͽ�g
�L:a 9��x$W��!#���e�Zֈ<)#Ri�8�q_p��+@��ꟻk���ƻX�]r�����ّ��{ښ�e�x��[���{�M�"�y�[�+��*)�)	IC�djf��{?@Yއ2�_�^L
؜d�&h�^:hi�g�y �������	�R+Do����~,�����*�o��T,y�[b_�;[$�"���<�ɑ�砿ŭ�~���b���N���HQ��%�&�6-®g�=�k�*_�̓� &��7珒H'N���njy�`�HOu���q%l���� �W��эdV�d���N����ɭ��k%��ݒ�Rϕ��^uZ��m]ׄ>J番~䁹3,h��;c�����P���1N��<f-0J}#V��k���?8_�?Y��.���&` '�719ǝ� D<�ɭ�;q�1�ژ�y;W$�2� 5`
Z����S�fl+��S�D����]�F��;��^Vw>I�p1�S�i�Bvue;!̫��4���/}we�����..�h�r���> �X����������t<t������ Ÿ�p��&&�2��2,'���m�B?!��3�T�����à*Y��<-$1m���K�`ܞT�fY��~2�7xx�O�����0�谛�
/��&t��-�74Mi¶���3�})�:���� )�ӈ��Eb�tv�iǻ=��X���H�$�f�[Z{�y�~/]��%��&�>#Rl9l��K�k*�Yt5/^���!S%Q�9����0��b�qt`2���?˖-�^0Ae=�N�������.|�k+�r���H�X�	\���{ّ�N�����р�o��X��_k#(��^	��[�/�s�&��	׸鰞
l;.J{QJ3	���ST�İ4H���+�P�A_9�5����ud*��=r�h��z��	+�`�RX,�6��Н�vߧ�E���4E���?�ʙ�ᤳ*a�ZKr�v=\$r�e_�:�h��aFj���ؕ2��A�u�q�?g��g�%��T_:Ѕ�AbR �߇�>�x�h��a��~��zm4��e@��#�q]���F�buT�d���h	����P<f��!��ײa����<(�x�5�������W�ROpݧ�'�8�;�.j3.���+�=u�3��_@w�-�LK{p&Ɠs4��vK�T��K4ʭ�uE���@��:t�������a;CS����HMk(��O%���ʾr�9�(,N���MubK�Wi`B`簝AmPƌn|��0][^��@��p-�*�l��W��`�Z��m�f��"
�aPo^��Tƙkx?$N�C���L����RT���7�5'��b��2��J�f��XU\��/���qF8�Oތ�=`~���9�0r@>�l9�"݀�8����\�a	�I$�g@��Y�e�/�˝X�#�MƢ��2��T�#@y|�?*������X�lN���}�����d��2	�0̓b�DfP�d��i�#�,�H��/����<)^�!I&�J{��ߴ�g�m�X�zI,���?Z�����ݛ��X������~��hcw�]<e"j�DD�bb�a\:�C���G:]G���\�*�9qm��9���l�F�<��)n�D�wy����ҏ�=Sw�zM�QX�>��3@c�+&�8�Zj7:�C���5_-f���z���/�
�5�S�t�O���ڃ��@��^����OT����*�q(hH�2��R�_�f����[�A���![$;K�����+�1&Njdz���.�F��&"|)B�J���B��t'�7�w(i���ƠN3AFt��[�eMb�VQ�<q$�M	��1���!"9]�!l�Lq�D���P0���a��b�/�S���1�6e?@��Rn/���ݰ����	�Ko�����c)`: �}����
�9H�l-����T��=cAY��8s7���;j��7�B��K��O��M�a( ��6�S��9	�uR�|*�P��R�Ypy������6�<�hQ{jU���g��� )���.n���]�d����j��c\����^�W���P�gm2�^���#�Z}�J5<�������7\���1�t)l����*l�0�s��������l��3�2ۘA�N�P*�`� w�j#x�v���.���15�_��K��m����ys��ǩ�3X��=j��d ��O�a}�\RNF����31�EF���[
Y��Du�`W��A~ĪI�Ԉh�S��Т�7D�F��Q�W٥D�U���}��,�ޤLw��JP،$L�4'���X0�b�
l?}�U��9����u�ï͐�fI��ư�bЈ��,$9#�Ɵ�L+��u_��0���p�����p�]+ȭ��۝�Bw��g����\�!�y M�V�2��aKR+1���� ԬM�Kî��e���[�^�
��mw��(	�ϩH9�������:�џ��Dv?y���P�\�o'�fSb�&��K*��s�bC�Ţ�Ҷ�x�8�Zf��_K,����C�aSZǇ��W�U�{h>߆�1 h��F�i��;U�1����Fv\���K��r1�z#l��_X�����F&$+œ��-'�g������2�У<]��>�È��qw��ރ�B^��ZR5�3����1���Å�|��b��0B��"����M��,�Е�ؗF�!)�T,��e:�h2|��4V'��_�n�8�-��?"�0�tI��l�҄���aB��\;!��[􌞑��è�Fy�.7� }N�Q&���[�le7N 	������	���*[���ue�t��H@` 
3��y=th v�dA?~��/׭
p��	���̬v��i���Ùc0�w���PP�� ���I���Zt���{��&X�P>N�")cFGX}���A��\%S^Hˈkܭ��E���Ga5B��p�-�+�[9�!��#�^7��k���͠��뱩e.c")zTf���L���,s�����y����/A��4���HM|�B�A;,h�L��ɀ�B���*14x�F�`��צ{ue��4�SX�+Q]�� ��>+��6u"V�w�r��:��x}{�>8׉3��EJ�YH��YD;��>����4�_�ٌ�D&H��s<�Y'�i�lV��'
{m�G(ѣ�RSO>j�Gųś��5� ���W>�J�p�®��FYC���%��PK<_]{|)�$0�B�-�-j�X�Y���	�!1*8[�Q�k��c;l0*��~������?�o������jv��}�YG�Bz�чN:�(~�R�m�Z:�a�IŴ����&��S���_D�U�$H�s�V�3�����N���@�;�/����)"�G�>_m��
�.���J�cI=���=�g83� 61�=��Ou����f'%?vm�`fd'kb#�+ָT���_{F�T% �%H�(#��9�' �n ��ى���Ɍ�f�%�^
�E��(6��V�[@��2X��s6d�G��N.��h��6�lm�a�"���1
�a��zy����o��m���\�J��,e]eΔn_|\�������ȸ_�.nX΂@��:���Ԥ?qSpA��恿��J�m4
<Oa�; 	���]��!�tl�
[f���?���$o� �VrL�f���҃xe��:�|onw�Ą����L3��W:���Xn����J�s..���7�$wX�U?�K�F���HV�tq�z�3���̅�I�����w����>�WX9A�)L��f��=�U���
�����s�)z%�����~���:f��D�����[ƊE{��}\#S��V����S�U����wZ~Y�wW��y�J�53�P����QR��0���y��x���:-s�M���Z쇦}D��!�
A,�0�M��>��̗a�z�~)&m��q��%��e��\�u�6��󖩏3h��6oI�P�x����%�S��,Vk��7�����*�O��Qu�Z�������C�(�~+��#����פ���k�5���Eo.�w^/����7�.+J��v ��1Zݽ#Fa�MS.Tg�N<�<D������q�\�����Ů��]��0ҽ	��W��W��v\$�8�P�CiǄƱ4�xeW�O��y�vd����֓��p��+[J�f���n`4ʱ8pʊ��w�l����K��S���9�(�Wа�RG�g�d��a�u�ߡ�}��(o��F^���x��Ch[���>�4�Np�_��M��jMB&�~�.��n�X�c9��%�۲�%%��+�%\���8죟K\@/��y& <�_��g<���SZ�k�q��6�k�Z�D��F:�4���Ě��+Pw&��%�G��ߓ��nv�wRle���
���Ry�������DwV&�q���kh�xPֳ6����m�B�	Tya��:�k(��������+D�҅�-Z=B��prKY@�ż��핲�OJ�崝&����q�kv	��t}���W�����y���n�2ELHN*�/e�ig٥�'��������͜��{I(�#��c� �t��,��=�*��3��⣦oO�xĴF��3c֋�ٳ��@r{^�.��p��yyP�y��a��k��x�+u��'8[N��j�'N�w��T���[�Ê���a�?��F��{�V�s��+�B�2��"�".��������?ܐ�D�2iІ���q�Q5�Pt=�4ӏ�qZޡ�>�����v���^����`a�(�m�/92�H_/zeV�屓e�&�����VPv+#ҩ���!���q�\�4����W�1��Wc+�����d2���,fXw.��嘈��^�TKL�#���Sχ9i������a�m�v���D�#��`EoM������85
�֣Oc��
Si�&g�T�O:����2E�~����������s
A�b1]�y�3��zQ9i�Vz0:u����O�z?j�	j�<�\������7�.2b5:Gl��=�}G�s0|QQ�����"�L��w�	�>o��h(�d��j�c%��n���qS�M���¼���̖��2��q^��sS���r)�J�,v,�1G��>`�ޟ<B�b 1bv1��Ok�k������T9����t.�?��i��QX4ƃ�;Z A�ɾJ!l[Y���fX�܉��,�8/'��A(��fQ���ET�G[m���yT	[��LF����M%���к�dދ�pr
��G[N�.�)%l�-b`�9������䩺;�Lq�!�6�F�3�HdV<޽�p*��@����WA��&k?������s������%^�j����ׅ<���5n:w�Z�i��6�"�ؿ�X��Ig�W�u����,��̝����^����1zn]��)@Ƙ?�!�=ǋ���9U��.>w)�0��~{�0��2[x� �틍��k���]����S� Kp}��|� ˍy��!��(�BJ�z���-+�rު�������)�ND��ű+�
�.�Z˻s��#���fﴄf�!�C�I���@9�9q�J¤�RCn9�t��c��g���+�[6�1�/�/�%�ν�H'3�fDl;��i��д<�-Tx��([��#Wƀ߻P1�7k�&*G�`�f���
���O�W���y��[�p�')bOv�HV9Y�>�Y*^�Q("&�(��c\�)�Ħ��;�j�p�"!Hl�.�L�I(��*��jR>QX�ܡ�Z��z5�6���Կ�P�N '�LI�y�i�E���=�=�Z��B^�-X<'1qw�AX/ۮ�z0�-��j�
��~I���v�ɡ)8e~���h=�n����ǥ��;���ݝ�#_swQ��X����n����xς�_�z@T��Q�ƿ�]�sh���p��v�깈�?:�\���N��=j��v����UG��
�]hM�9����sB�����c�ZQ=�es�)1�"-���
��V�c0Ґ`�h+�2[��}h�8���6d���?�=EOCf��v��l��$�Ɋ�����y�D��4�b��@PNz�.(csC�ܫx�C�0D����I� �^�i��u�`<�E�8�(���:���L2?�w����&F��U\C�婙�
�VB叫D����t쵒�=7v��I�R�fYh�����-#�ߗ�DQy�>���k��A}~�0��S���?Mؘ���˂�{�/�B�o��7/�c�j��(nAm挵|���f��?B��Z��?gz��������8���f��^�o��4�w 7#�WP��xOQ�V�������('���Q��UYݫ>��3�\weF�E�o^t���b>��*�F�:4	k|$�hcsPeb&Ar2��FvH�R����q���^A#8S*[�������ꎑ?�W.�<����;���Ic��z�����,ңP��
���or{S{��3o�����!���u���6OY�g��0�7~�����b�$��I��+�/ua�������:뮴�Ԟ4�M 7!�
~`W۽���G�=¹(��o@T��.�X�Z�=[�@�U��s61�0O���4OrؽК�7���;D��QpM��ȍ���H�窎������Snz{#��_��6;g�¤&!G�e�� U0'���䚐O�q����a��3-��_3���	ۿ��cY�U�ƾU�_O�4/;{�޲��Z-Q�]|0]�$�]/q3,4�٪ﮪP�����yU�K�\s�U@jp��J����z�?* �-�r|�(�HGJQ��pJ\��M��_^u s�(�A��ێ�!�z���:��+{�3N��E	��i�3��`�s u�����^+n�=0�mZ�������5� GW���a�,𧽐�z�s-%��!�9?hw��j}�8�����W�g��xqt1X����c/�NX�/$���W��c����ǋ���?�����$���Q�R:=��:�5�C�ל�?x�5.����}ʾI��4�].�*D�=���Ե�)�m݁(7�����w�-�N�s4d���<��1� ���0̛�3���㍰��>�	F����
���N��5Q% �hG�����B�9i ���z�u�� |*(e/�d�eG��k��n���'6jt�)(G9_
��Ɉ�6��# E�K�'��<�ã �q��I��FMĔ6.ޖ�4�\����[[ν��j ]� �қ�\g_��lY���C+��rVO�A�C�oF���R?5��B6F���°�|��[���*���`G��Yd����>�#A�%�L�ʓo���a��f���ꌜH����wqFk�8+�\��SV�|Ԧ�Aʠ�p�ὗ�ם�ꙧ���_2��MQ��@��1��Z1���'`��/Phn�=���J�Q�PU���Z/�@�ӹ��g�bvp���j���vyT�g�Ss�������@��-���kf�pi�>��j��K�.yO�
�Q�\�>��A��o�2��;���m�%�ۆ�+~��2TJ,���^-����@�����z�1CM�R�3������-�|F�����Lb�'��9w���KP�+���!�;�<���+ 5q��;��nV�����բ�]��?�c7y���z��1�2d[���$4i�GI�'�j�#��Y�C���7_
���5����A�65L��&	�<wK-ReQYtY���
e�"4�1r��CWk�NJ�M��Y�AV,�)��u��վ�VJFB���� {�Ď��z9�bjaA��?�2���Z%��(|�o[���?���:'��$���#Ȇ��o�!����	�!��4i����x/��?Y}�FQSPn| 4�0���2
��t��IU�7��c��Bz"���<=��S�O���`�z(�����n�=��n�L�đ��J� O��EO����*�<dL���Rt��4Z�}�~̢͌aװEMD4H�|!�v��\t�#8�p��elK��>�Y�]�'ډ����y�P�o ��A����=�l��8�3 ���N˒#�<��Y2�sT(��=�3�Q�]��aG�[�\�Ky��#"<��ByʂI��yĮ���	�?˩�j�c���A'S�����H�pՏ�U��b]	k������_+b�����������=Ҝ23���i�kcuՙGٗ\�Iw�K�������mnn���g�.�/�Z��v������8q��H������#�����N8R�/���zԸ�7���7�!�,F�]M��$f�m}Ԛ�<ɪ�e>~�*��v;�#j�f�#D!Ee�4J�s \Ux���=&|��?8�Z�a��h��1m��kљ/��ۑ&������= 6��Va��b�x̷�N���g�;�_��VS1��Ձz��[ɡؾh���6��C1����M�4��B���j��B�b����s0�X%P��]�W�( �����`����rh�����*�7Kb�(U�G$��}1=$r1x;��]!�G-
��5Q �к.M��!]�ޜ�n�;�ؿ�'f��Xv[���Jb���.m4�`K����ۋc=����A[T��J�(�
�}���MX��%!�^���aq�9��h9�v�$�9��尐�$���O�=��0�E+�\�XE�8CkP�z�ovI�+�*�z�Z��P�T1��\z��z5�<���f���>���#&�j�,l�\� _�OPPE�f�����-�� hv�֕�������6þ�H�z53��dOæ��>�bk`�� �����`~�A���}�K	� ֶ���N+�G��-躱��p/%�:]���H1�a�r��:m�6��k8D�:��A7�sW%:��SyY����n�t��i�@�X|�����@��z]��O���FH����Yb�[�\L�d*} �z%���I ,�t!;g�e�(�G�9��AR�LtAWG��S�;:W�Pz�1Eo�Y�V�_,_a�� �5��j.�l����fbd�A����=	Wk�[������3��̋v��ܮ	��O]D��,���Y5��U꿷���ʩ��K���|`s�&�l��?,w+)*Pn��+�Յ�?��7��}��x 	��D����-��!2��v�g~���V ��`��q�ѯ0��j!���k�u����3�4�09fꀤ(��J�����U&�tUN~��sӁ�ͺ�h{S������;`���ڊ�Н��*Ù�7����fB;e�JM�K���i��h�=�p���������E V��B��T�G��s.ȩ�Y��߹� ��G}�sr3����s�F�W@|<pe�	%N��6�a ,%�MCCO�T��h���8��k��ZƳ�V�����[3ȎM��T[^?t�Ͷ��Ⱦ�-nD�=E��
);��]>5�b2@���1xjL��6˷ɿ���Z��%U"�B�O�e�];yV�����{MB�if�,D�&*_
����
aa�,4(c�I���( I�8���B�"u�%���c��6�ޯ��-�3��g*K����~���5l�
f�MuI���V[֗ح��uF��fٹ�ł�_d���X�"���FPb_N�1���ݧ�d:z-e;�N�;^-�&��T��h� %_�y���[���ul�P�bU�d�B���ƣI�Y�����/��m
J�u�@�r5��^�H�,�I��)\d��z�D�/4B��t�y��뇡�h-[�j֥�+�ڄ��7l�]���y���������LY�(�Ols9h��9�v�_2���x;�X�@_��|�"��+?�]�/��p��3�G����o��x@�H��9�x����9�o840�'��O�E��[��*к�~":�jz�$���,vY����i&�y����2��Zo.2��l]�'�wi�펑A���`u7D35y�j��;h Ep?~n�P?�X}Z�&�@#����Z�VBm�`ȉ�P/�W�ʊ��5�2�����1]��K�vM��ַ���q��?V 7q]�y��?L �%�jJN��{t�R��-�MN��QX��I�����P�뱤�^��O#NMhc���N]��\Q���_x��=q�y7�	��zo^�Ov����* ��2�fB�e�5���/����aJ�[m�=~�:6�}�E649Uʾ�ClZI��?�e�Y2�/M�m$E9�����Ι�%��"�3�m&��;�Iy��7�H�K�z*t	��gV�x�P2��+��u�O��u[^fK�S(��ʩ��4mBw�q/��W<������D������5�?;oq����KA���~�C���\ ���̔`�`"c���VZy\Ʊ���up^_NO��7��6o\3��۝�J�wuw1�&��&1LC��C���q�24�3���#z![�%�⋕�����؊�6��Z���:�-��Sa4g��.��H_�9Pl�k���R5
�j&�2��l@v͹�h�,�xk2*��ʫ�9lY
ϙM�3G�.���Zr>�����kV��1~b�?��4�0�if��B�-i�6ף�x���3bS�Hי�oT�|�{d�~�,UJ 7��ӡM�b-І��27�=�����	�`�	)V�N^�M�(�3���#ɖ3����Y�亻�Ƨ
��Ue��*\;������,d�>�'��!�FK�Ȕ�\�=:<T�T<8�IΌX3��d��VpD`�l��d9��0l�%SK-}HkV\-���3�4\�d .�l/�f�˩����_�J�O�k��dXBr�xJ��Z��W��(& :x�̄8]��@��U�Duf��R�d�?��g�!q���ޒ&��*��pF�?��[o	6<�m��+� D�cl^�m���6��-�=���SV$�#��L�пEi��\�j9��E\�E�wC�'�p���+�U��p�I���CY�i�@Ѓ�0}�8� RU�{����V���ќ�PBʽ������yu��"�n�cQ�BJq#i�l���m�p��uG��L�Őo]�S@p��+�t܆�1H2E���jm��s�fp�@��g������C�r.�k��#E����n�C���Ö���<���*B镖3��J�w�$,v�B�������e���'`?r�U�u��I�`�_�\��E� �B���"�o�����^?Ku�^�q��U�o��1�٭"3$�I��%�t�G女ݯ�<á<,߮\t��,�ԋ&�4ʝ�널��V����ĵ��C���in�Q=�+���Rl���<��L�1Tl�e9`L$*>3����`�7s�6�����<��|��N�����K��.���N�Lo�M5G*��yt}�����b�xR�0�$	y�t�䞘�4�x3�Ҕ�O�㌂��0�ƥa9��l٣Xӹc1S{e�D����dՊ� a�����J����� ���a�Q��@�=R����\lՇH����6"�0]S����}eU��Mi��n ~�X���2;l�(oBAud���B��n��t:lH)RBKb�NK��n�K�ܼXz��$� |��t����l�c�-�<ڔ8S�`��2H�/`�L�Fޡ��4�4v��>�Hm��p8�(�m���'�d�A��d��j�S�5��4�:��e�n
��a�Řy�F��<�w���<�[[	F�H_� �i�&�Ȩ�3����~����RxKR����fDŧ�U�B�.av����}E=��cg�/W~�;����דv�Ppډ��Yf�n�A�/I�9���nڬ��b��gS	f9���0�uS���	�\tW�F5��%���������-���d!K�s^>���?�����$'����j] 3�$R�)�d"�=�洹���3j!	�[*R����b�=��mP,��0w���a��N�=l�Z��Ե��f��hH���%��M�r���� k�VgE��}V��gOPu�w��
mG�P6�{a���v�*������U�f��tX�M�
E(d��y��|�pc�������&�q���5t��:wyJJ�%G<���[�Y"�-��"���[o��� jqӍ������</�*}�ki �Y�F:�)]������柄%R��������R�_�5�)^һ<q=�}b�eT;w�S�A)l5w*�hEt�cI,���9OK҆l�H��!��q�ꇑ<�3~�vF��La�j�����_X��yۍK#�������@����SB�tJ����:�	�h"��&V�sZ��!��n*�{�)�8 ��������c����p�o�:p��b+J"J�Q���'AR*���x����}�6��	I�5�0@(e?�p�4ʣ���DnG�1}Y�i�բw�<jK���
�n��q&����?͆K��73�����E�.�I7T���)�Y�,�<<�Y��,`�y(>(*�w��C����z}
J0��%�e��6%�F��Vq�W��2j/g��^I~�Ό�ωݵ�X	h�b���U��DU8:�!�yc��a�n�ٖ�����4Zig[eא��f'�����B�LV���� �y(�G�L���XG�ߏS5pa�f��Z�D]j�6Sp
;�a-8B�j{iɛ��� ���-� �%ڇ�L���k��A	��t�pJDʷ���{�k�]C���/���ԓ3SL{l�_/�sI�*� ~�K�|�ݥ󨾪���bp��},1GbJ���[n(x��}�85�n|���p� |nf�s���;��j�/�ϣ&���Mt��,�sqL2�&:W����^���Ž�c��o5o�	�`�òQ��ұH*����� ձ�L%f�����;g�����q�t��sӢ��z�F�V��w��s�����#�j,JN�Ou��zsj%{��%	b��hh(���W�v�6�Z�cw���ڐ�<-.:���9����Y�e�y��z� Sa��f��D9��+�5D��_���q��r�A�ș��K�F�-%�  gF�}|�=)�ǳEDt訏�~َ����:j�?b�@lP</��^H��'��T)���YG���f��ݓ�ߞTd}��Qk3�]I���9�}bU6�#�L�"�s��m]�Y���e����с7K	��7�%��t.��p�]:~���"�YU�Fq���Z;$3��M0;�#~O/e��Ԓ'o6D�%`��Ω@�f�չz�g�@�T3Hs:>t�c
|Ğ�*�0�<���|���Y��0r�f���< d3�o,�u���K��_��`��_R�|պ���W/"  �WM��x��i����A�5`f�KkOW�O�
Q��|�n��>�]�F��"��"��ڄtUT�%Fj���x�8y'�G;c���W��6��k�y�)Nm�9�z|�H[�TI:����E)����:�ay1z�r���̨I���Ok!\���QJu��Ҙ��I�b�	4��_��s  Oa�9j��ɍ){د/c�q�8S��B�E
��QQ1Z�������H��R��O)��,���m��'-{}d~�j'T�һaG���{f��S�Y:u�2H�8}��Vul@��寏�R���{8�$�"΄�z`������M�� '!���:�0sS�X���Vv�?�I��g��N��;v��ԁ��1�<��[�>�.�=�[J����TͽoR�%#�����ˣ��K%,���S�����5�Q&X���4�N�!m[c�D̽z�.u��ckax֨��*����ٛ�n���9���t��T�E�+da�D���/��vM�WTH�&*@<*]�a"B�%Ǌ'p+O�gm0xT�,Rf�uu^h*p�LQQ�����Zb1W
�t����W�+M���c�F�^Z0v�38J�z��k����䪰|��,0�	���ٗ�Q��8���y���e�ǅ:B��fn�% �2^�&v�e/ �m�`���j(�:Xߕ���
wt;�|L�~4��)1�xk|�ܼpv����O���N1�U�ޚ9�	��u�ϰ�8�E\���9B��ߠ���1��' Ͼ?Ґ�
.ڊ�9E/m���ꘅ�YtPq�%#����/�7P̗0�:$��[�B�}�}v��f;0�"M�6�۫�D�/Iֵ�Nj�}�{�ʨ���c��B�1K��YCp�B����0bA�"�`}`e�N�ɟ���i3Bz���~u{n Q�͑80��?��Jd9S)�df�pb�?Ø�`ط� +/�q+���8پ����#r~��4�5:����Ui%���\�>g����F4�N��z�F@᪪��U��WDY�fX��f�ܷ��k�,ME2c^�J_�j]��(#w������33ڦz\������(��[��O
 ����<���T��Z��ըW����)ɲ���q	����K� ǁ�tِ�s5��պjh�gh���s	/��G@�^�[�k8�����:��I8Jk�ԯ(�k�#t����ۚS^+mږy[��A�9��-�8aި�zp�p_�K�@H�vX}��'ڦ�6�m���c�V�YlhkR9�߹!H:���VE�����8�5��ym��y�Hc1�	�x�г������}Sx��~/�QZ�x��2	�ldىp�®?c�M��ş3��&04��=��Q�"��P.!t��O�˰�lo���$��h�87@O+���g[.Zƕ�) /C ɬ��2�=�Ob؇��ؤb�6YK�/����D���nԏ���jQJϟ!�wX�a�Ļp���o���n�s�.���ճ�P�Y��ڟ,M§��T�S����* G����a�K��7�����g��:��U�{�)��b��oo� � �Ƙ��Ȕ|���98�w���i/K�����ЃQ�pJ�6��D�AX��"�"Gk�\��X2>pA��E�	5f��������%�*!��S�[�L6���W���F�쥦�Rv}ĮE���0�6����Z������i�1�Hdqg��NDb�>�9����q(j8�H����4��$$	�<�b��>���Re�FZ�0���^�ѧ��^Z�'�,��j�(0��c�GQ �����bVˊ1���SBǷ'�P�Vf�zN.�-�CN�Hޜ*��G��҄a��O}�ښ��9�]�?*�+���@��(Ȃz���9v��Ӡ�t�S0w��M�<i�?�zb�S�j=���μx=p<��m$E�
���V�(Cq�)F�J��?O4��Xx��䨌hAk�9�PT:��]_S�1�l@�ҏ���{���0�CN34A��_��iP��t�e� �|�!v}̶�;��?��E�;4l��p��i�����c{A��MOO�����QMp�,�?�vx˘"&\���8�Lw�V�ď�9j��\���$��?�R�����#�4DN:����L��@V�FQ�}C��7�7��� �M���UM`�� G���Àl��O��$-n\et\v$� O=�Į��'�>�Q�o�5Q�X��u���H0:��?n���'�KXF�,�V�V���<��a�=q��ٔ�ŘV�|3����C/���ugr�`ڧ�� ~� u�eyC��=l:vi���|���`��l���� �����r�͕��HíMFc{���]�̓!�9��Ä�ƀ�XPM0��i��ޯx���a��ש{2f]�#_���{6��1�ERm�%(�G�c�H:8��l2���yWEKGC�3�T>��q�� R7[�!n�P�#����Nm&Ɗx�@�N��c���,+R����B�ї'��qCw��e^�@��4��\!�>Y4�v�^��q킛�rL��XS�I��?\t1=��ƭ�	(�L�6\�R�nr.T���#4`�C��а��_����}�>Xz���
���9���Bnz�����%�FacQ���Q` 9���A2���3[����Ҧ��	�&�׿�rᱳ)#�9E]U��d���߫*��ܜ����Ԃeǰ�J����g,~Q)R�T,�8��� ���t;zE�D��\m��&|7�O�Vڕb�r��Ԩ	�� z�T]��g��zG����O�>���cj�w �s?Y�K��c5�YĞV��	��P(( ��T?pJ�s�Un�tCtC#-����%�zwTǕ��ΑB��j%�������m(f�U�l!.��Uj��r�}|sJ�	m��bsEy�b+���RW��܏�4ɒ�/M��x��D0�ν����a������j��)�K0�Q:�"����F��ϵ�B�����9�"���u�bQ�}��!�T�ޘ��<5��I�a=x�R�$�XY?h)�Mt�9���o���"���<�]DJ?�HY��~��_NO�����kN�����bg0�UD�a�:;iR~��51;����(�W'����`F��,��=��+�6{Q�җ��U���*
Bg��\IX���O���q���B�HlO�Z�I�K��<=�v��Pr��o�}�a��O��je���aW��������8@^�7g׉�Ã�B����]��	�=Ԟ�$H���y$���B����x�>11��«�V��4:"W�de�F�g�D�2�m��]�z�B�l>*�Ɍxus�)��ϫ��p>5��z}s��a�`�b�BUȶ1<��R��غ���I3"���u�������|+�o6m�z	�}�h(3_�'���x�2ϸU����Ҙ5��m�j&��W� 8[)�eC'�'4�^��@���0jjD�����H󸨅Mzl�}m�9����[\`������^x�`lGK��	E���������F[_>��:)T��"����딀�%��R��S��2�f����}"C%��{�p&���"�"*T'�"
]���13��%��'Q~�$w��HQ~�#�	��I<Sn�h\J�eeO�侹6���Ciu>j1�,��N�~v�^�p]�tt�KL�v���/
������K<��}�GZ��5B�͍�(ln��o�<����g`^��?��@��2�f���qq33f�$����i ���P>�2��p�N�@�m���c<0�\�e�a�h���B��*CX$��z�s�8�#';�NdT��d�� �n���oS_!���y�����i*f`�Ω�\���!��:Rޯ�@�eo�sd�-W�t�>������D��\؍ ѩ�Inh���mZ>�c"�@��sדK�ʡt2�."�1�����So��SE�UIJ� tR�:>�կ���uL[��rc�4��7�q$�4r���9�}�����ۤ�p_Y��ț�We�!����í1�8^�
��2����_Xq��q��Rk����= T|l]~���}L&Y-_Y$T�q��������ǔ�>Jl���f9羓 ��+�ځP���Auũ@Ї-xuH���tTt��eCϳM�2���àw��������G����k�[�T��Cg��<���3"Y���3�G/{8m�־ćn�3��׻��:U.�##P���R�e#��~�%H��ܒ�D:c���m�š����FkuT�ơ�k����{�^/��8�5�*�@��"��nHBN����#v��cP%�|r�@ۙV1�ã��?��Mb��(����6�O֓�W�����#tg�{��iYa�W�����{���%.����:5�q~��nc�g2o_�ra��c��PT�羅���))M�{S:P�0�2�
.x4ע�
�}���Mc鴉ؠ�˭$f\`���޹��Eb�ߒ�L���<^�`@���x]��*~d�{����̓~��g���@�~�^:�g-��,�O��C+�u�����jk���DV*��1�\l��C��a�X����m�eQ�k�#4��v�Dx_��|!)$��sB�O�z��c��7�@MrrD���E:�1ӿ�f�_������t�]S�2z���>��nw�mb^
�,�Ze?��E�C���VfA�c��C���Hd�a�iӭ� �e	}��vj!��������U ��D2g�s��G���ñv�y���ͯ6eaQ��A!g\Qu=�0Ә��(bΪ��,�?�X��V	��g�X/�� ��Z��A csY{Xޱ	���^`X����Yw?���Ya��<��~���}�
o ��

���ͱfLL���u��� �}���	�qϣn�P\}��au���p���U��\q����e��Mn���;Ǔj�:�>^c����o�4]#7��5]6^5��'����X�4��ˈu��!^��l�[�t{��F�+�:;��ܯ)96�>Z�xy٥,��J�������Hc��L �Zy�a��-̤E�ߙ���q ?����̝��H|�OA�2h�*�7v��}�>���Qmx��1�*�6IA�X�-��|�貤2{��?��s.rh%�����l;�-߰D�'3kQ&�̻\8�.�>µ���*��K���Cq(M
�i*�$+-�_2���(��3H[,==�>(/�F:P���j���i���P�."����I���ž�:7������mŲ�Eb�W(A�ɍ���+߫�$A�̀"D�n��İ�(�یZ��^0���%���9A�5���hjC/�^��5A�8G6	k\Y���H��P�����,F����(n[&+VT#_��-�(�\�N"�CY�6��ePV�z�$(�_�'$v���G��2-��u�<<�qy�3��S�.�P�b �����^?�DC��Q9ˬ���I�=��o+,��>=�V�>R��"}'������k�ot�m���=��8@�ӗQ����í�a���<8�<ZWla��v{a�|zKu~�ΞO�_���ݒ(n:X��l���g� �(^�����H��+ �eL�L
����Κ��c,�ϊ�;�=����u���@ w���i"�,4Tm��h� ��'���P�)O��v�>��]R8�ݨ�q"��a�N"yGX]vh��8����g��1)�.^Lw/x���3gYƃ��Z�]!�Fe`�m;𾩷�4��� ��`%�e�8���8cM	j�U)�(��.>�a����=n:u����VB��>��}��F}�,I�����͕W��]$�!��I��nOb�-P�n��G`-�t��)��_I��T�����d?��M�lES�=��ڇ�-r�0@��b�(�?~"|l�B�ŵ�)e�A�d�����̝�H�e��Es<�j�ލ�����J�K6���9�^u<��j�����FO��}��QR�(e�SL1�����|mf)<��o[�ڠ��[���w?.���	�0ժ	�D�/�C�"�qz��Dp�%�C���8Gd����u�&3uz���瑉���#m^ pd֖�걈aܻ(��e�*�G�+b����k��ʂ脗7B�Z�)/(N�����5�ڄ��՝_u����L��ϛ.�o�Ш�CPo*C[5���Gc.���<���U�7��6���uF�H0���h �����k0�1�n���%J�Ȧ�'�6V���n�r�	9���Ie��ڻ��"��]4*��ට|8+3D�D?�4z�&h�Ͼ�[
UL���Ws���hx��Mu[F0��j�a��������A_��MD�%&��c�c�:��'�C�Fj?��3�Ä���"TC���`�		�5����.�������������w(�W����r"Fv���nP]����>o1��؊a��o���s�É�����js��z�#�sOʴ-�&�D���2>\^�TS����A�y��rS���Q䈚�����G���=�3˅=Q��W�M��͸@�Omy�b9�j�A�Da��Q�/�<�m2Ťf���3&���~�	��u���~&;�&D�!�O�A����t�������E~�_Na���A�5����q��SW�c&��m�ϐ幵>\z���E(����\&�6��Y���2m s�h��l�lG�"`SE��@�U�X=q�[ߚ{ɾ$�EC�-�˴�c,����n�Lb%��-1��%m���ӈ$�����n�>�vډ����	Oiȹ/D�	�Q���o��}v��!î��
�:i�=l>X�;�q�ػv�(��T�}������w5kV˶ ���$�>�y3��	�f~�^�D����
~=���[�++��u�3Tj��Au��O-�-
����\8�� ��zMn�J���^HB_+�/ӯ�<��h9Z/ZG��6�1�˩P2����V�2e���)�ؚ:�����?kNe\CQ�4�����r�6����t�td�b6A)zDo�4肚>��k��9#g���!0������ŋz���6�D(�CM�JB+c��d�h���UyW�FO/v�{��_9ģ@fEw�]P�N!gh��e��ֻ�l���(y�ꏼaמ���1�e$�(�h{AN�	 	�3��N�I����+P[�f�Y���ɩ(����vova���n������Q�z��X"�?��=U�@!��O%���/�R�����4�i�Հz ��h4%B��H�����ʂ
^�N3����Iw �����]zh��
1k�@V%�zc���g�9�e*^�/e��u�1z�:x�PW� �v�<�s7CD pW" ЂNBT���~]�VRx�� �-^.��Ջ�U�d)27��Fؽ�"c���߫�~������6��tR�ގb�{t���,6����"}H�7���b�i�h���X�y��\�*�:�~�(2Qc�jLGp��K�9K�%Xi�����P�����_�M�q U��|����B0�|8��YS�wN3�G�T��4�-3`6��o�B�f�h���$��-�w�?^Sz �М~i�9���8�i
H�z�n�A*����Ʋ@��+�x��;�u�AHOFbW5�iJ��*D���5 ��B�[M��B�`���@����ë]�R�T��m4��Ոc8;Ȉ
Ĝ�1���^�6�Py�n�SS7��3�	�׀z,=���۔7�j�7RNt�兀u���<'��e��IM�j��}���:=6�α,`Q���L���p3O�*���b�V�,Ԓ��q���4�����ڐ����{���y�˄�YB7�w���:O%Xv��%Dn��L|����ڎ���Yp�zT˄�"���Ʀ�nr���5R�f���k����'�·���i{����΂�������O(�Lh5�w"��*���-�Ξ����7g���O�����6�w��
����@��U;m�M~���v���p�)G9O���%�-�TG��v���%��>�L���e�甭K�n�����(���?z���-u�c��-�����K��NJ��	�x��˔�..G�p �Q�8�a'~��.��*�{�jz�()�(����Ryqs�9$kv�$]%)A^��/���y������BxW���nE�;?�{n���uX�vD�2H��:K@��`�N�D��GY.�\x���S�x�5D,����F �!C/�3��vS�J�a�0���@�\� ���sk)�5�Y~�yO�p�	�R�aby����!ZN��g��ME�~L���\���7��T)��������C����û��{>ћ羄����O�B��H���y�������)鳧v��rA�H�w���>~v�"^X�=�����g��)
�a�OW��bW���%��	#���Ҙx�S�'� ��)��s�?^ <����^0d���Y�N�I��q�s~��Z��V��ǀ�#������5����	��{f�z�ڟf����Y��	p�U��#�E�ƹM�mĂZ�����2��X��%>�6���~Sy�y~�im\���KN�M��|��횲��5