��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��We�����9�b�vI�2�ȏ�����
G�Ӱ���L�`/���谙W���?�U3M��,w,a�*= <kG�m@(�I���б�OTc�]A�\�C�/h�>�����\a�1x��M�%��ʼ7���+i�N�.�q���;��4�n?<�ܹ��L�R��][Ո1Α+����I�\����=�#�.C���@Vn�#*�rN�l �٪n���\HI� 	�,Y��LD��d�\�D��W��
�Rx$�[d��SW�9S��f5�o1� ��U����F��ʤ���v~R~�<�����zqq��^�1���T ����Z�*�)��(�c��V�6Q[��a��L��i�Iܘ�7�W�����&��iȹ�Nz�v�aǳ��X�������;T-fG�w�?�����,�ڄma8Р�/"%pM�\>:h�����·���<����u����m*R�k�:��icX��m4po��3�#$�묾Ct4&�dҡW�6��ϋ4'��o�.����*݃#:
����}���1�����[E)0���mR�-T�"�-�2�X�JG:wY#�����c�A-=7�x�+ۅ.d[�κ��a3�Ym�	2�#w[��sܯ	'�i��1~5��}F0=1���z���Q�����?�55�W��+(����s9"%�n����	8A��GG���?}� 
��]����K�Ш=�P�Ccς�Y��`�p���{+?��Ҥw�Bʐ{Ў&Q���qӼ��kb(u3�*�,@�!"��DqKQʄ7J-�E����8�rԢ��ьX�0����Zu@�I8��fa���@�^c��k���x*��i�tpG��&=4�T1$��0t`B�u#��h����N�,���^Ѡ�L׻g�6�D�'°9ߙvܞ�2_Bv�>1X7�h*]�4��`FR4�c���s�%�:���r�P��vR�_w�K�*�����YT��_��ܰ �qR��|
��hS�>��f�0�a�I��h�5Q6��ќJ���jp��uR����-���v��F~�]�_e�@�k��W�d0��������䳆Oͽ S�	A�y�!1_N�:i{�m��6��]�-H=L��F�G��
�ʗk��f������ �)
(po1���?�TR&R�T3�o����_���ȿ��5��W�b�����>�7���g��dI�X�g������wm�P����{�M����D`q�ZR+���������`��������:2%6>*2��],{��ނU	�c�ay�j4��C�\۴�	,	�P�B��!�\JM���Lf��q�G�����(�5]�w{8�E�f��Ǿ�,��Xb7w��_�t�Rr/7N( c�!_����>Ğ��Ь��4�&,�sM ��"�`�R��f?V�{�Q��Ey����o*O��v�]9~ԨJ|�1���pϣ����hր$��|url��[n�	>ۀ�1�A�Icq��iqqX��?�j�%��&n~Sr�1��w"��Yh ��)�(@et���HE��1�P�sW<�E���ݻ�)Ñq�����P7�����, ��)Ll
pЈ��AH,BG��G�jO�Y��c
��=�Y1=Ƀ�����*�9���?)��k�.`��8b?���K>aO�_���V:��G�-p���_��F�{^8��zg,Q�U�.�Uv6v�ܲ ��8��՚
E��Ku���_Tf�V����<=,r��[u�{*��������i9����L����ꪭ1x��������["�V�<��{�ϭ�.+Y^����/�7$V ���@E�ŇGd;��?D�/�� ��j�\gzbD���\��eu]^�i�(k$���FԐ�?�凤�#8�B���S�n,(n#�Ќkg�޻��=��}����W{�����ɩ!��?zY���o޺,@~��<��| ��Hoꨑ�ޅ��w��x(Ҫ۵�܉LS{�(��4Ox�2��(�p���P��n�)k��<��&i쿲1���D���l��.�>�Co�z;� B��c[���g:���.�zÑ����e@�̩/����.�x�N
���'�1m�?V6	�Q���S�]��}�}K�'ߠ8e��G���q{GD�<����tfibp5U��!(D�ں��_Z�ھlO| ��8b��(�S�9},�U_f~Ji�ׅv8�"�
Y�����Z;��|%�n�$��LDaA��T����"_U��\_de\[�De:|ő�9�%��=s�b,������y���ndڜ���^�~{��\��x_N��Q�4��h����3م�3�q���Y�ڼ�	���*jl�>UvG�s����� 	�-��~��|��X�b�׬�=ϝ����u \�W>h��&<Z0�A�/��;AP@��r};Pĺ��>h�n�����*�^�t��2���ՇJ��^�6���!�OR�`wjOe����a턋��ֵ�g/�c�!���,�	�Nq2�;�����~�j����#|�E�ˎ�v�$���f�/,��n�*�N�E��Ή¶U�J�������2�w��u=#ȅqk���DŨ�~[�gjӮ�q�7լ:@x��&�8�A�>����0h�O�#F�o�� ����f�O1t�1�F���/ܐ��	e0��n��7�pZ9'��1�$��&���J���g'"�k�B��|1{=�����i�=p���krMo�=r��O7J����)�]��*�D����Q��R�N����`P�~�,~�D����h�݄cv�uȹ�*��>�n��5nD�,h}�а?�Ҟ��/W��{p�gH�z�U1�Ë0�1k��P1 ��N�Ӌ����Ռ�g���~)�	 ! �7���b���V�t/lVư��T�5�������Y���� �-b���=�O;8ӹ�`�/��&p��=����׺	�U�p:�ْ���� F�0�8N��;eO10v�%(�t����A#�6���\�?�fF|�k��?�r�#{�K�n���Q�!�� z���������Ɓ��x�s�^��f����)F}����A��J���3�X��Cq�/I�ē{5�L�(�����{�u��N~��U:��ߟ?��tzߡO��]E�%quj5u�1�h<���,�It{6�cf7�эn���٢_�&vA ���>��>Gr����C'��D���=�(xϡ�����o
� ώ>��a9 J<on���O�C�9��x���g��c�?r�ͱ�`���1�jVI�B��r�jy�:5�qy]����ސ���J�)Q�z�i�u	껞�{�U�hJ/��s]�İ��s.ån�q��P��/�N�5�Ŭ�
�b^��ths����%�r��z��;L=��x�D�@ǭM���GK�;9�����FK������R�2ox��n�á�!��/ſ�<鹛�[˻�`��q���e�2�8U��]�2R�9|b��H2G�]�Ĺ
)2��H�7����~s�*�K�VUvQ1�R��Eʥ(b�Vܱ7��b��@	���F���G�-ZM/�Pl��g5����x�=)�!AŦ�LA:���0 ��j��(��[̍���ܝ9gH^��[���k������r:�O����������>Hg3l(s�����W#�s��0�_��Dn��t-�y,Z9���oE��36��/F��7����`��WHZǥ0)5�@Z�M�ꕀ�Ĝ�_��ϸ)������y�eX-��lFP@��/q��B�~ǈ"G�'�{{ZR�ϟ �o������.;�������π��H��q�&��s�Ѧ��j���rj'��h�~`�QHw����u��d?��t\�������6D��?X�Rj����ĉ�oUw�pX{X�D�Q�WX�c��[�w�L�P�>㺚�� �)�~bZ�� &�5��A�c������u'�ͥUKk��-�K6,�O���"��_�y1�	_�y�J�<9m�s�Ż����ӿ�?�{ųu�;��������I������՛uF�P�č�郅�$cT�mֿaZ�ׇ9��@z:�Ɖx4�f��.���{~�b����h�I:�nu�E����x�J]���l�g��{�׃2Lp�,��kV��IQ8;� a��]�~*��_�8���p W����t�n��� 7,N}�/j��Y�h�G��6X�2��F��7-:�-Y�{���IllTs��'�l�z�T �u��d�q$��x�0�P�H����H)w u�� �㸇�A9E���̟�l�����L�<]�:�XS)'I��h8	���[kL}cm	'5���nX0��V�xd���M{��p)�1U	��s/9����F�⳥���Z��C=V����L]z/{�[�� Ur�6X2���³)S;U'`Ia��^�>�=�
�h�=�"��O�C�z��(7��&�t��0�l���U:�vɶ��;R(G����w	-Y(
��O?.�ٱ�H��Z0d��b$��l���r��+��o;������C8�+Ɖ�e��e���Ѝ��  :�{�+!���ȃ�#��z���Զ\�_@BeJ85;}�?㨴�� L&gt�*��mxrl�\�$�sH�7�(Nl/5%�#ܪ�v0J}_O���,+=��z#.�E�=�\�j��T���4ŏtvR5�t�p/ӯ�	p�R4�@	�卿�]"���G�m��VDd0��w;�d6�7�!
А��a�/�5�F�{R�䟩2��&i7C4�%^�⓽G�G��cc�$�~�7j�Z]�}�x�5%C���G�q�jM�T�'2�b�ʭc΄6_����Fz�-�{��~����[����'�-&�,��[���d�+�����V�6k{��ٝ��ڻfw��c�[�����~���Y$�*,�(��=:�t���Y�E篡0���<�KVb:�B�t3G^{2����p�����W�hb $~����!�Wa!���L���s�����f0����OL-�O���o�wg1��� �V�y�'�nS�������US�~�Z?3�a	�%��X�������Soc� Mm����U,<�MO�Lim�'#����l82[���!��U���C>�\q&��Ӈ[3漆3���BI(D% �78���K��M�*��>�tǒ84��0%��cq�&�����?�����iQ��9������?3@�� p�w�)���G�v�X��%V���A^���Ѷ�ht��3%�3E�~���ai@Z��ȴ]:��+t뺑䭌*^�a��G�7K���h-r�M�DF��-���q�`A�1���hR7����mgw�<\����?L����y=t�FN�o)��Ff���ͷ����ԟq}���=����B"��uVn���$�� ��+2?�>r�?.D�/XU*x��yἪ�Y1��ƔEp7e�W�"ۭ����$cp� j���b6��~Qz��ӪP��_���1[Ly��&�c�)
Mk�|7����NC�[�Ń�^%,��u�«O@�ZJ��,�]w,20^V
�۪�k�Զ�N7���D�ȗ�s( ���n�oG��� ����C-lj��(��X��3�V"����I���&��5��x<��P���C��0���p3�G�y���2�"y�˙Ա�̄���/�q�O#�����^�uɤ�a�z�r����c$jP���$�SI���_��~�!6�)p�8"��=gL�Q�/��f�H�5z�/�^�-ټvqH���A�i��rWX��U���S����{�س1Մ>U�슶�=^D@�5DF�:��
��3Y����o�wg�g+㩗�s�w���։(��dg�w���#n����fܑ�q�?�j��g�2za�`)�ǵ�_(��]���׹n'�ɹ�7���H�=0`�;�s�M�*���w*1��+��+hv-��Yp�2�~�\m21�)�e1Xݞzp~�pf;���bV"�E� �pCv����P ���
)�C�����HS�C��;�ٝb�P&�[OƟ�2)x���RgDM��$�t0�Ҏ�$.�?�N�����vHzwwZ/P�����C����I��$^�8v5��С�C�p&�^�4�\ �����䍾�HeR�����LQ���$M��=:992V����e�3��K�3#������	��#3d��(9P]�%� i=��Pw�t��k�����O�����="=��lԵ�$�n�UB���u�]��]�x{LR�0ʶW�o�-��IL��>'=��|���[�E'�v�lt���g}�`�-4�#�RA9n�?�v�$0��KԜ�U�z����}�v��8*G�[���N�J�#��	~�1���,��Y\co�EX���r��s�����Z�<>����%�8����n����,uj$�D�_u
�������C�#�@���^�.Z��9�iӁ���n�Q�7����]('m#0�E���T+uD�3x�iL;�K��]22R��@�8y�CW�ё�lٞ]�#�rހX��h��^�8����f��0� 8M�_�b#�/$7�o�z��m���w��$����u�f���A�	��S%�d��co�%���Uk1��p߀Dt�X�Z�'�RH��;]���4kp-��Q��1֤j,�Ew���c@J�;/j����5�BX
��d'dX0�漱��?�I���9�¿G���4�VrB�t���˿U	���pTiTÂ~�m�X���= �d�;����G��]A�J������>���*]����-�b"��^�<f֞�-���f��~ӡ0�i߈��Jx�p"O�'*�XH1VU`njY:��`��.k����~'�����("��	�xv�s+#%�Q�4s{\����i��o~,|�����<�m^��F�����6�T���[�CA���kD������N���y#��k�->����D���L�3�ӏ�(ߜ�����=��\��i��n��pQe�OIj��X�<k��{��@ȍ`��W��])G�L�8Ӿg�yAw�LG����_}�G1�~w����bx+��?�QΫ�m|){��U��
��lzE�{�����PE�hX��Ƅh�k ��`L�
T�%3ڹg_D_��QjZF���5�e�34m/�>��Ζ�C�4�[�4�c�(��<��sn\��|�m D+�m���>���0��ͦ��+�G�����kP���&n&��:�Me��Kߠ&����ތ��Z���B_�eRh	Pfŵ���y?p�Ӂ�վ{���h�87��[~p��}]����c�����"���M���w�����k�?غ����ɴ3B=��#�X�"���F�ǤN9�0��(�q���~��z�R�
h*x��<���VU��P��s�\´{u��Z��ӄ{������?y���J�����佼�̗���R��P`g�����ϒ��!�E��Z�#u�����v���
�*C,�������O���~��4m���n�{�ɬ��Gq�����ژ��t�,��U�0���}�'A*7_�&�}�x���B��Ԭ��_��t�XKZJ�L�~�O�(PV)\rC3yͭ%n/|�j��̗Y�ƣs�pS�F��-�Ͷ�Zp�{||�g8��KD���MhA�-yw��e�!�����#�M/�3��z�-<�SX�i&E�W6��8����|y�W�����&�i3�B3���~
z�/�G"���
��=ێ/l'�y�߻ndE�����
u�hǼ4G�&�8,���V��O+[�����s�ih��~Y�_M�Z�E eg 'f�w����Qf�{�ؘ2��ň�������J�����.b�rwx��!ج=��68�8�$3e\~�L���2������� %�ie�F!����/Ch@���4J
�h[�L#������=�g�I\L���"�sc8�m������w�����[uFq�����щ�fm?*ƴ+�\p<�]�o�^���C=��Q�x��e���@��x%��]P� )`^d"�C�S�����q�v|9��3��S��k��k�.$���T��*�^�����盐L���]�K�`0U���m��,�`��3��5��L�(��A^����m(�0�UCY]4�<������;S�����|���v8��!��s�N;���o�hHb��k���:ƘGP5�$��ި+�+
/��fE��ٯ �,�0Ή��g���z�Հ��2U��]�B@2
�)��qu�Ǧ��nBQT�?в3]�m-�}��QbT�:U:E_HB�i�/�=���O�,�?�y9���۽Ñ�����A�9������A�2g�T4[��9J�r�Þ$�H��o땑>g�59�}Y⬗��H��!^���g<{�pVӛ�Dyj����7v��sà긐H�0�6����MzL0{>��w8)m�C�բ�^	`,��c~� �9��8�谉��tǦ�oo���Ly�+Y���B`[C���nK�v���m��j�D�s�Y�͓�@�l+ q�-�f��k�U.ud 0��:���ۓ��76�=kg���{�}�_�?�Ҍ��n5e�w�V�<D��������� ��_)��1Ϳ4���	����Z�����s�n���-^S�Z��r���zRuc��?i;��RS�lωS_=�$30�?�|j�r�/�#C9��ߧ�8�4~�%e���6%̡�%� e v� �Ye0,jh��?�RT��2�(^��9���[������q��Rsf�)U�K\��u��ݫ�n������q�(DAM����-�W4`��;3K~pZ���g��B���]�dc
`��r�SШ��̀�Q?i�馠�����"2vg�A�b�`�Ə̭��ng��E�-����-'h��m&TLI=M�7��d0���Lz�E�QgJ/d���Kd��߰6F���bH���+�ƕ�4�����y�:�.4�����&C��ZP���?�1��o�oR�� l�=^��=}L	V�ȷ�B�4�U���s=�ml�h�����yQ��� n�A��e��>�"�����r����
�{��ŋqAa��_�h��$�(tk�Y�`OQe�7�ŕ����L2���7�@!��#keS��!��Э�aP����i�����b��vM@�~A�\v�gu������%@���Gc�kF��3�MC��˭�����E�E:�Fd��R��{G���l���!WȰ|�h�B�ᔜ�ϥ���fQ%@t��ܢ�C�Y�ֆ������j���]X����v2�&=�Z�H~W`���]�d �F���9)6�_�y"��QL�Q ��/��u&�I)�畡�(��	J_��W!.�{��صO���g�|��STF0;����6��aĄ�t�	P������!9�U����x>$Ӈ@0S��:(� ���F�؅�w�8]�*		wӿ$���m~�,Q�Hp�qhW�,-�*���ەI�`͏�X�� hX�9�
಍���P�,Y���:A<�p��;r�4�b�b�jp�:�80�ܔ_Hp�Q����e�u�&�' �d����uᆹ���qV���s��2M�E���I����O�"�.�M$��Z�نJF�9{y��0��f�������v*�r��-o�^����AXߟH/@�E0�RGUU�u��D��lG�>����.���j���U��pe���F��}���C�-s�⨠�#�U ºK2"?&�-ɝf5Q�j�94Y��=2�YQ����[1����wI�w>~BB������ɕ����72�a=������fD��x4k���Ov��׸�C�&���R\[V!4�F��/�o.���Mb:w(A��!ѩ��S����~f����ר"�}�)�C-i�,�Iɵal����e�QF~������V��3�^k�`K���B�sKJp#]�(G?�L��Q���r�bE7v�g�}ޡ"����p�оH�JY_��11��s2Ro�������x�Ol(��Y�G��*��.�m�.����,��񢪨q`��� {Z�^�r/�1b���^v#+�5V�.t�֐���%���1�z��n�o��m����З��x!���aw�Y�{���あ�g��O�d���$��MW���Z�L�-Y�Cq��I�˗d9�R����S)u�A�LN���i��/!T2��>�?ѫ{�����l2�� �<\��z�������F��n��=���G:�Ѹ�Xw۩d'Z�,��J�W뇝��u�I�g\i��o�&,vґ��_F���7�j��i��"w�=Ţ���/ڧKu�"��F^v%�Q���r%�U��d���TB�)4����{C}$��/ߘ=Y�.�z/�m��-n�r/WOu��G�X�Nd�h��x���V���z�h�������dX�6 `nW���G��^*��F�ܤ�ƻNG��	�$~@�1)Ȟ����S��6�#�HH����W��.c�pT�]}����YQ�<e�(��#���/"{�Z1:���&�n���q���+4	���+f�إ����f�ǈ8���T�g�p(�v"��[&��j� rR��8~U��eP=��ۦ�3q��V̌�CNנ�{���G@��߆�Y~U0��8�(�A �"��Lt�m}���D�X2$}��q�g���e|q��-v��ܞ�Q~���>q�����[�q|{��rc��=v�R��尺R�*<���ЗҐl1����Ʒ��!�U�y�ң6��� h^{W2+�J��R��Jm�g�(Ms��ߓw�k����fQ� �=�93�m����ÌJۛ��8 �G��f���0�p$[5�S`�=X��nCz8�Xr�1m�3� ��'��J5%gw�J4��}���D�Q��ׁ��˝[Vd�_��R��K��s�n���"��b�V���k4Q��-���q[2mU����i�(�<��T��t'�n~>68/��"���><g�d��4�+��4�!�%�:��Z��������X�~���K�r�m��<���a����&{ۤ&�i�amL
AqG��$�{�1��,��g���IT�C�c