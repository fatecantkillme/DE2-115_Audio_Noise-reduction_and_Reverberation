��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<i 0*j�_�;w�r��nUv!��i~!5D"yl?0Ȏ]�?��#�p��`6��7���7�.SF��+�5HB�l�\�:`�X=.���j�!���@��,��w�O�d��v��gS�O�:@�(l m���7�/A��$@�х���A�n=-bo�����l�#��Og6XxN�W�E��YN8t�G�Tp ��#gMt�Y�k9L+�?8�
J?R_���5�����y`�M&�2��	ٟ5_+l��D7��
��J����7�kU����Ց��!ū�}����w��(A��3f�b��ɚ�2a�qpDT$ڼ�EuS��<}�����w��@�&i˩F4�jf�Y=�+���I���ofl�R$�z�h o�cT��K>��7f%A��O��>���κ-;-R��L����W+�7Ià���Oڳ)���H��/F�=ځK�h1]P�I�F��"D5��*wQiN�������ey1��H<�@�Vr@
��&�Ϧ��9-��B�9���E�+MY�C�nEIX�+�!�ʫ�N�~�i5�I�=Kf��lZ��@Q^s�(�oI�;
Y�S_���ۋqǗZD��俄��6����}[[�+�������K���\	.}�Ή"���#�"��>Tڟ�(�Z)�w%�kg`�3�u�t��\w����j�Ƒ����ݶ֤��O�/�J�F�����J&�ܮv�줗��Xc[�� �r�4�L*5)x(k���)��+��n���R'�%�n�s�<��@GA�Y�i8�*��ö���I@�gؗƛ<r��"�����rG�Ed��*" �z��76��m� �V�#������AƷi� >�(ղ��Nc�,���I:'4?\��?���7#��9!���ur���e���Z%H��~E=�w�%E�+<��
}��ވ�m��Uhm;q^+���������Y"P�sPq�۹�oM(�̷�T�"ی!���~/b���X��׈�\���PgV$ѐ��R�(x��`�j���y�����|�[�
�]wX�nulW����t�rw�� {sė�1Əpa {[�y��.��$�!��LL�u���^;]��0��r��d�Ff]ݬ&�-��d�#�0����k(��K&�b�ch��J�]�k;K��0m=M{[y�*`��ڋ��}�櫃�j��e^C��;�T*ԛ��\5
/���0�{�a�:F�2�|����h���q_����+Lg����"VT��No(�4�z2����F6����t�j�)�مoOJuϝ���\��E�"��vN��]�ȧiz�z��.BX,p��U^Z3�g,�fyh�Z�� ���-�[K�a�$!SM?>Җ����&��϶���Ͳ���$y�	Sĥ��~�v�*�L��ח�[��aLS�?�
x�K\\Ų�Wߐ�(&�ϔ��}Wr����^��FF�|�����|���)�N���a0 ��E�����g3W���\�E쟈h�^�� ȞE3 Z@*�����Ќ|
�*��$�MQE
�r���X�o7���:B��&���o�|��nua�-�CR��*�M��-�,�FÚ;hB���$V���^����J�{��+��� 踟#�X����L�����%��o��g�X(�EZ0�	���E5rC$��q^�m�
�6��P`�'�5r��ځNL�rE|�/������+^^�,Pq�J����C|YG��"�	�ч����������4�/�KӠP�:�f�%��Is�iBG!��Ψ��؛�%�o3�0�#Y#�M���ؽ��m��7��$#�y���%.X�U�s]�tw$��ּW�k��1�/`��Pi|��g�S��ͬv�Aj����5�Ǟ���Lw�iFE���
�<Q@���f�ȦPJ�ģ6^pq�4gFe���YD)�F�)��.n���k�O��9���)��u�G�\��>�A��aٱ��9�Xj�|<8��{�g\�Y|���"Dk:����1��#@�$�4���h�<I�4u�+�1�gBpw�r�6�#�W����k�Х�!���iN�WwP��1��ͬ���i_�{"��k����l����������!��
�ފ�+�Q�8y��q�|��+���+>������� ��}��/o:�sP2�*�(*O�M�2A#ӯ�@�q� ie���g���E{S��uދT7$ô����JZE@�꿿t��Tm�H	�x�*�;��f��yƞ�'��z����h��{Q�+�*��������}�A(�u�@�a�Bt9�'.�Q��:L���O�����2�Y�Rj�J�������q5L�{�Gjt��n�C��,-g=M[��>�1_��O��tveT�#XkT�𰂡j����~���~�9�x�P+;���j8ݐ� H�8���)��
��Ncr�%M����8� �4۪N�ÉW�����7����8��p�:%���Z0����<z
3���l���[�Y( ��5^K!�)1�!&�^�ňT���MQ�x�|���}%k�x4 ��UbVK��M��$2��g#�I�Im]�˺\:<C�7x���F�9	��Nr���97�r���'i,!<+�W��S�6ѵ*o�]I�i�XV=�3=�\����R�Lʴ��g�xbX�옿����jĒ��_n���蚝�r��ȑ�(��g&d y�F(U���:�3�J1�xS~lp��%���:�{6.Pc�I��{�;��tJ S�m�Ct�=�pi����$��
�ʄ\��'�J�ܦ���b5�9��!��_O�{��1�E���F�鲼���
"��E� �c�Boi�faK�5�0�Fi�==-mָo�3�YԙR��55�ը28��O�1����P��2�˵�o����^0-MLX���ghLA�Gю��~"��������q[�i�Z3\�|�H�O�LXr��s�P��\Z����]�=EG0*7$�7��6��G���GeV�� ��2���`�|���aAD�0�zf4p�=�+MW�o(���VUm�v�2ŋY<���	����<������C�+(sFk=��@:	�_|IW��r��7��6 ���g4��P�/%y�p��/,z������	��9�l�M���5�p�>) lt�=�iZ��_A^�������ت�&��o����p�&��^u�c�Ƈr��*ճRe�l.�b�c. �.�Z�<��@���<1�JF����|"�k�/i
+����d��=%xQ_�M�d����9u��Zw�ڗf�����m�,��k@�� 7&������h����$NU�vy�4�y�3�>t4�G�N@D��+�Ь��o��|>�8$ڎ��SW�I�;�<�nyd9Ud���o� �nd������E�8��	4�kă��6�vw����Y�>����¨%X�L�98b14Q�2F��f>1�Ly��4"&:�N������,|���r=���O�NXQn&f2G=l�V�@LD{tl8��`5Y����YW��Fqj��~.>�B�$����6�<�n�g��@q���B��7Wl�P�����N)��
�
�((��� �il ��"v+�}�� �a��˖��q�k����}j�`>�c?�5Y�v?��ѕ��P�hw�4�H�2�p]���hAc�'�����I��S�@�a�s�o�j=H��	Xp��x�K3��*m,�G>����1�I��]����� 1�JL�|�θZy3)��S�=Uc��t{���}�7��K�sVw��?�s���pQ��~�+������%���S��%�F^)y_7w���TեI����#W�u�L~���<��*���>�縰�g޾">)��CP!���n��v p���Bv?��fa5�,�%���/��h�5N�Jj�%Hz���xg5����3�Pxq#��L�r�>U`��-j01��!�s�2������n����B��E��#RTI���x�iSYN޼~���la{�7�N�u��0*�{$ens�3} ����(�.�-T�b;��XC��]�SX3 ���z@�}.8�3�>���}:��� ;��3�f#u䌳��,q�*�A���Hu\���F<���B� �%��&KE���=ħ�X�Tڭ*!��;�;��2�>(<)�r�����8�	Hh�,��##Ͻ���H�CڸNJ���#�Co �Z�>ΐ�6�{��pBÓ��&�����-��E����$NSQ �s&ZԪ*aU���B�,|��x�3],5�z�b6l��������h��-￥O�_P��\Xs�;vN� �?��#�4	����X'Rs�>�f��$��b�h!'��?M�f���ќP��oh�' �\ɾ|H��� �7�!W����~����5�X'`i��faj�%a���1m |���;�ҡZ9WM�m3�v�v�t�*Qd0���y�{̆�w�M��	�K?&��D�Y���r6��X9hT4�1ʓA@9���F�t�[�]�^胂�n��\3�	y7n��Zz�n��L�i���Z�6ㄧ<�XBvp�9��I��|�*�w.��X�=�����=!۵"9{t���[��)a��r�,��Q�\��P��ܵ�CѶ��c�q�*n ��i\�.��G}]��q�Ks�A�s�9�Z2�@5C �����zJQ+YN������ �O\ػ���|y�.0\�t��t���y��D��N��*�'��J�&�BZ�(���fr��,�d�9�_�AQ~��:���.Ā����g���-��򄶲F|T�&��l�<V���Y���U��n
�S-/�z��3����%x�V0dC#�S�fx�0_Gи�B��k��t��lF�H�H4A�J[�U���xq��L��.6Or1�Z������5i�E�x>,g0�z4��x�n[@��F�fq:~GeE�û�y��lI���eb��~k������&�����Z�ko�<
�[9R�����^�B��bp�n���x��=�Z>0u�r�fk���1~�qv�l]��������ejM� ��"�j4ԛ�2��+yS �Ī����O�Z�C���5��d�ʨ=)D���18TX��i\yR��(�+2о2����Eۧ�b��x|s��{��4@�"����0�����R]�A��B��P�����K�p��Qdh�g�Z�'��I�+?��Ɔ����m����fi�Lk��6�T �#+�мO�	0�C[r^�eA���)��z-Nf���F��4)e�)Ƹ�e�V{�Y�	 �?�Wt@�JW�&mO��b����r�C�����.k�q�@�^j��Q���y<3,M��/�����o6�v�h䡬ڝC��ŝt�fz{�K%�P'�.�og����S�F�R�(���D�$Òϼ�N.)����W�Y���*�j��0�ʐ�e�0W[M�$��#�i�J���*���'�ǒ�σO8AC�E��	i󞩇��7D5�K*t4Z��n�y��OUi���n~"�Q0�V���Q��qyL!�q=V�z_��R�w�����<�%XR�/AS���%�k羻3l����-F���j���^����po�mn�P;"���R^�`4�*��eިF���w13�DT��^���?-�/w�.�Ap*�B?t�qā���'�'Em�P���3��f+ei����||��֎u/1X/@4��p����&:���Z��l���aȇ�\g�g��k�NUT��l��)!3�0Fw���LZ�X�"�E���59q��>ڋ%��!R?��$s� �|�zB�P= kQ3���IdQEM�9IJ�gb�s�|,@ ��6X�ѿ�����o��^��m��?oP����B�͠Mu�q�:���x,��;�-U��S�ϐX|o��w|�z�{~z�I�{��ܶ��ſt��{&��T@�c��c�{���Vj�faX�g�T`��D�dũe�?��+�F���*��u;�b�v��tu9�[-�gw?���*z