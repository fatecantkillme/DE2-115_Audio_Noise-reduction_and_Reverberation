��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<Ph���כ�Q����Oءp�y��t:N�8��S���Y>�}��x�t��Z}�}{"G
'�HV������ʭ��l�/�Y~j)W��f[E^�נ� pm���N"m�~���3���I�_�v�*"��k�ٗ���������׮�#\�j�&�����=;�([s��-z���^��t�Q�W�w^s%3���_!��fZ�,xl��L���P���h�9�����oS$�P�ݱq�w֟����|s��4H��L�љe�4i[����w��h=���B�u�q�S  ��֘�!�^��LiM��"�$��0d������d�����WP�����?�(��=3'[q{�W�CűOIC�`77kF%���Y07�~�cn�Ұ��r��쎩@f�Gs����\}]��Y���eM�YR���+8|ⰴk�0⍦+�P���
4Y�������:܏!*��C�	9��L��J0q �	_�?'��c(|� 7������`�W��$�1����X��Ֆt ���-Z�q�Y@r�p�_����k�!�`�Ƌm��W�s3�_���V�ue�R���N���В��r��a}���+nw�F
HM	�](*].H���P�:;��K\=�3�N/q��˽sT�a�\/�0�Y7��1j
za�VR�R<�|E����r�qp�:��?� n�ß;�EF0������UcyH�B �\+���@.W�c��P9E<!hkl���71/rG��`fR������$���n`� ���v0;���tN��ޭ�E<���L���`:�����?O@W�-&2:�U�h�j��������t�O�S��� �c�1ք�Se��k�@�u�!L#�-�y��G�>����n���q<;�F��H�9˟e/"Ԁ��`����`[kJg�x;�eɦ6�WX%;��۸ph�ӻ����&u�������Z����'�@��_�-�t˦��^k�:&�J7i��.�ϏAw���}�w�X�'�,o��xb�p�����^�ᨭ�1�g�H��Q�ZW��&v�N�6t�3~��a�&wo�E�>�H�����"�6��1�Ǐ�N����*E�|˽��!4X(�O�����8M��ɕ��H�nȚ2�6���U����A�th���Fc��wj|��*�1ñ��09�G�o�7V��2	�	+ ��x�z<��{
���%�p�ŋ{�Z!XL���լ~��=���=p=��z�ͽ!��3M�up�-&�V4�z��L��B\�����I�q={\�T������L�Dm��U ��?�� ����Nn��z_��1������x�o�)l]@ЦˡW��^�(qp�T��&�n��쪼���Wӿqzأɾd�N#t�|��膝�a<
K��ކ�ܠUq�����.G<������l�ف��Y.�ʶsy�����XL������m0���\4!���;!���E�w�h�zFB�^&"�w�4�:ֺd4���a3���@.�R�����R ��?���A���J�X��J	K���M���Hb���u.�5ʗ�,�Ğ��C�ܑHO��-Z��o���vÏ����1��Mی�`uw�.~�$��
G��F,	��"
+���]p	�}��+�N�}8=C~� s5>Z�;�����U�J�҉��9�Cy����eD�۫�$J���H�9,`��,>H%K�N5yt*0Z�uv>���'K9��$�	�x��B���7��s�=9��H4A�c����\�4�X�$�yK�E�S�(X\]e��L�������ACrXG!6�/�9��H}7w�s�EOd�G��"n��B���a5���T=�Y�V��o(���w��j�+���vH��?�uݬ3��ndF�����O#�P3ɲ�Y�y,F{�(�ѱ����Gy�}��c�J(x!�
Nf!��"�_�@����m�b
_}��u�\I�/�Qgr� �G�4��٤�r�xa��8L� -�S���ڽ�j���
�;�>Đ�rŠ�Z<d/���F4���,����D�h]wL=���]xWN�W*���e*��J�����s@r��Gd�jzqj=���F�.��}�"�즶p����"��3B'������l��B�F0�Xi��,˨����l"S�b��]d��-��R)��C7u��d4 ��?��j@99dU�H�)�?�i�zs��"�-eZ}AI�>�g��֦�2{m#��h<��=k�41Vc���˃o ��z����n[MD�i,1�Wj�������k0�7���3�g��p�I�ŝ0�2�X��ģ�/���%����;��(c�0a3�����H��L@�U��9L�W�<4}�Kْ��Ph���g�RWn��I�v�<��g�p�Bk:���+��E���'����y����u���pG�ھ�Ώ����W�b"��r�M�I��՛���Vw"�W��m8,׺��A����as1~(rG�͇��S�e�����5�i#A��N�d�.�
�?C�X�h���'q��P���5�}��88�G�=�/�oj?��O�q��C����,��cL����(�1WT0��&<����t�4nc;�TϹG� G�s�k{�Sgs�GE��ʏ�BZ U)��#���N���u9�,X� /�	K�h���V�3
 ��X���Ϣ� �=����5�1���(zt�F�� �.y��fE��r��5o����4��h�Vb�l�6�LTw �{�ћį���+[|��z(!�oJ�o z�k��a��2��L�Մ#�kɞ��=Z�L��@�ry0�)�,3��v�ܐ�»Lo��+q�,W����B�q��B5������c�P�F"k���45������*��pU[�M�'sqt�)��cr4Yh��h��[~f9�eJ�����-�{sb������;��긚\��APE�%��a�)��j�F��e��^�nB@�3���sQ��;����2!�H��g� \y��Z�&>Zo;�!��:~%�)����gE���Zh'�W�W4!�8��Щ�W���������&M�q����B��m�El���6�ZV�k�"L�0<: Bf4~�'���8feg�@K�bsc(
R ��)�A3�.��'��U~�����*%�����Rl�ȱ���z��O���=b�ٻD���M�{�y�<%�O+�Ab
�0=��v���5���m"��+2���^�|^'cg��v�%���C������X���hэ�e�4�z?��4�%}�������s"�^�xzL���::_��l�������rz�I+���_L�c8t-���,�*�J�B�ҭ�Y��Z��vh���:���8N���f�"Ѯ�h�Ko5ۅ�Q�?jt��j����9��k�B�t�5|L��֣#��R���hѐо��>f	�S%�^�d�֩�'�q;5� ⮙�����%�/�Y��z�Dm��~��Q:�/B�h�TLOj;���'��O0���/ _������C�Wc���lxN�sba��zYe8�@Vᴯ���{��pr���GIN��&�`�̈́�������� �͏�Q��jM3f?w�RhL���^3��xX1�ϥ�bQ8����iG�8@�zdZvm�#&�J���{��b<��W����	�@�J	'Ʋ�ޫ	R+*���E-i4Z�q�~� q������w�/�9є��L�ںn���	`P}���ٯxW�G�e ��h��{�J���V]�> �T/<���X������Ҝ�k��O�{�t�:�瘸`���A~�G*�B�D�}���ő�E�j(-���gy��i0�[�D�4��_j�Q��7��}��L^��� ^X�i�y����]��l'������!�(�Cf{�J[��S �����uN 2ִ�~��Q�:~\D�����ue7�ϤY�eʃ~�"�2�y���<*�b{����!R�y�*n�r��Ɍ_���ԥ����0iis�I4�-�M�}[�N�|�Q$�k�=��1c���=����iP�2<05�AW��( :��T�Yy��A� ԋ\��x����V�K�n��}7���tMO�����tJ��]�T�w� ]8c�'R��K�=��6\���	QC<ȣ����>j�����A���<��r��gu���8y �t��܏���H*i �S��.�b��By�S7�S�eB�Vy��{�Y�7�h�"F�U`�u%�L�ԉ�6�T��`,\T��N�»��;ya�ag���X�8%T�m.t�8�2��v`B)��6]�n �'k$J��h�ui���zC�E��[΃�	`)KE8\�b5�w�mh~�l���!޳����W��9_��x]���s`c����֒���Veq��<�y��:�y0�Z�r��~���O���B�y�7C�#�.m�o��KQ�h���-����f**|E���K��ʜe3����7�tk���kt��0�ɍU�2�����������"/�Շ�q�C�v�V�8�uA	��qo���v����T��j$�G��$Ò,���D`��,+��`������PX�}�����|q
�k�BG1A�J�����]�-�t��n�.��Y/�*?	���I�Е�A9����L<�(�W�v��cT�����؎�4�?�T��}~?��o��O1���/kpv�Y�e%E9�^T��>���u� ��q����DOuz��$��@�=�Ϝ�Š8��{�+���\�� ���4A��M�s{Ȁ^a���$�x��K�R�Y�.~���<qc�WkA-��=?73G�#p�S������s��᪕�ϳ�?�t���$x=x��Ӿ
�B��N�!��Sh�����L�L�;���h[-+� �˘)�*��`'���u��*�]���^Ή�E[�J�[��Q�*������?�a5|�%�gp3�v�E��� �nYKc=;�;�q�},V=$l�� �tJ��O����a |��֪�സ��>������8�?�U�T������;��P��ۨ�:d��m��;u�F���TX^WV��6���Q��BY����b�8QJsչM��=�A3�\�N��+d9���z56ɰ��]�M��D�����g[S�����$JR.K��;v����(AR�X�z�ع��=��+:����:X�\K���#���)ԍM����l?�|m�C(��j�ʊ����Y��������������`\�D=�pnx��$����yN�� ��<MZ�?PJf�����$�U��qkl�/�G���d
�[�N������o�Vʯ���k�7�?�yc�ҩ +�����mv�I��<��-��'�g�&)��==���s+]~h̒�8�#�����[6��E�c�}}���_g}8�Q@��n����j@��.���+���M�)	/�[�.�@����t����$#�-��_����!�9"���*WH�]�t-2��Y���~��8)��`U�M��$��c�vd@٧�Wj�Fu�E5�͘	��ߒfST��7k癙�f�rQ����ݍ��F����C�^�!�V�͍���ȡ�}��J��ö� 6���������'~@�ˣ���N�l��}��.�۸{�U�PI~�5]}+KI����l	l��/ò���-N8��d�&���b�i�n���V�]5߀p�.�]zn[&ʇ2 30����[�Ė�9����,� �uǓ�E�����/�t~����d÷_4�D��J�W��Vs#J/..��Gv�y��$�`�,=,+�qA�3�!��W�2nxTa0��UK_���⌮x��,ܐ�n�`!���}s��ՋQ�	Ӡd�vg����B�q��d}M������e�:|�|[�����	�n�t��no$��o�Ťc���r��R��>�_*��b���y��lI.����^��i<�h�=��s�/�P@��Oޥz,�9���P	�Y&��)	k�P�q�N��ӽH��u)��'�.p���=A�Ĭ�{Σ/*.���{wg�fۅ"��&�!��0w�n�u,Y�w=����i^�	�cpl̮�| T��_���͆�S}��$����C,�չ��w���#���Q|X%���ҦOl5O�`��*��/o.W!��~.�d�z��Y�4h/�i�G<�Y?J�D�lO�.[��9���x����T�ݣ}R �?e� �R��%e'�~;:|R;�����۽�"�<_�j�٬$P��7�mp��������bD�l�����Ƨ?xϼG]�\;Q�P�qa(�TN��4 ��	V�K����2����9��
ލ���D���L��ui�(��*�6���ѠX_�,?�.�R6!Y�a��O�1{7�����
�T0�7�k�S���Ԝ�$/.��q��xZ�h�$L-�鑁��PȾT�/;Ռnӄ5u�ts�|z��u��	�
:�P�Z�������v�'%�����|���H��sqqӿ��K�L%f��0x�<_�cQd �ŗ��ܷ3���X`)bht��h��Ƭ�q���_\\��TO���qs�=�� ���6̠%$��_��縑�������4q��\�θjsj
c �m�0<8� � �
�q�I�����kX�7�l�Ϫ��;�#��&\	Q\��xJ�<^��|�M}v4�\n�!3�����|�a]:�ء���@p���䵄�\:�Y/+R�^S�"�o�F�x����ͽID����̱f�� J�o5�/?��G�$�t�ѥT<y+J���@$���0����0�r�xX@xmʐZ��h���W�9�g����(�/(�iox�]��1M�3�F�*7PMrư���B8�X�Ӡ�1�DT�[�G	r�����+��2nFs��ip/�� ��_?�ӳb�"���ˉ<3ÙD�:@Wbڂ� i1A�/�!t ���xS���M�G��Tj?���ʟT�T��s�V<Z@�eV��U�S:�KI�Zo�a�7��u_���>�����"׷O`����r� b�*u�?�n%�/�>�M}���no�����Q�.S6#�{fB^"V�m\Gb�46�+�j�(.��������J|���l%y�����Q�zy_��"�~nZ�SnX�t�����Qx5|7"�Ɠ�&����^q��ж9�i�OQ*=��<��3S1����P%��닊:"=u�o�i���b��@�U]$����y$.m��~g�s��>(v~Gj��Z;���?Fw��[c�9W0�#�	���[�c0�Z��)��
�̖y�\d�d���@�)H���.*�����%�8N�nq,x�>���C˽��$L�=(DR��l0) �L�E ��S�"��$����J�L3�:�:g�<a��X�I���
ު6�p���Y0���>����oi��p*�Â��2�[hv�Lm�G�h��et��<�f��f�Ak���@��+lV�K�\;�&��
@�٨�ٚ�ZBU��EH���S�K������/���'Y8����-Ƞ�KJ�D �Υ-Z���1],�x��X�cK��7^��-�cLF{���~�n΅����N 0�n��q��"�x^�3���]�!n�������j��q2�65��f�"�=/i�Y0�!�n/�(�	ʋ��I^hRqIS/hj8���r>)źY{k�J����^�%}�V����{e�"��IW����|)~fqwx���0��9�;&���^h����޲����f�Dt�/Az�����{� v9��� 5��^72�娗�g�@��Usp1o+;�#R�3�_�mQ^��|�2w��°>���7�R�X��2��i��$�<
_8��vzBA�~�a�N����U?B9�����!�kR����HC{'o��b[��^��W@�Ez��:(�}2�+LxG	��C���ֺ�B��t���� �U2���b���J6�y߿t��!�_��*	ܱo�	����+p��T(4os�li�e��Y�
%{<��P _��4	�TtF��`�Y��c1�-O����0�q����CC����5�ڿt�L�@�%�)�Z� sGuJ����t�>9��������g�WY�4�o�&���CĖ�!B��\�2p���x�2�Í��5� w�\պ�);�o�@S�'��(���'MÚ�\`pÏG�
��q�ZYt��}�B蔗�0��B�x��n{�����<bKh���k5_U�X�>��e��������43BO����C��&�
u���Z��,��lt|D�yw��@~��Z�"c�E ��U�H����/��Y�C��uk���O;4*K����c��K�hCDZg��f���\���K�����Z&^#��n�{ך��Y祓�g��C��NѡH����}��H�;��
�0���:�|ӟ���\���v�bu�o�Nt,My�����z����ޅ�Y(�6b����袤�N������^we���Smi�)X~�W�OT�in^�#�؝���nt!�n�����I����{3�i��YR|/|�xJ���qz{��>�3:��Hg��w���+ew��q�<�����kV2+an,<� ^C��i��,4o\�-ܕ[�[�3S]�b�se�2��e�G����>��a6��7`hF�u�Tg��~��0���7M�I� ��by�U��=��EM�^]��侈i��;��m����q����4{��9#`�6�6���Z�#x]�:I�!�Ncl����[�R�$�|J���K˞�Jli�N ��䈖�0)/2����d+nP<��}p�\5J��s�x�̇��M������u�w���3�G(� h�n'�)���y!>	m�hN.�'DG��|�V*98t�QeyY�����2����>S��q �ó��M&͑����,���_��{V�B���H��Ѣ�t,Sre��s%y%�Jdr�)�_ kfe��{x�R�l�Mgn]f*�"�Ӌ[��~G�z��P�,�?M����K+։a_��!餾4D{�z%@`vΑ)��2<�2%�q��p��#��}�lytk~m	�i2�Iwߕ�`�& O���(�̝���ٍP��:�h�7�����~*[x3y���4�J�W��}'��	9�S�& ���kU��O�c8�@T��s��2�nO��H�K������s:o/k�_�|OW�Q�E1Z��#��r^_��Ȏ��!7dgJwa�x����T��6D�)oQ_��84�����Q��T���9&��=�R��R��c�lx��i�ePݻ�x�
�܎F�ub�a9�b��R�.�e���B6kAs*�ڸ�'��6��UrHJ�_���gr����^������e9�Fo�5�J��>,���;����Js>v@���!h:8���q��ŁC������[��,�b4��-�+\�A�ͅ��51�~��C�?�*��`���H 
nBֆ�����`�Ѧ�Ř`��ك�c����Q���
������rX�j���\ٰ���W�&"��D�^A�A�����*"2�₡�E�2'a3���{ݎ�(ӑ��zU���l�+B���jrY;x��K����T���
K����oA�z%yV�D.�5�1;O�QY�=�8K+HB��� 8�pѯ�./uع�_XB�}�NB3�z@���~ޜvp�jF������5�EK��9��4��kd^��.Cc�lG�p�Cz���qt)����w�nW�b`7��̻����|�IF�����_��l��Q�ܹJ|�-�Kz5,<��Ҩ�ه��^�oC�+u�uMGk�(���5(�K�;�2��Lx���o���|Z��hm���ܴi���]�/�t^R���N>p��u13�����!��O>��m3ᾟH���T������=�WΡRf��]�P�@M��}�r+�)�u��,Ww�p:F�mM�%�DuT��}�"
�Wcc�)��7�dp�x�����rd�L��rO�%H�R0Q*sќ�#��K�b@�1�u"A���@��ң��P�9	��R�W���Br�oY���j.�A-P3&g�5Jk�+k	�M>P�YL~Y���M���d1�PE�>����	�TV�a�D5h4Zbd������.���
s.��/��m�0i(�	j���N�Y����&���i�*��-�$�*OD�#V�R`,6�HI$���vbw�)7nc|s��/�?d�b���O�v|�����>c�06�O�6�8���
�՚g�����aZ�	��K\a[�c��8u׭@����oX�W�,�ҿ)/s��N&|��M	6$���=I�6��e�j\��m���3�	_:�\p�i~�&�g���[���p���vj�'ؗ��vꌳ��SkS1�Z= %�;�1s��0�oou��%L����.a2�H�|�&;Ȉ�v"lq��MбC9�
������<HBqXd,'<5$kU��sa����/x�h�F�a�ft8��]�`�}��*Q��?��m�2�	��ʭ�VCF�m �Z0�+����O/2>X�&�����j�Af�I���7��̚w��;@���P�����dSc���=L�$"�����ōT6Ĝ���нɶ�����ۦ�%z瀳�XQ�J�]������$���M�K�����T�I������O�������Y�#��"%�6_� ��D��1V"�~#�����Ш����(�P� w��M'9��ML��0��ax�³K�����`5S�ݞƤ��įi?EӅ���T��-	;���|�1V�m"� �>y.0�3�h$�}%���K���K]���u���a�M��x9����(���5�����C �����5��.@T�j	��x͏� �v����P�@���|���	�����k���*U� �)�r���hVȆ<��M-4���{M˘^�zmڱX�f^��i�0)�/Ak�<C,@!�������v��ž���'�� ���PO���,�4]���9w��X���9��dATA��;�q�����k������@�3{k�c-΂���|ا=c}��Wmf��ˆ:�S��s��o�A��S�xω�Y #&t�9�-�RJo����\�&:���E_*�2��Nl�^
ǡֵM^b�tmc(�����/�M�{e��
�ض:���������6��oM�Jt���A�:n�"p��CR+��e�:���0��4�!ٔ��"$.�z�W�O����R^,eO�M��J��Z��Ŏ"kM�k9�*j�'>��ز6���T�$�0�ޟ��F~��p��6q����L��ף?,���I�_E6˦A0Ϟ��ƈbDR��A8ꔒ���3ƪc4�U�fh=뛟��G,<־j�����PWYLr}��{���)	����)ɛ|�2�%\�J}G	���wCXLJ�k�"ֲ��!�R�*G���A-�&Lh|!�=�B�v�1gW�E�B��^@��8��{!��(��Wш���2���H!����`��փY�<���\�JY\ʤ)o�Ǵk�������Tx��E��)X �dB7:��}�V��xF��A�MHqI [ʟ�����(4�EҚ�ѯ�[H�*��-�;�����]��=Ǭ���r�����W���B�D���m�TX�E�w��Ʋ�}����3��	��E%k��w��U=-��FG�*A#�yS�����,��Y^�ʇj�Ӯ�
n�ri_@��MS�wfzZ��!I��I�	�|��������}WY�d�z>�Iqxxx.�.WyϢd~�
�r�lF��{�YH��V��E�Ԭ%�����-�aO��D��aT����+�ϸ*/����[�M���-�Gr����T�p���{�́���2�t\/�������6�-��g��⑚o5�2�:��P{)�o�Fr�A�<��,��{$��p��L醢$���G���x�>�U��B �[%QN�BW�� e��S���{eu}^�*J�<u���-�:j�C��R����t��j��	�~q6?�!   �V�'P����ի�y�Ut��P�`�(�K���@������&f��>��\��̢�9�]���)M#�a�k��{�%�e-V�7��!O��LQ�rI�	3�,���^�?��Q}��MA�&����Fuz�� ��X�6S����*��Tfj��ϒ1�(Y
����ܛO�`	��F�a2�):/^;�Z���hq�`u��#�� mFB,GQ��&�j��W6������ �S\XN~��H��3M�T�Y[ʎmC��cߡ���:���Nn8��]�Y����6q������ֱ�:û���c�K.��w�f0�G�um����l�s��oT�� �U�0Q�$m�P`�µߕ5����9u߹�h��R�Eu�'�8麙�T�];*���$X.�j��4>�z:�x����;�U�!g���.��zFJ�u��k�2��~�*]��SXx
�x���0��o�<`��u���B�xT�-�#}��ߩRcg�u����M��(�@+�y��4�Y2�,�u]�r�t���+ �gZ�V�=���|&S1m�B�6�'dCC�N��M�5�J�ֽW"�-$���Uc��(��n�{���P�2��_^�vm�qS�KY��"m�;��}� sk�٫�?EsrIx{��i:�ycï��*��,$����w ���e��OM^p�P��YZ
iPt������A����h�-��U���8�h�u�-"�{��x�+��B+�L;�𴊃���yv�z���`��q.wq��U��<9�}��5s���>��'~3�e�k�U);T�a}�`��C�B�]�T���,��H�ql�x[�ll���3�u}�ő,���fUuZiA�XcA$��1]��TI��@��,�]�z�'�N(��J�/(��)� Ê�y,8��i�BZ��(�Ș�e�'��y˴��I���v���zZ6�mw��q�ŵ�AT8�v�� �j H�P�39Љz^P]�23jB���'�k�e���.���|���͗�A��{j�t?c7�I���F�l�"Q(;$����z������H��OA`έ����˥�7{E_�t9O�LI���Ám�����?!aSʰ�!�Eoc��֡�U��y^�X��!XR�t��o0)"�!�w!HGؾ�Nս��rB�Ⱦ�x�ƽ��"d���"�3Ќ�#�c>63"�]:3=j�8��gN�R�+MR� �0}���%A���[dg�K~��䮧\��}8g/}H8i�����P}?��36�} j�_M�>�'�~$J�ߖ��n�=��F^�Zr�׳���\yff��=����	�!���.Q�V�K��R吾�6���/���PW `���2b&�⪯��塄f���8�Ѽ8d�G9`��s~ш��4�A ��HG,�FQ�9��H��є���s�����_��㬂ovH���ʶ#|3C�0c���Nû�r�)�~�N 䙎-a�s3����s[B���N�u?�f�H�\>M�a���3EՒ��m���%�M�7��8^g�U�"Xm��1-�t����ҝ�2W�,��+T`?��-{�E�=�V�]E��JU3�-h���%Σ�c���L���#���5�'7 p��9VQ>� v(�⁗��GY7�kr�����+��(����
6R��{���J$����A��S ;�Q"o�6��/p0�Jm��� ;y�K
;�v�!�B�̯:�Q��~&�R��]�>�!���ɧ�ͤ�����/�#w�*��3�JSiE��-��T>G�@[�6�;�����?�d���X<�6�GU	��tw*x�/$�m�{�XC��l����7�tf�X�������E���q|�Ǖ��E_){�c6
�c��I�`�.jRXfl��A @�����u;�/ad��	!ك�>���� �|�s�_E��﵂:p`���W��z�0��:T��M�8�>�\#��Ih�6h���	�9�[��n�.\�9�DsY�h����Cn��S_���(��\�<0��L���V���'��x]�.ɄG�A��֑�{��/��ٻ�|���ٛ�M��Lh�����qx;���V��g��B�L`����Y�@;���)[�K՝+/������Ȳ�+�����)�y�'��gE-򚌨g�5+��KǜH���{�V�v	E[9�^��=�TԠe�'4b��{&�*Z��k�=H���m��,@�9f��qM��`�S�����Ř��[k���d��E���hg�P���g�n(5��t��ݺ;����ND���ꁡ�(��-���#�l����pD���2wZH�I�Ӡ\{a H�]L���ޯ�k�z�)Ywr�c�2��y�4��q�ܑ���T<;���H��4�+�S� ��z��y�F-1��s��q��}r  H1�{-�IdJ5�LWiU��ʰ6!��������fo���+�=���fr�d��������:���}�8�	X��k�_��i�|u�g4��VDEK�h�|q]���Gt��n�Zu�EZd"�'3ї�%<Ǯ��r>������E��$5S�l��4]��$5��A�����e���K�0���^�X�hjt[G%B���F�o���!��\�Vl��S�o���)�X+�dz\��<�T$��, ��D�{շ��i��&�3j�FF����G�Ӈ���<C��9Ծ���QZ�+�e�Z��<:+�!/lnc�y#f5�ͬ����*�cn�]6��Ik�M4���sֵa�ן���Ů�p熞��R��az�����mB���k��Q�����	�n�К�N�7��McXR`G���>���S�O��'�R��>#�7�˦�r��N����*29{,�.�}���'\�Rrix����P[A���1�O[�g�ۇ�p&p#���_0Dui#�NM��V�"%\�8�$`aj:@�����"x!�\Vt�5�����LiG��0�=��?A:K�i(:��y�۠^M�}P=Y�`��Q3,�AV�<`�f�Q`�'���a<�fG�.���u�∆j��|q4��Q�����nӄl��r9g<�������ʦJ�(�ZZq��7.k��������%�`	E�*�m���i<�r��g�y���Q��i��\��0 K��/L�����y���R�L&�]���k	��?#^�����P�CJ�~�:R�-�.7SF�W<A|'P-k2��hy-Y�3�����/��z}5��0�$=cOn�Yh� �TDs.�ͮ(�
{W/�$Gv��3�Р�5`�XtA?�'�*	"�v��8���;�`�q��e�n���o�X>G����@�Y�@Z���9�*Ԁ?�L׏}���,Ų��늮*�U�/yeh����)��Ō(��:�K^��v���9��2���?���p��	^V�s9.�X�9g[[�v%���`27��f���m���.�1g)!��
�z^@Vy>�������0�%�1�pH�z����0*S�ƭ�nIZF�	�!�
�Yk��O��f�r���u�� x6�8�NW������q�s\sjl|�����rw����>ʙ�S�<,[����@}��8a�C砟��墁��IT� v�tTɴ����P�	O�\�ߒ'��O���&��Ĕ�B�����
S����_�[������k�Ja$)]�m9 Z�k����EGa����ga*ܦ�l,W5fE�	6��J��,��߄>�V!zm����ǀ�ZJ�f���Uf0�#���Ԗ�+���u�"�(���u��}NEY[�tI�x�[����[��]�#dsQb���%vQ���8w�r �}x��f��qW~{���Q*��7֜T�7j�� ���
�&ج��������M���$o����Eڲ��|N?5����]:S�D�ǃ}����߂����5N�c�.����v:Rc�=����ܤ�h6�cKP)��
o�$!sMW��Jc�}hAf���YҢMxO�����]���>U9>�8���m-��ɋ27���7�M(��$jW�g�ؓp
���Km���w%�z!Tt�U�ާw��q,��鼫I3��T�-E���Ø8�b卐��^ 0�N��ª���B��8�ʮ*j�~���^������jz��{Q~��b�cL�� ��w�e�Tp�T�9�Ai�&J��]��8vH�ۨo��Y["t��y���P���ͥ�у��	���wPM������JZ[r�@'�u���5��LC����񐴳��K�n��4����|;ph
&�6�ql}�@Y��`y"-�k�����h��c8t�rb~b�j�+��h���=���
+�$U����fM9 bv�+��L�����oW/��þ�'�� ͥ(��v����@I��T&�Z����/1J�X���J����#y����L�Z�,�Q���1�[*�Ͽ��&f�8Λ\<�`O?xІ��60�A	"�P8��B���7��Ŧ����Wu�ƕ���X� �cT[B�+�N�ߵW�uϳ�;�20t|`K)�%�'���8l�+�?�w�O��l��,���>�W�ʷ�L�	���M7"�7�ჴ�����!�{�T���E�+#�)��5z(�L�*)�.]�sK�qԳ���M�|��̫p�0��ۨ����6&��|W�)G���6/��������ʰ�/OP�#��7,0�޴?�˥���C�����G��oXi���u�!=�>��L�p�o�}��|$��>�#ߓ���w���� MKW�>��):��U0߁u�.�_x��>�Ѧ��H�He4�����\��_��Q����/��������)l�Gw�>�7�� �<���-c�����
բ�����v+�p:ǩ3�5Uع� ����״b��o��@����6����}��j!�"����3�l�n�Cz��r����jMp�Mt�{A�����
C�� d�#��3��@��il���SA��%�z����NE"��I�������cQ�|/{t2����6'Z-O�<o��G܏,��PS������ �X�H�T�褢�1?m�����_�'�h{N\w���u�g�;+Q�8y��ƶ��H�[�"�����T�"�,����m�+x������(�����IZ����f0�<�ɴ�q��ę�W�e�y�Xu�h�DhZ?F)����8誂��2.��X�s���Q͟�����DJY;=�7���q����É5KP��C�SF�?̭���������!q�(,]��d��(9�F�����)����E��z]H��tO���.���EjE�lem]���\۽,��!a�	K�OzҭO��e �@B��h�ad_�%_z��ⅶ��:d1B�z��&�55{OE��K�|i�?�?�t,*����6^t2)���M_88A�	rd�^��b�I浏��� �O�&H�p�N�!��%�oƆ��=s{�醷�-���8_3ғ��Y!~TY.-�w\�r(|\���cPV�!�䌜&q��;�Uu�Q�/�8b��͎F���(�T�n(�fS�]�`����ZKa��&�w�nŶ��P�?��W��~G�ލk�����ֈ�\(��2��S��^�+�o� 6�dc��Z�x�O0�Tb��QLD��:+GJ�Z�,*A+l�>�3���;Q�������O19�%{��vt���K���u�[A$&=�4E�R�L��ޥ]0�;�L�3}���!��Y��x�8��F~{`��m��OX:)�X��G�/nl�X�D���/(��-����K��ߧOd?�{w��T���+��?k+t�������&��ux)#�x��rg�0#����(u1�U1�$����$�����L��[2��^��)4��rR���������B#:ɻ%��]���]����F_���_+�<�_�^�B,����]�^oC��������K�P��T�
ˇ��"����3{�D����wb�f��G���J��Ac=���X��# ��ɷe����1�$	~��jN�������V���x`�"]K;խ����l��d"�ε�{>'�v�i��L��r�%�u�[ޙ=�$�F!9u_^):4`���>�_�pd���Rs��á]���!�2���6��|%/��sY@T��0�6�id�E���f��w��{^J{�}.�D�쏳Ҋ@��6 ���~���R���D�}��{R�~�k����I@�P��ڒr
�~�����Z�~������ClSR5�g��d:Ih��O �XR=W�eAO�C�#����xH��1�����ͳv5��*��&	` �]C��x]8?%W�7���ӄ6���GaF<x	3�S�&� ���Q���ܱM.�3z����_C&��:����������0!(-��SP�����|��;w�}��H0Q,yn/��W`'>��ɯ�h~��W���
�B����1���*�?�a��ttBv�eST��SL=�V ���j�;P�Q����?~"�O��������?&A��Ǒu+s.�9����bթ��3Qd���$ɷ�i��|�d�X��������:��
����GTn]$���Ny�\;�h�M�Α����`�?)�r��Z�l�T���}W��AYӾ'É��_ g��9�z�,���tYA�ņ�`>n{8L�k���D��%%l�y���8�W�����
����r�M��M���`FJ�S$H�K�Gs" ��ߒK�a���"-�6T
�!�糔���.aQ���bz�ߌL��#�s�G (6�����켴w��s���Z���ǜ(|���U1iV7��`Z7�^�Gǹ*@�gE:8���xwيf� �P$�~�}����]���pL�\���c�RC"�ǅ*�H��r�9ke��Eb�p�a�P���^��ݣg�Jg�ʨ���%��@ѰmZݹ�V��<��7� ��1�h뱧}xY�=?R�����E��}j-�U�Ď	\�%.<�V0c��D��m���2�$�?��	��)�=��[����
�n�yIi�,�f�s�pV{\��,49ߛ>�-y��ū��?�Q�$���A6��94bM���S6R�$����.T�x|n��W��x�ĥ��
�>���k�(�3xK����V�k���`�S���V�133���G�W�v��b��l�h�;%@����˺M�C�a�e[a.�-Z�ӏ����e���T)��4!S㍋��E�K8b����3�BJ�������4_@'���7W�|�e��ʧL��"e��.�e{!J���f�7�yf��i$o�66:.���\�Z�A��@�&a4��g�����zǉ�	���P�#�h/lfC�|���/���<�?��S��N:Y�C��9Sũ�@��W�]��98�o���f3���@G��^�#��}*�
��Z!6�KQu�\ܸ]��M��Ɛ��F,�/=�!P6V�b;�-]����-
�3L�X�P�X��9mW"�c�k�����"harb��/a�/�����6:�%��&3"�K���)�T0^`��Q�d�C&����T��z~��&^����l����z����MzPbq69RƱv*Xg�`�24P��ÖN������n���A���|�Úsu߹<ɴ+0{g{B�F��[�B(,�79v�q�ʬ��4��-��ƦH�>p9G��
 �P�OP';�QuJ����Ð_{y�$C�ƂU��0�-�na��P�#)M�0�<c�Xm�j?�F�[�ZG1<�����}E�^�1����YyJ����\ˡ��=��ch%���SK3X���z�O�����31}��%`.rO�vh�&�zKC����%!Q�pk��[5J���Se�.j���qRh�L W��J� peTw��������u[�<ԛb9lQ�^��7%N��ӏ67�~�~��ŦX�zJC�Rc�/C�Ǿo޿�0����vx���}�1={@�8���S<�CKꇂ���!(n<�Q�\�����7ө����^cr0ME?��a͌XTAw�Ce��Һ��7ȋ0+**�Of��:2�X(�E9��ug�����)M]�}��7���("�U2F��r��*rԴ�M/���e !�nV��4���>;&=ɨ�4�2���e�w���q��web*ζ��¢�n3�Ѽ�ӵ���8O}�v�u��^��o޳aj?��'��)	Y��7K�����%��?���v��A�<�l������f��k��7?�~���Sep#��x�٪�K!h+���"�z�E��C�f�'NI�sDy
�T3-�MO<���+������-T{Sʁ9)��Y$ 4��,$3��%����r/�l�k��u���.DM��42�B47鼭"L�I�2�d����T�D��\v/���IZ��67�i�v�.�B㕮��^��7����%��y�Kp9��Q5Y6���&��]]�U�s�)��#��%K���7XZ^��f�<2�"Q�+���\gV�f��$�a��3ck<(�@z힮�.��� 
���h�+5��e� �����DX��۷~\����x.B�OA�	j�3������<t���+�:��&�X/��!fHv����_�hw|����~��Z���,[;�P��*�J^=ǢN6���N#f_)b����a���g�6��~�ے�+�D6�ޥ����X]|a�֣*-e�{��Ʌ�9���&�"�xp����7}��%�k�9>*��1��wEU�*����WfY=))�e��āS�vVH����Uԓ$��ֆ�������]V�8݁� ��&��=l8#3�2C����̿؊�}�E�`��M�7������o%�]��L1�q����`�2k}�˝�u��5�"ݠ|fV�r-���9 ��ٽ��Z��Uq������w�.TX���}*]�3�?�-glQ�J�E�T약�?<皹�Zt���Z�ъ��rr���I�A4��qy�D���l���:v-����3$C�����2�k�r� �`���PA%>�o�tS�N��l�P��E#��g���Z�}.3�j���NW���a�G,�x�G��Y�����$+���5�����o���/
�s��/$��,�vh~|��3ޔ&�Ҩ(+���r*���1
./�K���g�cQC���Rq)�N�98���F�Bj�P�\�Z�z߻k;���$���߽.�
�",W5Ig��pX������$v�%ۿ��tK��+׳����K�a�i7��M$nV�p�[�s���)�����;C��ߗ�}�Yq�d��9�4i'�f�%�(JL��)���P۔�,.nW�J�!���v�"Գ������:��,1>�&�.���zXQ��e�w���0o�D�f.b{P�$h�>	��q<eM��	�<܈��#�fw���H�84��L�?���k ^����D�t�&w��
f2����S�raǄ)ȟɇ��QE)"�p)w&�do��'����R��5<&{�b�m ��J����C�a	�m^�A��˯
�G[M�Bj������U�g����pl���+�C���/"��)zd)H����^J���'���[�Mk%�Vζy��}���UA[��,i���+�ɭ��(䜅. �H�h^r#�oMU=wqjl��h)Hǲ%�̆����q��5��ĺ���-�N�
Z���w�%u6�n����z�8B�<u��3]`����N�5����2�Ϝ�Z�x O����`s�2��m�BԖ����@jh����:{��B�VE��k���ͅ�cރb;��h��>��Ң̬��Pphf��cxGbv�������6q���u�-���)�^;�@�ׇA{S��Kva.������8��m��U��Z-�ț��a�i�����x���p���="�jB��k��N�w�m2K�]i��d�i��[�U��F[�K�H}��)�|��,p~\��@�k9,^Bϩ��̈́
�����Q��[��k����S�v�Z#NF�v����,X���R�%�ɣx���>;�ۮ!Y���Ob翟�f0KzM�`�șSg���7&t�hhN?���KK/}�p#	Z/HL`�W4��`7�b�}V��sC([Ǐ�p&aH���-�d~V5&��<����W�tp�>���ߨ��Y�B~^_'��M�%-d�X�l8�i�bˢ��R]�T�zFmk:����,[����:Du�[F�N��j�AZ��9��7^Qt�g��v��uw�@���~�8DmB� ���.)kG#x�R���J����Ch����m�=�5і-���uH>�}��Q
�-c�tJ5�_C=�ļ;�:�rHI���Cׂ#�u��>����fN��p�5���;��������g}vM���*�k����n��̩�"&�}�kL�'�1�<Q�;��3�rt}}�_�whXc��j?*G��ڢ������)&����Q�҇eA/g��W�֖�t�.y�lq��y���m$�����{ ��]�ƀ..hc�Fѻ���2[��!؉h�X��i�ȥ�����;��j�%ڣ����VH�ޟ�W)�-��b'f>�F�5�@�m��Y!��N-I�Y:�Szb�q�k�T��IՏk����j���	K�K:����Tv}���v"����ư?��ܷ i���I��T�N?��1��v��R�R3ΗZ��¿�C�z��� ���<pވ�b�ú�9�k=�>nьS� v6W�]������[����=�ɐ�[�����2����;󿎎:�^9�����R�z�%aY��[N�E�Ԁ�I��l�[>.�3��]��ڨ�@�,�p�o�2�a�~߃�+R�JAw�z��&����Gj���l$��E��@�bg�*��GZ94�}��T$|�����	����_�bBV��L�;�}��(����|9_4�)E�	\���đ��E9O��B�z��p����l7
Ol��g׆� 
��, �0��v�i�C�*�?�W�>����6<�����������-w�N(*�ȼ���`� T�ۏW�x�5�6�r�R�]y]��b�.0�=�*�m�E�BV.�Tr48
3zMM��_Y@��'������I�Zup�@�*ձ�Y�j������?N����b�a��>�3�8.u T��zěј������fi��:gP�Hm�{���i��h�4�m������R@jM��+�>Ѣ麯���G)����;�%��",R���m���+���{o&Uꡫ���[�2!�=r!��{���H6{��?<��&���)�jI[;������_�y&P�� �||#��
��2�����<y�+��	��P
kX��#�,�@`��!"� ���[_K� i����B/6���l�A�Z��޾.�Ϸ���|��g'�λvQ�FrY�=4��W�g�$#8��0�)�����(x	q&c�c���Fn�n@h�|j����P��"^/=QZw���	a/�I��������a��X����LI�v�bSA��U@�����-�,�q���u3/�v��Ҍ|�OB��I_&'���UoU'lL�r����Z�bV�*��{LK��?b��X-;?�T�a_�g���v.O�����9C:�
��o���h�/��4x������oش�?��{aAG]٪4 sJ�w�mqJVak)|�߄��}9 ��
@5O[ⓝ��g�������dԝ���h�V�
�Hw|�/�+�C�X�����'��Th`��h�*��B|ti���Z�hL?v�B���!h�L��\�5�!k�ך|�JɨTލ�d��[���SEC8$9C��-�X��p	�S��E�=o�mt�O��f.�ǉ}^t��@��T3Gz$�ɷ�G��>�������9$;
��ݑ�M%�0l��R~[�B`z7����ʣ���fA�{���nG��o���Z]��d����vZ��#=�?�����裇1�\k� `Z]W���b�� c��j��UڡD���<�&3E� Ȿ*t�2��v�goȋ���&�i����*�/�G��PI�����lPs ���r�d�d߽���T̹�T��§�7\5TyPC�yf��OE����}��2�a��)�W��fAj��bT6�,�H�a����X��q\w����I�p�����0Ɏ��se;�ۜ8�4/sq�i�������E崼�C���Ӧ9e/�������ߏj$\���g�?�>�#7��P�7'J�y���n�$�\��	4�<��z�M�WZ�=w�Ɋ�!폣q��2�b�}���V��rF2��Q=��D\�d�����%Tr�*_;����IP���02���d��Z����Ҽf��D
{,/{*�,�>�sx��rMiZ�+;>�L.PA2��̞�6�Ncq)��OF��������:��B��r�,�}�Z��cD�F\j�9�e�5x�����/�f�MQ��q�Fy��?h����H��q	�wTR����l��P-�Ǻ�o��=�mՋ�+s�\�sD�Κz'�	�q,�Y��� ��!�PGc��ݩ�΂r���Դ��+t;a�$%�dv7S�f��zP�]s����}���h?�Oc��hr`�zA��Q�Y��{�R��s��RsuA�(�1�Z��ǮY���D\լ|%"��$�-i�T�J�	�+�jB�⌆h��]D�U��� �6���E��qm&M�$�Ԍ�hܧ@;jf�(���|z��(�=�2*�O���C[�l��?#"fF�f$ꥷ�W��of���hf!}j$�$Y\6�.�����y��I^����;�^ã^���1������`:�j�e���/�k�WO���4�"U�\�Q�߱�þ��-���n�-G"�$V=S�)f6m��7[v�}��Mᕐ�dB�.�����T�rQ�+=.��iP�#�7ޝ���K�������]g��챷R"Tb�SH�x�ᒨ7Pm̯J�5D�]�kr�~ԃ�Ï�R=?��Q1}OX\;���E	T�ķ��#ٮ��ڼR�|�:�/�A*����ԙ��bT����(;�����0_��9r�tT���$�9]�n��2��bhGT}c�D�B2Xs�2vkH-�1n�"@_����=$q���,K�����g�3$j�;q��Q�/SV;�6'��qS�wE�5���;qC�T_0^���Ҋs�"����e����R3��j{OF�M�Ny����@��R��x��Nfӧ�����ת�6��\C)�P�y@<M��3�,"學2���=��zյ7�yd��S�L<�_��j���:��o�-����c�Y���=�6�%t0_���@8e�A�B��m�ߨ�]����,�q�h�@�����o�N�2��;��)��J������h��D��·�"�{�[�4���O.;.�,~|Z�d
iD	(�ܛ�({���~bT�5K��%���./C/��*��;��i(��r�(�(�JM<��s�i��͡�k��5Y���5�ԻI�BY�-���M�Q���HZ��ww��\q>:)��1�_;�K��5����ς��,H�����)�SP� �A�-c��w�-�z���i�;ߓ���D�"tC�L��9�3�e8��ֆ�-��{/�'��j\(�'�o��?u0f�r�nv ���ZX��~I��Ї�7�����R����4�n��c���@�����ө�Xⴧ -�ѩ�j�\b!�ܛK"�����#�mz�&fW)��pl��:=c�/�^�h�L9�D��1�E4��>���O���lϺ�(_�v쌚
K�e��f��ŕ�߃w5G�=QRA;�l��������\M|8%�H�Z�����P#֭��"*�K��pp���``Ghz^�H��Aj���B���&�d��%�Nrh�2�U�R���%�s�_= �˜�-���
����~C�|��	�OUg;k�k}3��}<���"�+�r��bH6��	��%�$p@~R+� 3���Ô�� ߲�&/w'������C����97-|�v��?`��@� 1UN��	c{� �_M[�o�f����KjRg���E�?/�P��b>���fM��ܭ���x�[ڃ
��I����ш�(6��s�W��<��1r�N-#V�y�=�"�_*�����Bl��ԑTF����;dx�ߛr@G��癲��CH�?���;i)mE�)�1��W#�Cd��^�}�㦖�,Z�Q�ܘu���V�v]�Q�Ʒ���=����bK���mp���Ǫ`�Rbi�x(�|y�:y"٨ag���]+����r^4�6ʫ�"@��m��f3�g��Ak�]�n#6g΂���MS�9���@��a-s('`�@�X�r]Ǎ�������?.��X���As�^%����O��2;��Z�le,�*Ë����MV���k���Y�nhe߽�y{�)��I�h�_v
���C쥯*����6\Ra��Xٻ�M���s)�$xPփ�&��������{JR�e-h�@W\��H:�:V��]dyS�Y#�߿�YQ&SeVo�K�dk�URJ�p��8�e'��no�����3vM����Q.J���e1���b�x a�v��C����m!Ǣ�Z��[��-�I���'���^���wq+�V��:L�c'qn``���漝�; �D������|a�8Ɓ�����_k��o�ԁ�@�������+]ܕ�Ma<#T��+I��D�i(v�b����U}B��^��~4=���og�!T�K�/0f�`��|Ӱ��WY��4�����[�	�N(���?�H y�1��ɳq2��h��UA��m,`o����mƺb���q����S�d��rt(��7���Ƙ~[^��D'��n'ig��i�sZ�k����bA�e9��`7�Tͽ�_�����[��0�L 6��Ǻy~���MZ>�O��#g`�#��%&n�,.�5��g�Q���rk-iiZ�Z����*� 5���~�6/c>.��&o���&T�S�=�CA���В�XUDD�1�I-|H+F�gJ��gh�g�ۅ�:����m��Ŷ��[@#�Jn�-w���N�y�����E�C�u�B�|1z��u�?�KC.�D��g�s��bn���JG}�rM���c=��[}��_f��~�4 Zf掺-���\k:8�� 3|�$��ӹ��U��O����aj��aΫ)����C�/�C�yfUfn{���N�"L!G�Gce�4\�q��وjCc��MН/�C�i�����|/����Pl_#�t	�h'6�{��V�ݬ�3����Oz��V� mB\[n��x3B�I	�̉�D�f5d@�y1��O��#��ҍq��������94�x!�B8d"�
@e|�(��3˷:F���?�d_1��;�N���˫�͠�RZ$�-Ab��� ���R?��[y�M')^�8A�g���#����j�"�,����zz	��
͚^b�V���߉D������K�D�p��M�k�!H?A?����1��8��:Ѡ[����q�"�K������Q7V�y��/wgL;����>7s,�Dg��nlf�%�l���M�m���ǒ	�t�N���v�з��v4�Y���I��?�[��(/����N�b��G�72�h�ls��	���ެF��CKtS��"�`�$0�AT�6��؆2r��>��d3��+d=U��eOO�'�*0��U�C����;D@�xH��W�q8�� ƭh�f[x���V���%��~h���P��zZr˨����f)f#�k�������#�����.V�Z	�F{=�!����M����ۅ��軩��ڢ��:
�Ց�
0u�@���2�]��k��q�cM٘��A��4��,i0cZ��`LZ	Ē�u�̮3�g���;V�]���k���,�,�L�����x.2�I��h^�Q�� �Zr�Y��-�����ZB������hm-���R���сn8L��J=�.+�s�x��.`��h�� ���gJ�e��1���8�<�tvUU�u�)?�f��#XZ�e�F��Q��S�+گ�
(�@�N�ޝ��`7�9�Lj��k]_	Z�D�H7s����hK��c}�	����}k�X�4����Rab��՚������C�B��4J9���vE�
�s"x�cs͊��qv@-���;�u�ֈ#����*"�l�Bу�9�M�j�×U�`��ͧj����������K�BP��f�Nks,��XYC� ��g�-D��q^}�{Zx<Gs�'F�Cu��}*��Ѭ�Y���?%����OOv��V�KT�A�Y�3NUF�2��	�%�����g���-L�'��3�����	�����}��@/ՑF`�\Y"\c�,-��]��:�x���:�'��N����� .&n�:���P�i��t�=[�[���׾�^K�[��p;�2kdrX�P�Z�ҙU����9b]�6I�#7��������X������9C��4�����o���qR:�0ZxCH7�-Vc��>M��6���6��"�f�~�$��
\{�N��?��b7����"m�xsI�������t,����4;�g������WhDsI:���.ۨg�a%���׮x��'�Oݎ'�swTb�;�~��t~Ê����A��88�4��&���ܰ��{��J���ԍ���\��B��{10#������a�^P�h������O�0G��	��j�^��k8�/搼�e���(�*�������EX��|��mT[(b/�?���b��(] �6{�܋�ʾ�S/�O�]�g�Z�x���C-~`j ��B��!�퐠,�.߆�P1�PY��m��ZJ���m2a�R��;���j�|�Wݗ��L���(Dn�;×�V��j�Bn���,y�-��K�P�[@�{�f/� z�}�n�rn/8��;a^��;c�Є��Un����E�d���Hv�:@0@�mgL��~Z��0\���tѥ���[1���Jи�C�-0�u��"7{g���캄؃�[]y�jg"�`��~h	Zup6�Q<�| ZV�Y���Y��%1C=���3ɂ�w��AA"�)�3�@�],�=D���u�]������VR�[��r�~�չ���8b�	��G��cPZ/�-����������`�l��z�+�a/X�U�G9#x�������3R��w�(�Mj��0I�yU"�_��4um0���8�E��2���Y�p�[z~<�!~k����%C�Y��g�r�N}L��,��D��^�n� ��/ύgz�;���^��e��Ym�8���*��/����a׬-�,R/��C���f69A�����JI��a+�Z3�Y?�S����u�(&`.�� ��+4J������2˱v�!������C!�\�ʥR��x���̆�V�w���ڪuv�o�_��w_�(��6S��CL}v�Kɼ����f��[����}�Lq�q�ݕ7B����=_�\y�Iah�P_ET#b>�]\����u* TZ�N�P�*n��#����,�JTܮ�_�Q����,t�w�'O|�L��u�n��dW�O�j�����r֫UCQ9���M!��3u>i�ʝ]��E��SS1N�{����_��.�4�?V����i{Rq��g���^ʟ���e�I�/T5֤<�ŷN��#X<۩A�ߺ6YH�A/]0�KzU
R��⾹Ec�~g���~8��VI�]Z�B��Ґ�EŞE+�q�
��%��M��Z���@�g��S�O�n���C�2����s���	����-��jAύΤ��!(D�w
�g!L<��r��G���n�k���(�Oi�I��V���+@I���YQ�Oa=dvo`/Z�`n�l����{X�5ܣ�tvG�1���Bt[��כ^U��V�)0uat�A�F�vt]2���X��c�-�s�Ċ\�#��B \�~ �k߳����W���!"*��~&z$[���`��G�`Owgn�]S@�C�3��8R�(t`'X�|�±|4�ฯ�� Q�1�xL��� ���J���dY̊��Γ^ŏ���4y�A怺$��[��B,Z6[Y�S��M�̵��-T�o!2�h�>t��1�{�����p=T�>��.PUpP�W�)v�"w�B�H;�	fs�Q ���ݿ�?�|T��\�8C��y9�{'��а����5�$�~\��S}_*�lU��c���*�pK�����1�O%�يt�|9н�Rc_%�;�� �����{���W��Mx40�� ��6����;��]T̀��+��%�9걔�C*艄Gf\��eN��tO�O�%]v�EL��w��"cVT?n��ܤ�j�qV+M���:F�Uf���ƆI[�#�l.ZꜲf1����pmǺtR|��ˋ���?^��8����H�Ap�Vw;�\�&d�f@@��p��AL� )u
�[#d��-�7|n���ؓc��7ڒX��B�<V߫N�ݹ}����:����	I��l�9aH:��;�q�"\7$G�!d~����+�#�F���4�*�~:��K�m3�L�|/=���P�K��Oi{Q��H_�\��o�[=��� ?��h�S��&���:����\������K�ٷ8>�7�E��?���$�P����,"�1]Vp,;Ho-W��~N8�3Ӈ~zV��$R��
���Ь�e�C�H%����=�8����w>u�ȓx��}�]3�pn��ul���:Ȫ�]V�*�-��ec����YTci��Y�-��w����_ة�6��.BR"+�J��%BG~p��δQTRW\:#��nPIA��(�֙��V���&�
�1�ms׮���zû{��)�`d�A������*/&?�ٗn����BY���x��K�)�`�_�è�k�Z�×�a6�f�2-��`#���*X�'�vU{��g�^���	�㝞���b��s��M�'��_�&z����b=���x��t_F�Ց�.ASH���y΄�x|���_L&2�B�1�Uƨ�i�aUI�������d�ޜ~��Ow���+a4@���EZ�lԁ�%+8�d|��\���S�p�V�'�I��^!/�G�U����[y�:5�2]�K�$�v��A]����W��a���I~Yʨ��YԀ�Q.&N���A9u���G��*7?��7�g�E����Zz�/�B�s�U�_}�.wL.m���wy�����kb����J�����F��.�K��/\+=���%���yiݝ�g�����U�d�@Ŭ2�D�/
C���>�5W�\+� κ�}mgî6r��iX�`�6C4��B��i��т��6��q�4�wWK���n�꾮Mκ���(|���rgX�uw&�|Y���߯�2��vy~3-�=���6ף�b��p?��^OV�>��Z)#�ZR$�a���Q���
��g(v��.h6�.�^�	��B#��Kp �%8�A�֧�!�Q�����^a���oI{
l9������*C�l���k�����ar'0mZ�4�*c�!�������.J,��A��.�&=�~�HKM�6�,���"������� ����\��N��ɨ��M�)_����n�p<�%F��R�ؕ�\2�A�Õ2+�5�?5�f�q�a�ѭ�v�uT�B�K?��"a�_��q/4`��Ց�dT�b^�Lfy:�@�n1�����o�ݛ�?>6��f���N;�!G�:�h��O������-"�@'�y��h��h�>�n,�7
��E3R��q��:6ħ��E�:�}[\^�����.��D��'#j�asT��S�j�*|@��+~@��m�	�69o�$�P�u������n]�e���{$P-CNR�쁯�)s�j�r�/䚥������"|Y��L���jA��g�m!��:p��b�`���R�� ��g�n5�ݣy��l-Z�·�u��R�pou���CrZ��LT9��{2�U��;��g ��5Z{Bqv��ZR��(�r�Z����26xY<��x}��G����K0l1Y`����i�t�l͟?8M����������;�q%�+#��NF���9�a�0�h�4J�E1$j�_��hY�@�C�>�~a0���J��G�p{@I݊��
�!� ��}L�@T�s�{?H����k��� UR��ᦧ6��?&hBw�|Ц�IR�x�XY�
do1�ꭄ�I4uP�/z��|�#�81h���Bbߞ;V+@0���r�3$cbN�xB'e�j ��6�n���=�H���L�	�	0jtHa����>_j�_����~�����Q�G���
���6�?����@�l��$ҫ��7˞	d<��Y}����(��E�4�eA�մ^�Iu'����������jrWT4'x(~d���񏟓�#�՝�S���ӕ�A/Li��/��bů�T��=�lӁ� *���6z�3�(0zSF7��> ��lc��օ�'`��3�0fL�?�^�-q7��^��Xr;�s/C�C�*BH��C��H�S�[#HX?��ZIQE�/���O��F�u�L��R�)�e5}�����s�r�d��m�Æ�r�ٝ�������PXw��JL�)��#��P�-$��}���
�U8+5t�`�P#��,��]u�ц��+!���&-)��R�I�AO^�/����D+�bVC�;4.����͓�w��2�M�x�|P��٩VwE�k/ޝkj�������걜�!싂Z1h��!��MR�X5y�n��KJ�~'j~�*�񹒇i/�a��@�%�f�x�hbzE�	k����Qc�XxvZ^��\������S�~EL>���@������T�~(*�����K@{�~�^N3ĨR��%�A0�'i�x��*!)��şwS��&q��ѓXnS�k�QE�"���Q��X�]?���b/�(Է�r��C�fDR���z�v��u����w�{��SӚ��+Ԇ�흂����a���q��D�����!VFK�4�t�� e�Y�{�
�	G�^* �b����_c��s�IP�-���#h��,���&@��z'>���s���ZÝ;v�t<��?���2w�;I'��tur�u����py`��Р�C��T���m��C{y}�?y�;._����&�k�۶%�i�-5��(����p	'���P�3	46��ѝg�@�/⡄ߌ����~����Bĳ���Dp�l�)ܳPL4﮷��(#�zX5E��ֵ?��i�`X)��֮���2:��\�^���Ha�]hAP
�C�3�X)�hÂV�7�쥈��pΒ8�@ހ��J�W�w��\��XZ�Snr��p�]eE�P�O��F��gR���Y,�����=��?n�^W�ȶ�s�Ǘ���U��'K�+Ƣ��b�������,�ҹ�����o-�$iN�
���v"�\�V�,�n�x�R���S�ְK��,�x�}�w�Κ(Fjhx#�`ܬ(c]�]Ou;��/'J�B�ϸ���a�д�9E�L���cȷ��|���G��oK�����N����l�Iy��x'l#���>!4.u���/�E�ҎaH�}���L�ߊ�(�qA����
���-�c_	e�g��E���������Ҷ�ʹ�w1����*���Aj����U�-��%s��|�c�d?�(�t|�6�,qap/.�/�`aW��+�r��,���aKn\�Wp��R�і 	rԩ�.WQdB�A�~_V;W�;�3�[o��5�_�*W��R���4��W��p�w[�Ban��n����|��� �^���û�hqOnŕ+�4���D=o[c��d��oe�\ƾ�����U�8�mߊ�L�b��=��1�kV��4%J�t�w����m	�F>��l�a����g�i��9"#i=�]ob�3���&6�-��⡱�w�x�cG>�C&��9����{B"��{� 5�hk�o� ��JP:鎖f��W�����UH���2����x\���mV��tRo^z���H�������T2tO�C�7�@�,����c�Ry:��4{�g��TX�)_��'
�ev%�r�k&� ʼJ�bI��	u�y���l����@7F�e�i��W��,Y�sX��:O8.��������u�������\N��{x"��#[�t����1��U�Pw7_�	8�!t��g���2
ZO��}��E�6��4�e��B��>�j2Q���u i�X��*�-��!M��4����t��*@B}��o�T�`@dc{޷�i!.�T�����Fޝt����]F�&>�Nt��y�A��t���,M�"AK4�	���N.9XZU1���f"R�,P>{b�u2����/c�$դ���]���S'#wM����'9���f�K�Y�n)|�{�UQ�� 2
Ҫ�*D玴/{��n�d�>(�Y���~� E(����ߛ��0q�U��f������� X�w��u0s����w6q:�z�
�90/<���b`EȪC!$�������n�V�fNvx8R͒"ӕ�E2�Hz�࢙��GMq�B;�EW��qd�*^�?w�άR^�(q�N����ҫ�mkm�/?!*��_[�b�HE�:��F�ő͝��5lTX&fk�f�k/����#K�D\�7
u�	ʫ
��M��>�Rt��_p���N�ͫ�d$�����8���>����/��\�M����R�2�I[��T㒨�b@��Թ�l�9`���&��Y����U�PEċ�3q5�nV�_𞥞�|h��\�Xl�O��}LV-_��#���9N�� ���p�!(}	^DJ�O^���H��<����e��1���}5I���#a)6t���3���{�D,\�I�]���|�0�w>U!I����,WK>��e��W�\���JQ�@v]�����Ej�s����~�� ��x���H�#�ȭ�����b���6'!��3�$��7%{^	�}� ��S;'��&)�E+#��p�Rn���Z���u���c��`{��<"��	դj�n�8L5L]) ���	�2*���>N��3�0C��	�7j#{`�U�1��[�7���H�׈�[�0�����D��&R��R�31�fU���$`J�z���Jw�{/,+��>R�ZX��|�ekXP�:��K��.�ұbmy���q�M��|͛?C�Nk�EJ�a��G99~;n��2A��N�#�ۤ[c��ޓЂ&��.���_wh��M�$���zsG�ZU��`Ԓ%)z�o�Q9�2�s=V��U�$��s��~g�D>�:tpx\`�__A�hQ5'l�V���j����$>i�ڔ�vטSt}1�2�ߨ��џ���w��߄�Ԡ�~����{;x����@���=d��Љ����ה�b�n�~ͷ)ڐ��ƺ���*��0��S�R�?���Xk%]u�l+BҶ6v/2b��|�MWe�6P^o0E]>��ٛ��cP���)�5i�`�&+"����1# )��il��ϼ�=l P�A�i�*�e�oDj��_�'7#��*�L)�MW�+~�n��_9���qI��dx��Y�#�
�F�G���{�Vnp�Y�ܪDx�����n�>GAR�k���N��G��EfoQ��3�Zk�('9���p�4W/p�Ps�	�Й�$�'��g����/���m�9�ָ��*���4���/��{6�w�Xs�5UP����`�^�G�/��M�ѯ�FBr+�C��v:!�o�c�۳ဴS�4����Uk�\�h΀Ҧ,@+�V\sqB+:��Bv���: ��rK�U���HӖgG��UW�s�Ԭ������34�4	� �i���8�NY�W|���k5Pex�T_삺�/�ߴ�5��`�O�'� S/� /���)�$��/=�=�nu%��,y���+^S�hO�U��d�j *�1��$�m����W�F1�ܤd?w�t+o�)�����VI�]���/��n�P#�O��-����az<@ѝ:�0�;���*�vm�@��Whg��_�d�����:����H�+c�~ߔKb��h���'������k@քw����l�#��8�?�!>ۜv�8u/��T����5p�{U��mE�6��uǜq�S��(Yn	f��l�޻S��r����vb�3bR�Lg��Via���i��3 �����[��l�;�/�jF@�b������x����ʳ�B�[�l�b�Ԝw���6u���䯰���:����ŋM�e�V�YTLC�,�D�a+��/��&W9�y�I7�+����?	���k�Lp/�IF����n��ӣH�D��L�2
ٹF1ñ4������UN �t咓��m��W&ˤ	�O�h����+Z�*�3>��1G��$f�CGJ�)&�.٩~w&Ϸ� ��Ø[Β3�[���9���:�D��(��_c����^x0���G.d9N�]]��>��W����L�Yc�e<�i��0����^M�#]����>�e(4	-^��0�B�~Ҙٹv,�8�h�8�,����W�*�)���&��Fb2K�;�:��Axj@=���EG&�� ��K�"�Q�tx4�ژ�57�:��l^�&���>n��R(i�1�W�j}O v����@~�\4�l�׻����~��3�Lˍu��4�m��yǡj)���}mp;UU�t�v����<&����� P�cji��,Ĭ"�ʗ�	Rh,><a��X�8�흦�𔜾ť��1A
5n�Tѕ(�\"�T,��}�,dO�"3=��d�̠�"���V7��DB��8 n*�f �Ł�=I���Y�h�nNe@�p�E]��4!��R�����dx�h�]T{9�VG�|����M��u"�Er���K���d|I!��	ڦ|��'?���"��Jx�ˏ���E݆�X�T8�/n�@� ` ���V��LP�*N?�F1�y�z+.^���tG��z���V'��SꞩjEM��K'���/g@ks�5@@��!f��k�֔��,n��]��We&El�(�Ə�$XI��Yu�	C?eh�p{]�`n�����RZᒓt���\��"��z@��H-��Δ���Uz^���"��oSՖ�iG0(=db:�t���]/���/�X��E�\���(maR���~�|�y��4��3\��㹙lM:��������NG+�B�C�@��d�K?����5���l�Qқ�����qX8e��%�T�[n�N� �Ǯ��m���Y��f�(U���+��xp��-��vTM1m$]�.��g�����H�7�s�QE���R�{�=ژ�ʱ��N&^�T�JT������WB!��"Q���9]_��`t���@���*<ib�"����KA�ᅞyi��!�h�b�Jz�fE���b?<�2�B��|�^��M��[?NM��?���Vn�ޣrŴt�4.��s�[��q
I��k�S	�H��l�]w-+���(�W&VZ�95c�l��J��`t[�����Y�h�U>���T���Z��q��bWlo���3����m�X31�G-�	H��E`�}��v�Ϥ��u�Og B��)�ͣCi��Q蘹Pֵ����k��́h`I}�`���jb6R�ä�!���#kkӶ"��!�@Uz�n��ƀ��_$�6-���MF*�� ����t'E�O:u BP�.�Y-zq!\�^F�N&!R?	�g��S)rPf�n+�6Cg�m��a��ԍ8�G���Kܠ�e�����Op�����-��^
rU:yת�o/K�����L�{�����5uh��x�� ���g&��3X����ɯh�ȑ�Q�
���w]�i���һno��8�6�����q;�4!?���͚wX�S��&�Ů�7���Ws���v"�`l�bǲ�TұU�/9�v�Οt�M��{o^WF7,Fc5��wQ�v����3I�ܨ�`$i��`;�E2��Pcy�P�O�����+9���4����o[������KG{b��ς�<�אj��}{� ��A�$h�}޳<�%�<����l#<��79�3j,"��pG�wGs�w,��7K8\�T��6��S�(����>Q����.�"����2����z9�N�(��0��d�M۟F����=��kr��y�5c��.HH-��6�p�:D�+y��Êj���KP�&�5\�"�ĎK\4F�0k�6THb�vd������Mv J��G�u)�����	};���w���'uT���S��lu98�3��� r��Ⲁ,�9�!�F�ӭ���|�j��>Qa� ��	�UHjQ��&+>�7P]�h wDe�����-Ny��m�j��O ���|��<�J ����2ġy[&m�>OzkS?i�����ӡ!���h�U�%�5�G=����*��4�V!�-K�0��O�$���lf��P��3~���Y��g��h@"Rw�⥯$��<�e`Z~n{A4��y]ޗ�un�L_���Y.�`���вբ��$�{a�K�v��������I=�#\U�.51�̦�'q\uT(�����#bU"́���V�3�iQ�E4-������o��O�J��Bk���6� ��v�r�N�Z�n�]G�����ʝ����s�fE�`�Tl�;����Wm���щ��RW\�/kR猵4c�10ޤn����K�L�����El�bE�<�	�ej���+2M��9��eť=����2d�xĻ��,c��W�uu-I\�ۼV�S�lB*��n��5�}��pZ�r�(�m �J[�	���;_�����)�D��Y��9�Bʯ�m�����/�-^�Å0��t�@#��� ��E�����$VH�����jr>充Z6G!g�^_�$(u�ԉ/_�a�R��4{���o�y2�~)	������g3c�*�k~�"vi���
��j�ŋ���G)�� ',���_���aޡrE@�ҫ�ʍ����jX^��|8�dNg�d�a���R����}yR���l�7l�rV��<��YОl1��Ql��L!�&��ߟVb}��˃���
�sE�<�|I��;Ǳ� ���>�NRs�Xˆ�ʤ�oF+�?&�������~%ma�t��]�K���<z�O	[�'�}���h��`V�Vh1�*w�P""�"p! 5���Wu�yZV@p��:3!�Y����_���~x�i��qߑ��q����[��h��iG�s���d(d'̕9:H�D�&\��Kjr�%����8X]�)._v�j� �e���+]dN�D�Ғ�I�,Q;]1�o�ˊ2��I���M �L/,Z�v'a0�$�Ji4BB䈿)&�?�I���fA�e�?����i�]�	��o'�
J�^eӲӦb���!�
R|�ʯl%��!� oj���YQ�Kz�77�n��$�!���RR52�ܞ
�z��
�x7I�?�i�}�$��%��F9_�ި�����O��3w��q��R8�����sp�]������!����� ��0�a�Z�Z,$[�aϠ�Ozim��P�?���9�������'�Û�݉s���� ho�$��?�z���_�nn�j]� �B�����0gvz{ �92�/�����X�TBa;-�o����L�C�V�J���I�}p��hVGJ�j�{�}�̷��=X����x��>�����*h��U'�u��Ho3���QG�3P)����n@�s�8޵��>����>�͜,-�[,I��4�0yQz��՝�<L�jLe���a5��+��f���fO��U4j�'���[�{tZ/�?ޏƮG�&���j_�8Mwb���F+�o=w�d�/�*��_1�.�/?'O�K�==n2miw#41��xq���6�I8S��X�xH�I#b����4>���W'h��C#i�`-8;���5�^���>01���>z*Z����e�C��n������H���n��$��#��]�[Q7b��n�]�s)v%� �v�mr��C�zlr%B	q�P��+3銅�	���?����H�*�?����i���#���Xjː��b�?��cJ�6j2b�^�P>?;4��XTn,`�*ո����`�7�+�t0�ց�S��]S�;��ը�4g���)���G4j�v�:۹�'�rzG�7D��n���i������i����ު��EG�Ni��I&� 12LГ��2X�R�.��RH�����=]��kȓ���(����$�H������dT���Ta���T�?G�sE̊��s����r#I�[��2����=6J\|�<�Ô����!Rg��rJ��#�SmVO��o8"0�x�:oz�����.�"xS[!x66몿,0z&YY��LU'��<�q� �Y3��f_�*���h�
`�8�`�[Q��^�>��פ���y�O�Ė�Qx�=c�yq&<>�af���%�&X�6n�,g�r�~���hLX��R��Z޸at}�؃� s1!�!�l�KH�Ņ��,w�P�Nmc5����m�����W��7��l���ؾ8R�����,�i���-�~��l��Tj��KW],����ߔ��K��P��'?rZu���z�t����� a�6o��S����A�W�T�O2P}�e��+����a�m�a��;���u:�q��=P��� �f���y!�v����/���H�;4�v��z�M�������4[=�J͆���x�ؼ&������Z�y9<������r��R�7K�*��:��/�<����b"�.(��g��%-zw����Њ��
ysCv�)�[�P^���e4�	sl�B�o���&$���L$��(�V�5b=R���u��n��=ppWT�u�N�T{�R��}0������kQ�1@;p@�d=��BС�����3*C$�.��Z(U��}P��4�'�3�庛���^��^�ab�;���t��"e&a�eu:!;��<vK��Z݉⎹	� Q���ص����w���T��#ߚ�6.:�7�� ����#���L��I�[��Uw`h] f��MrF�r�D��E�X%G�iRZԖ|�c0�{9@��;�a�]Ԫ؁"��_�!�aY�Ǡ,�p�Q�}����K	����M���$�KE�O2wn �)[�Rp�܇�gr��������TmW���;ѣkz�ذk���"�
O/�{�`hm�?(��>����h,|�j]�y��+�4�<%��4�2����
�[�|�M�1z�8�/f)�b%&�u0qVVM/\�;C'��!Yn%O��Cjoq?�)U4w�^e┳�'���Ő���l�M+��a��#��fa=A-R>D,���ݹ�ڕ��_۠��y��|v��#���y��2M
�UY���4X`*Y:k��w�h��1�����3п�a ���5xx6�".ŋ�����ˏT�V�0����@���j�������|�Z>����7��H�6��xӅ̈�����Dd�;y�#KN�1���2x��ߠ"RV�� v��O,��Cp9s�i�W�/\���߻���dV��O�h�.{���\γq�O!��G��Uo7����ii�Y�RX���!��6��b	�#�pg��pս�� ~q^��*�o�cv��52����X�R�w�~�
���^�y� ^��ݨq_��E>��y�m�;���?{�Lm{�!�y���Ҍ2��/N��> �����:y݌.��:y��&$���-8��������9�[]6�����ĉ�RKk8�hM�I9x`K}N-�Ì�鿊��;N�@`86�� K��2nHt�(a�g.�2!���w$�7lW������ï[ 6��'��"���Dym�WmI�7�S��x��r^*�e�O���}�Q�)h��1���������_�0��a��W2H~��5{xx
���dq��[#�؉g`���	T+[)�8ER#�o�o�,���GTO�h��"��>8�\Uz^�1J���I��3Ӟ<�\5*��xT8���kd\��s�0���`/�m������a���q>r0��#����4hp��~ϸ�2�-6eH`<Exj���H�a���6E��+9n�]�� �����|о���!(sf���}ۗ/|����c'�nAV(��/I�-#_�xC���h�� ��O�|C���z��Q��� ���X����f!\�@�x"o<�SD�C&���A�#�0YQ�i�&�r���)�D565M��t�ܲ���!<c�U��Ou�������D'��H��E�g.z1��o�ң�p&-��}'���Pϗ��bR@�رJdH�ubh��z�2�"�����ܸR�P��v���p��hحiĉI����·��+%��&��x�u3.�����B:�Kظ�.��]�d�(���ł��DԄ��:+��,G�ܶ�n֌���R�f�۶| 5D��&�4�� �x���D	��zAsK�ˣ"��79�}?���5Tѻ���]��U��v ��%�@\���5d.a�,QZ�sU���7܍ϗ��\J�㕼xW����<E׮��Oi����/�?x��K���}��q�C�nhQr�Kz��1���C�����*t�<P���?�}�<4��B�ϗ�lW����p���<��2���;!�����ַ�U�n����;�vQQT[.�_N"TI�/���i��4#��� ���N���	��S��/k�#�y~4)���H7g+����5�9
�	u�Rkɀ=m�u� %ʁ1��ƭ��� ^`�j����h8�{h�]JAr��BEy�~ɡ�ƷB��q��F'A�B��eb,���(ó��G�f�;*o�/XL��;�n��W�>�t��-���k$E�9�S6=!���o�'+̖�2v�ӛ���=Ͼh�P���(#~[N[�Q�g|c)8� =I��a���+��!pt�`�mVc���g�e�=<>��>��E�z����õE����&�Q���ų*��e8��i�5fj,���fOFfoU���M��6IJj��$�gCT� �O	�O�2�'���`�p�H���ɃkS���xi>���C�ѤaJk9\�{�>��Zٌ�;���-�G�����_��'A�p�ƽ /vl��x�w��yഹ�6UI��7�n��K�v�xO��!���U��AL|_������kd��ǩ_�Ή�Kk��li�S���&1��a�ɜh��CiM�Ϋ�|��R����o�z��Y"�6E����j��(���`��)&n3���݂�~�XB�*�s��%�" e.�σ�ݯ�i��+P��K9*}0S\�i�K�l��y���~Q�	LI�>urK�'F;�O�|�τ�^�@�.� 2`���~@膄2'[gF�M_&Z뭋��L�Eϫ=�#�(��5p[�/ӳ�k��R�����VD�u����8&Gu�=���%on�D	N��w]���(w��%�-�ͧ��wm���9�W�Hn�&��3����Zi"XI�:�"���\i��ϻ�@yL�����I�14'g:��wk$�GόP�����{����ry`0Ϙy}?'�5��*��;5^�Ydj/��{��c��n� 3�L�#�h�ew~��۳,��</$t1�n{N N(7F�a���$R�?S�P�K ]֦՝3f���i�#���I:�p��"�"nЬȳ&�mo���g�9w�:��#9��'�-*��[f@)��Uk�tV<�V*��cK�F%E�k����K�S���gu%ښ(�G�8�E��]���iPl7��n�	{��$���&V�HG�O��2av	�����I��
؉��iy�?�����ȇ.-�;1ks�^Od)(�NHZ�VM#p������ܖ�3��E���j�c���ְ�mS�۰�%�v�9m!�n��|���l�����ª?�`)�\/P�bW���+�Ԥ�8�������7�0��z0k�W����%�`��Wҷ�d�@K8����vfM�Jr��	� ����u��i+�#,eI���w\�C��`�t�*� D��V��G{$%�G/X{�0�M��'�f�\��6�����ծ��ݔ�B��& ��>W���V���0���� a�E��T^��\�-E��0Q�}y�KЅ��\��%��=�M�w���mu��cH�<���gZ/]��`� 
d*���lf�m�f�f3�?��%�JpNxR�\R��X�T#	��(�l&ߏ�.#�Xn�;��������G�΁�UG1W#���#��LV���x���-�W��bp�>�"��r�`��uTgg��h��c"�����o !��G��X�@L��5�.G��Ag�b�-��f��+'X���O�FXSx0�¸�}� Yqrp� 3`^TK2(� �C!ܼ�����`2桥��T3�����J`����������[H��H�D(0�{��k��=��X0����&MAx��M1�睭�[o	t}�xa�:{a�w�����m}¸;I����3��`g	&)���ķ�� !����2�Z��񡋔1���z�2Y^�gG N��^����w��0d��<eX��ap�h$dш��-/� ���6�`VV��[�ݓ:<��"��0��]x������	4�ݧ��ܯȶs،�君��X�e����2��a<dҽ&{��L�ȨM
<V��I��7�܀ѩ�r�I��x ����[*��s�{� �
�G�`,@���&Oj�2��{Ә�V��%o�zྕ��o�ٵMWR��V��P�vK]�%'����yZi��|x�j�_��S��U}>����"�s3��G#f	ת��k�R��,lRG���'�<�8�J_b5��3B�S��%�E�����L�J���1�de����[��D��&ˣ?|�)����f#t�5�0P�(���{������0)B�3��nH�0T�>�s>s��V�ʩd��4��A,�J\"�oSH8��jB��=���	�BQ]6���M���
U��B��fSp�)���֠j���$�E1G}�����������՝�g-��J}6f���u�j�v,Տj� �Ʉ(s��r8���-��,����7����3�ף���.����R��`�[��H�&�a0�h�Y���9�r�����ʊ��)b�rK�	�TA@��-����,.��>��Ӟ$s��3@��_��]�/[�gSQ6����d.@�D�`�g2���ƾ�'�k��ۻ���%�e��j�����z�QJ����1���|��lA�$g�ʴ�~^4�"`?id�IC�
��{ Jpז�y�nG�۽v)3��q�N�xة��		���"~юC�=��c�L��/�ڌ�����p�xb�VO����(���y�t���o�#��BE��{"��"b��<*↸���\�a5�':�4�|��J�^����?���b�pY<��Yʄ�v��e�Km�{M~�����fp>q��皾MSH�U%����D/�2J�8�Ke|�5��_��H��>��S�v���&W�����*c߆���n�麥;�V���� Av�y�QB?k^QR��75�X�m$NP�_�y'i{OaR|�^J�IT��ɖM�뵢�+HC-J��S���l@�:K�unoh�r�Y�v[)i�Ӏ9�|�{����O���βpwZ�ӽ��u4��vD���&�N�Lm�G4��Ȑ���{
��Þ7]w�^�ө.ۦ�N)����"�e#绣�Z(/t����8P��|�<�c�[� $�eσ{�?�fN����D9���>5S �c�
܎��A���]H��3 2��/���UX-�/�;$G�/ N�e��
�y�
�����zr��N}/�@���m��L"<ginPH�/kQv�7��;~�2��x���T��2L����4��{2�&���>�J�\f�M�j���iPJ�?��K�: ��ː��i�J]@���r YSu���y�����"þ��WG�7:�!U^)U�Y6984i�#.E�e�9���"��=�ǰJ�Xd@,D9\]�qWHT�sc-�#����>�v�����çg�D�p~��L��ǯ������ѓʆ��LnR0��̓�O|���2ƃ�Q/>Κ(�96�̜%'����o>�H���2�z��5w��`8�)b!�~�a�����tȋ��Qy��|�u6AcR��;^[؎XP�����9:ԟ-G�xY/���>��E�&�GB5��AE�څ�i��/	Hm��7c<���cS	���������1��ml�E/h�PQ��ڰ�I`�� .�n�������i�?�z�)�LKD*���!����GC�R�K	2���d�ۜi�o�o�j��ߚ$�����{�+�K����E��ljw��M-<4��2��7��%PN�`�wl�(}J��\2[�'}}�,#�&�D��^BeH
���9}�Z 93��%��NC��}vҭ!<�](�)^sЊ����QE�Q����;��2e�0q�$�׽l+�ˣ��c�� �����Dzc�3_�]�V��J+cT���/���l5摍R/�^9f�"�A�(�!�L���M0 �<�ţ�9(�r�h��ԙJ�Zb�3�1R�u9u��XC����A�F���a<_8�N;���I|<�|x�s��߾�rv�zŭ���	i������?=Q)��$$���`�����Ј�Rº�w�#�,J��čaɛ][�\���P[@�� ��G2
�]xէ���ꛗKұgc�I��7P��ֆ�vP�r��N̞��������L�!�/��������2se���E����Ę1�.�{o�D3���4���;���Ev��@��I@�DD�v�%��xN(��&|zQmA)\kXR��1f~f�2B�5��l�y��������p̘tw \T�U"����`l*��-Ҷ++aX���~j����^H�ݑ��[�����,y�������r~�%U�OWF �����O�ϔ���,~0��I4�ϗ�ȥ鹂M�H���B�3D1Q1�܃,�oXț`�bi�.}!W~��k�s�"�,�����,�16!d�'+<x�͠EHe2�����)m�>^Y�Pbc�Pn�k>'��퇪�aj�[���bE�0��=���*�H�4=�R��ޖ���y'�]~{�]Ir��e�p���rB4؍�Y��
�|�a���f.�+Ó��~
@����L�H�{7�*���
i��E���s�+���a�����T��[<���P��>���/ ��i�O�w�/."�"���yϘ[-�F	�q�(�э���rA��W���_�ǎSj����y�4��{%`��)VVW�65��HbnZ4�l� �J���*���;F?ce��_(0h��x�ք_2���8Yf�`�
�B��GT.n�6л�b�����j�d~�\ߟgx�kuc�T�+���<}</��$� >�#~K���P2e%Y��6���W���f����O���zdTQN���Ow�{�	7#��!@���gB�u��sq��r�a�L�]��HLz}ZfhN��b���$�ʔ���!%��-�W6��-H�л�3R��}km�\��i�P�C�f_��m��c4�}�am�ʪ�Q�[Q��#��l����	��J?s���D�m�mԶ}cc�yy!U���*�,�I&9#؞����AKR����چ�ì��H����Fe6����������	�xN�i�oRO��b��J �ޢ�<�|���6���nI�{w�UEP�jӾj+s��z��� �*����
�������tJէ;�Y��̍�2��vW1X�)������Zxm0���D�c�����T������z
ULGTDמ i����X���)��Ƒ�G;���#'
G9Hȗ�2��$� �Tl�Lʸ(���@�tt,tY~�C������P��ƾ4��-� &jH�	�
=�1'w�\Y�|]'0*R2o�������@m��9�E��m������%+ޢ��q��"m����a$�ȳ��n��@�g���^���#߃��}x~�p�*�R#�h iW���_���M�A��J�M����<a\Y�%A֡�����㤖C �+���l��!�jo�{�z���Y�s^bc�d]>s!{zg��]���ҷ��k�1i���߫��e�b�[����������9<7�E9B�1������Q�5��#�5��A�ŉ��Y�&ɨ�6)�+p���뗂���������kA#8��F8n���������ه�΂�!2�.�eX�`0;A�
d��L,���pɾu,
�9��:_EL\�̡2�s�a�k�c��%UiR��@k�U�1��2_�֒��mtk˅�F<Pm���V�̛�#�ß�����)�_�����o;�m'��On�̴q�S wc�ާ ��1��aI�*�ZL�~���1��;�`�A�����ԩpFqlP�
���K����?���u#��x^m��Sٿ��,<�������ʈ��)��X�}��y����`����m(�sj;����JxQ��?��3���[�.��B�HטIQ	�~+,D�������tv��+y��q-}̂5x��p#�~��[�׿�CE�������N�����y��`��P����SSQ8�֔�S�gu���H�H�I��_��(HQN���	?x���l@�w����{!���n<��B��h�l�:r9CL��i�Ծ�\<n�č�u��q��~���2
�}BO���(H眝�ջ��QMr����t?����@�5ϼ��]��DN�q	^�YH\%��Ig̳������1�H7A~{��ɢ�],�;����b(�ᶿ��!n֞�/N�F7��R��%�_$��� t�l'�����S�pJ�Ŷ�(�>N
�N+�M�:\VALG-��vP�b�_�.gZ\3=B���@ �x
ܶT���S�������5��g
�%���yw��,.�z>�z~�L� �R��EN���,�L$?X�v�L�M���'���IjIpZ(m��!��Л�i
��i��F�
�w�ᬘ�%�4�	e��H��:Ж��^����*#��W���V�dH�쭮(il��H�1Qr�6I�1Z+��	�ܩ_,�_�.8�5��5�I�����;(��?�ɏY�%`V�L��c\SG63_����<W��L-������d��]1vl�'r��s�Nu�V�}��-G�n��M�����`��^ce��d0���a�B��2�^�siUW�e�aOU}��e��)�`��Ҡ� .���P'z��qQ��0q�=:YI�S��E/���4�cV�k�۪pӺ��g��t^���}A�>�����-��O$�`��6�5�"�VF�U���o�¹��� |z�؏���[í�NĶP��I�ߤS.
�n=Qu�/����)�伤��S����,��M�bt�(k�}������o��v6yM�L�F�y�=O�\�jb�ǠB�N�]����O�o']WH��ƈy����K�"�i�	'���R0�dwy��J@���U�~�����O�Me鴶hd�(�(>�Q�}�yC*��?� ��bD�VW����;�q7��ev�� �9��n{��	��4k�R���[��C�/�z(Ć��!�8j��%	�/�#�E�IdS�AY����۔�i�����I�y�!��W�ڼ��V�c㭽�1���	X�^H�;y����]�c�yiWp���K[� ��t+��3(?}�-0
�õ+mR�o�h����䓶��-���/-�\�T����Ĕ�2d��:���: �w���S�����xI�J@��ϩ�j�i�����}�hi91�iB���	��vxb��~���T�4b>�B.h�b��T�g��:M���InBݮ�����r�[E�oyꈖ�p3��o ���N��x\��b{nw�]���٩=<�>h?oX��@�&����j���
Q��s}}��c�"N��.X���lI�,'�*x����.~�d�ة���vfF����,Pq���0�F`�]�x1M�={�Z	'�$V*�]��������C���H�f���@�{(k�e/Tp�>�3RL2#�d��y
k��H�UAGJ�]��M����n�rP	5v]��|l��fA:j{/֜Ms���*�r�-Jހz3 we�0T@�:��%<���9��jGվI�]��*&���ht�옇�||��Ao?��p�qϹCC��?>cc~�x�g!1�/d\HK��d������F��T��Xu�-��>w�2X��ч����=�Ĕ��:Ϟ�g'`k�9�.��7������|f�̽E���WrM��z�2QF	 21��SO����Ps���z�n*u�#;?�z�ȳ��҂:{���z����p�FOjgPHFB���%��J����!���|��1u���Z�ҍa���c`P�\��c�����KĞ�e�}�S��c��@�])Ce{��~�T�C�Zv`R}t,0R�D?���G�G��ힾ��_�X� r��X�8"1�`��ȌV��� ����L,�k!�lw�R@�&��E),�����O��;?m'
��P<�/�Z�,UV��ܣ����s^���RM8�r�l�!dAf�΁��K�Axz�%�r]5`���]�����a��D�\�Y��#@���l�iY���=7����x�[k�cx��ی.���p������k�8���UZg�F��)���yx���X(�
"yO�Tj��n7m�cJ�6��p���>O��%#34�/��@�t%��i#���-E5b*�9I�0� ce�X����O7(��<��Y�m���w���Ã�	p�2$�w��/�/���`���W���_.�<%)��0�Ė�f��Kg+E<Э'�y�R#ȸse��'���{�R�[����H��8�1��گQwG�D���������s����������5�&pdS��R '/ۏ漮O_d�/HRv�nW�".�VE���iR������:�M���	}�{��(8�/��	������ݲ
�} 
�F�4`=��xz�?$uDa����0�����Y����U�P���n�V,Kb#��M�z�'��p�z�u�Vw44��DR)>M��((���o,��-�Ih�ǋ.��1R�N�_��#�U�F''!@��6KFE�8��2���v�P����B�JB����a����1��Vm�s?���ZSR�1��9��������;lZ�%�����U�v�L/��:r�|�6�s�Y�ߦξ����Ru7VSh��>x�������b.��#�g��3���:����d��&`��=<6���q�w'y�$Gj���!y��4�䌿_U��e܈���z�5�W|A$)O{�`��N������Sm�U�a�hpϖcv�w*
�$�z��g��<���I�[��k�����|C�]��?3�P�Y��9��Ԏ�eÆigU�_�Q�n�:��C�� �.'��'�$̮�U�wͺ+��n��ߺ�>�h�j<�r����4�$�EUp���g��G D�ۏ7$�Ц2'Zw����K�nv6�&Z������$t��_if1����n�.X#�v?	���W#�o<����@�*7������V�� �7��3p%]Zuk.cF����k����W>����\<�#��Gcܚ��ɒ%��#�>E�a�+r�������z��b�x_REi��iq����GUF7'�,��r�����Z�� T:D��f`�6Z�� �L?���u-`h0OR�3I�uP�l������s�n����F`I����ȃ�R��<^Z�f@�p�����D�iJ���1����!'��M9.� ����І���cO�=9�<h��%ʠF0�IL�n
9����}q�Z�a;&�/d�^�	��Y��Ң�Cnx�J볓��� H�c-�%�R% $��] w^b�w�-u:�L���?M���1i&�K���圈U:�o��D�r�_��c�?נ�5U��.�)CQ�z�(S�7]B�Q��������T���`��j��vћ�eMc�z�Y��0�o\�c��)�������|$�(��	�Xo�ռ�~1��"U���bɉ��HH6�{��0҅Հ��^A�,�mXS�;��
mK���ㄝ�z��z�H�<Wt����T�)9)�5َ��=��ג.������:d�h��V����l핓���L��|�}��>{Y�Y�YM�{t����{zS:�9N.#�z�Oف�������w����� ���,�����+���<��g��?����&�A�Gt��΢s;��Af�W���0�&�_��1��-��bG��O�)I��$�f��<d����F���>�A��4�7�����'����@�2�RET!��j���$A��e�nC6v�O�[�/�T�	)��o��9�ɔqi3�3�'�\�f+t��ّs$6���yy;�9�<1�%��K�a3.v�Y����:�ϐ�t�pF��`���nG�&��+��ęO�Q�=zH9t��-��w׺ r��Y*hr�fS�T�^�$4��`AQJ�u�<�2���A9�Z�ӇɪIp�=����{9�ѐ�P#rO��9 �	7�Ǟd��?�V���L F�� 3��ڥ��g���yN |M1I� ��;��n�Q�u��F|�8���j�a��P|�/��k����yޤ�b٫�$���p�"�/v4&|~G.�/Va`/��&FB��1�sZB�>�V�?�.y�X̩�;�ԥP씕Q�$\�-=M ��	d��c�-�� Q�V�0�@�zrQ�l&��u�WI��Uk����U�w�*�td�f��N���.Z����J /�؛�)?/	��Y�L���]y�m{C`���Ĵ@&jr���I#0PWB�� 1�s���Y��.K�0Y@r�tg���yG=�z���P�1GkÀ{��/~5u:�z���1\���o�����qBwa�ی�4�t�m��a�[�Wj�5�*@�S�0�?Z���U�=߷�xp��)�t�O���ɡn`\��RĔO�ܞ������m�hv���<��@���q07{��a�S�l���o����֭����+'6��^?*����뮨跦N��]��-�&��x�d�jcRi��26�J�6�/�Z������~��xX�?9]��}��{{NM�	�\ߙA�W�A�_6}f�S��t]����B���,TN�as��)2�K|K���e�U �e/�*��j�M���P�6V�eUdf����`.�#hk6���}Ŏ�g�\t�r u�Xk�m��̕��\l�2�R��K8��S��")�%��%���T�UM�n��F�	�v��Z�S���X�3��f�A��܈>9�LpS��S۹��PG}\��������XU��B�w��X��Z�S�uOT�[�q|�C^�������
���@�o��������}�����ø"��6�Z���#��\���e@���RA�n�y��	u�n_�h�|c�:��mAw�(ȳ��� H��y��{�%*����3���8~՜�-�s}��*���������b,#(��E���C����(��ܿдaw�6�#�~6ȁ�CiJ���'	-�'�Q�CI���
H��r���Q����B-�tu12��Lm]�D�^���]�5~W>�[�1J�A��������8h"�2��l��M��i����%	QZ�9ت%W�}P�����s��`q`�� $V�����0�������f���r�[
�i��	X�nc��}�L.99=�M��K̍���D�4��A�=o	)6XLo%r�o�5"���%�}��/�����2Ή@ENA�:�ߐ^�a�w�@�/��a���l���s
�&RE���д鎀�M���j�1�s�%��P#d��PR�s���.��Vp��r���tp �01��Ѽ�,�ip6�x����ƿ�B������Hw�[�</R�+l��.F��v#�Qo<h+�ߚ8��!R�t�M:�D��T�1�����ݔ�O�3:��;Qӊ$r�>��u
��3��,�o4*7�B��d�+���a-A��ˎ�ۅ ��LY����;����/�8�J���IA^S�\�}ɑMt�������Q�?��F��i`��Vp�Y�,�[Xz�G���u��sUu�Z�ªaS4�L��G�5�0XQ���~����Q��Bnږ��7����7�Qi�y�Wn��-�q9���G=��]��������|��k�Se�P�Ӭ�ּ��FƵT��������<	j�aj;���Y�*qZv�k:V���������ۥ4�j��M����1  �j\p�/��pޢ�Q�R�	��ù'[9�iŐ���_~ـl�I���!X��z0�vF���yu�Ul-�Yc*�P���m뇤�����~d���Z�4�F�0���
zr�e��9�d
e�o�k|�
�YF��n�շ/����s�]�S�z�*�<.QQ��OA�o��p;w��"�>΢;Z5�uF==��X6K��ާt{8���V;\/Ep6�Ӡ��Y0�h��L |�E�)�!�A�EO6�%is�F@���8�͖��@��~׌��;�#r���#�J����bX�̒fנO�=�Ǣo�f|�j�9�=gl2�s��S�DΖ�Cb�`�44����?tD?M�ӷ0מ�/m�n�l��8==�T��o��H�&���}���3��Y&��+İB��9ѪP�%�^Zt*;L��������@�a��z���, ����KJ�L�Z����6��eWI68LL��'���+5=�֢gc�'\����Y��/��H���8c��,�u#�O�2����aߋ��
�r������B����2��H�Պ�49�
H��1��S�ۈ��9�3S�&�ă�a���l�V���MFh@�>�ZNŮ�f�M�b8	u�&���5�0��W��_��;(VO�G;�U7Gy$]���;�e�\�E����;^�L�t�O���Yᝄ�����d+�t4�2�pW���я��%mR�P@Z0��)61�׻�Q�g�s��U5�6B��#m�6�)IB��c�^��f�S]�QWOd�ၕ#磮F�]�5�SV��q�a5}����ʯ3rX�<聾K�X�4��W
{�fL9��I��`H4$� ";����] �U�h��䱸��|X]�B���^�8����#HƸ�EN<�(�\����<��|k. �)#?��
��@>N;��9�!j�{����[=�4(��{_�8��#(6��L��UK��Z�~n -�N�A78��5���4q��$��N�|�fg�u��T����-C;J�2.B����Iz��'�B�x��8~��0^�;[mᇷ@,7é^9k��=�!n�c�./*d���F��o1!��i[!V����)k�8_�oZ�d���j㰡~�E;q#J���C�t���,���P�񤙋��4�B�I��(��o���aĤ����(���5�	2s��"��<X��I�jr�t������n=7K�#�3 Ve�
]X�q(�~}�{ԏ&��av{��Vn��h�;;B2����� ���;O���>����u�j�3 [ۼ�
����~Q'3b�I9����
�3�^
�����C)Y_ �r�����#��y(�V������O��- peM�pi���>R���9�{�k�D^(z��0%�4@p-tL>͘R®�9!Bl�e��K����,pt�'��l[���t�Z�������I'����:����y}�����JSw��9R:�ɵ���bU�:���$A�]��&@�� ���#Od툚� XC�X}���s@,_��}�F<r�%�(��t�F�ޭ�4������cG䚜}�v^-�7�ӂ�Å�0� 2SO�R�֪N����!8��5H/�˄0_vJ�/�!�7�"{0�ק���`��Iu@�3��d�Zb�[���<�8M/�Z�$����e�js�{p$:у�P��X�: kO���Ν��%��u)g�B��$ŵ($Z��&���/OM2�p긏o	pU���Eu��Sйú���L<̎g��)+8��y 3[oa`��)-�� ��W�"����2^YD�"�:��~Uҿ7Q�����y����T�8��źEB��y�6+n��e�\;Mfﶈ+s��
t��C�2����6��߁)
�+a��$��n�?xnj��0f��-jb��b��+� <��8C�9�v����Xb��q�	?:��S)��U��]��K(-�h+��~�4x��,N������mh剔X��>;J�0�qn�D�%Gs��JE ����v�0��t)�d�_%c\3�ʥBE���G�V����Ŀs����/Rȃ16`��0X�t1��!b�D�Fa��"����u�5f��O�_=	�
������Do�F}#}C��Ss��)�4���9�3։����O~��4�y3�����.�%Z���b��=P�n3C�]��:�@z|\5�o�"����kl=�����(�8ˍ�����ₜ�<D��Z(��*�S��D�֬_�� �l)��}n"	�^3B]%��?��$�i�+r0kg(�L;�Xl_�u��>��	!���\�9j����^�~�~��{�~�ez=*�����W�[�g��ѩ7z����va�:�u:��?w/�}�;uC������sFO΋�ۈF!�� ��Z�|;�9FP�Th�]����d��=�g(˲�+���?M��حxه�ʐ�L��[ YQ���gu��Z�-4(0}��dI���G�ڋ]�ꮎ;#�.-����x�*���`�	�~���t!L_;E56��a[�A�y�>Et|ɨ/,;��E:���=ƚ���'.�����ԧwD�l$������'�ta��v������x㢸���H��[ܛ$ށ���_�8+����n+�z���yƹ�r��xG�vfI�)��5�2>�����@1Ja��ӑ��S��!����'J	�ґ��"89Zv�Շ��Ķ�+�j�Ǵ1��V����1�Ѻ�h@����Q�$��4�sty$�M��Ϥ�h�,(W��Oj��
i�rЀ?fjw��&x%���n������=�����yp��"���'6Z��y<=]b�:5���^ꉛ�����`v�~�a Z*!�U�?鮚����Ԗi�B\����%'�ZG"�eqx�A_! �%���Ӱ�ܭD D �`���C��;��a�o�O'��$wo Su*q�?ffǀ�����s�Kd2��%r�{v�K�:�7����6L���XŇ�P�%��R�_k��<�s��5�{/cC��0<�F�`R��?VN5��S��;�$�[/�^C!W佑"��� %��,�ߩ�c `iGvD�0D�i��31t��Pa�ƩЖ��:b�ñ���$ts/�O�A90��k�H���1�@�
�8m��T�T��Z�ȿ��sh�U�;�|�����x�.ئC���G(_��K;//_�vk������=��Vp�K�1d}m��?zl�#u���|0��}U��b)V�i���M�]4�G�����!�.#�Y����_qO,��j(�}1?1'_��7�]Ô����}����:a��n�oe�խYg+�;��j��?W����>��@)O� �ϱσ=�W<(�:ξWuxcg�,.�s�d!�ǉkxp!fͺJ�z��η%��,����ӌɼ��2Ğ#�o�&]�B�ʨ���C�߿ W�K���$�Gt� ����%!��]�sH`X�p�b���
5��P��C��%-�@l�>�	>-�i�>qC�)�Y{���mZh&�$"���JP饊iK3����O�Ӄ�u6���:���̖��&^�q�.�fM�f��@1%���)�]G�[NN����VK�~W^�_-H�9<�����m���-��:�vW�$QgH5J7	E]:Y��jA���N��^P��;VK?Q����/A>cx)C*��M�'��-|�E���1ph�x�~95+�c�Ψ�3o7��.���m隣����`<�D��f[^!��=���Y�����U����w���d3xU�,�݈�q�E^z܎nu�`��L��ȫ^lN��c?rUC��[�ü��ʱ���K �E��]�a ;ŀ=rqߨ�y!�#��j��t�����W6�|�� ���>�Ȱ��,������Qy,����xW�����:���JC�/�ǤqH�Z�E�N���Kʐ��	�$̯5�GE��N;�i4���C�SKFU̎�����#�N��� �J�#ZP
><^.Z0-/�Q�ԭD�p�0�le�G~ӗ�ha�=���J%L���e�F�A=���A��k�@��S��6�	��7e�`��P3���ۉ��7)�������8�g�H�w�����[:�Y5ݟ����=�U�):yY��rg,�6 ~`�BMX7*	��:�״��������9W,ڤ�N�	|�&=�4�/��{���'��W�E�$����rAmyiN&�õ �yj��"�@��b=)�[�/kɗ�eH~���y���m�LL��^x�*�e�s�����b��������N�H�����ʯ�}�Pn�9�ζ:c�A���F�$�p2�dX�d <#N����bw?�3��j�<���ڒ���l������\֡����BXy�H?�8KnЩ��%��ܓ�5,��PxNO9@`�}����ț����:�'��t#���qї+���w۶d����uĻ����<V3�Oz���7/��@MW�7��8e�[��@��qt3�O�݋5�����,MK��;k�����%�7ѓ��&�1��P� PNH��}��=Mt�Kk��"`��8��5������~�n>Y��f2���Q�Ԇ�U$q�ҟs���?����k�W��7�g��� �/QE#m:7k��u~&�z�� rQ� ���u��O��z�G�)Y0�H�mn7��<�q����p�膕擺�bYl�MU!��E2��yiW��T�r�ވ��Y:���WB�8�l�Zt6 gͼ����2�@�����@��˾���ɴf��p��v�'6����F3tnvS:K4���-�tE	�hZ��c�Mr�2��F���I\-m�V�HL&Yka�CI$�$3�;���W� \5�T�eF���=�ݫ5�,�L��T{ɞ�����Z�dU�68��<3r��/W�X���V@�J��?#)&wHc��G���%[�%��J!6e덠�E�����P���N�A�4i"��}P�+hu�y���}]>��Dt����
�(���[�*�4�C���4ހ�I.��c�^/e�����MSU�"b�s$�� �Zd ����.E7+�Y�� �q����;9�p�ɯ�������GS��J7{S�k�D��
*�
�:E�@,<~���Wu0�K@���#|�ހ$Y���:Ϣ��:Cg�POU�g6h%BYjc�1C��7�Y��
\�4���9Ы�;���T��.�Ţ���	�}uMsU1$��bd�Ƈ-��k��8n�� 0jx��y���'�g���<J�z���E;�\�G:�$'|��aH)/B<����G�M�����	�m�o.��V���i�dǽ�`'b$YLX!�Dg4����俅E���A��=��"J���t����r0��ϹMF't�LA Z��Û��6����}u��Ѝ��+���/��<Ƈ��	:8��R�N3bIhص=n+뇁zV�%S�ֈ-Hv�N���}kb$�y�7�y�l��	���}����q��b�����b��KU�j�$��r�x�S���Ne�:4A��7���Fv��ʡ�3���҄�8F\7<��8o����q�͹���,�?&�t�`�i+
"�"�_�;���>�))��L�爐�p����E�R��l+cv�A���W/�N���(���Xy���;�f���rJ�*��-���^D�s�ěcv���]sa&�e���-Dg���_�BX>�!����	5C�i��Vx7"�ۅ����)dX�@p�t�5V��(7�T�w.����0�D*�������\U%Km��#�Jֺt]��4�douސ�_PM;��nK{E�kݑ�drVR�:�hxu�ځ(��bo+r�ɇ��lS:��)q9� �S�G������`���셴�S��� 	t�����.�{��ya��p��H(�VY�l�5��=���������7��A)��g`J��ˏ�}HsV�/X�J�[�5 َ_�5��+4�*A2��K���4���p͖b�ٖ���Շx@Rkw�5�C�,�M�=[�l������s�s���ɬ�߇Lٺj��^T�@��09,��7_H'�퐺�)H����]�*�`��9b��Ή�����������ɻ�<'��qW�0�R�
����>)��%�"�"��h]G`E��"�DD��fL|uT�P���c\���WmnB �md���[�6Qy�^jܲ���:,g˖����)a�Mf����#K@~�h����X`�J�W�9�Ș�fi�Q�Q��#}��f05�&[��X�A��jnn4C_�WS�Q��$��.%�v�K|]�4�&��Ӎ�;��?|x�����3�� �fL����"� �CV��` �Jf7��_�f[*7;$+�Ikg��x�}KlT���F�6��Y���4Od���m�NT�\�7�����u���.!s�0��O�l���A�D�r��s_`K���f�L�.���l�x8v�pqpބ�N�bϿ0���5`A�=U��U���2��]�??�_�y_��5�HՐ�d�a��ݓ����z*:0�٫������W[�a�0&���8{���c��V�F3z���qˤ�n��i�}]�����@�B�F<�9�i�#8{�Zƾ���=	IzY����:f@ )E�&�� ��t�� ���vZ��w��\$�̭�d!mW
��۠ː���&�G��|���@b�� n�>��a5�j�P����f��@!$L�ntݲ�$�%�}D��"������V�B[�D��d���w`�p�8������-��F�*tr�^�P�v�����l�������׮ (�V��8&%	���܏Lo�o�z[ �	4�������NIE�(:)�*e���hi����'
UԮxˣ6jiK˦f�Lj��Kf[J 10����C�4�"��<�47��bHn���p�88"���u���xPA�76���1 65i���2��G�	��g�=9W1�D��y8U���L�U��
�-!��A�7�*t��!� ER�}d�r\��җ�k��D�!=R��<�d��Fw�E�,�7���gi�e�_�Ӏ-�K��N��!@Zl6�Fs?��rl�[g�Bp�_!� ��g��bK�f�d�|�]��,����w�h�o,�<ѭ}�_�8���ã�W?D,��0����@t���)�"�v�H��2s$�w�:&��s�8l����tV��[�W������9e��X��:����!?	D�����-NK�:��@��Q���/�����lwo�4�ڹz��z�
60xo����fU�u~(Ig�m/�_ā�$�|��4[\9�-��r�u��X�-�0m&H�4K)�V>���J���ɖ�Ħ����e���29{W���KĎ'�a��7�pULWn��z�m�A.��,��m%D�;W�'���m�]����?f�o�M}�?n|��SX�;�� 3��޲�UM��~X���2��Q��=�,S���*�)�1�~[v���n¨�|�O.q��~��-5M%�h-th� �LH����b���-�(�U�]GZ@�a�����*1�i��|���u� 1x�Ʀ�tѕz����eg5`P��Df9>�W���!M�VXT���0�H��if����]��Ӿan��Rk��s����7vt��!��+a�?��R�ݹ@A�������������L�	�9�4[�po�`�����������I��,}�.6��V<�� ��1���c��xgm@
���:>a'\Ƨ�U87m�cɟ��z��䗣���Y�Ox��@E:�Ӆ� 딩��j����Х���o0���.jWZ/��O0�}��>_&DL��ե˨$��V'4Yj��q�h��Ǆ�/ޘX(��oP��+d���1kd�1��S����ɄX��/�\�;YXE�+���Z�z��w�����J�
����<w+C���h�3�JQ)����B�v𓢧��l5�5K���R��Rj�'"w���d���Ya�
i��J�֖ G��ځ�tH&����q��&����<��xqV��e�X1?ik�m�"�-:���Y����)�B��N6���|�$R�3$�G��gw� ���yŠ.(۱�u���ꃫ� sMb��$��>}�LG�$��$����GcQ�����s�!��{��(<�l%0!���p挮�Gm3Fk0B�xқ��`.�������sg?��Q��+Qn$�j.Y����4�����v���$�5o%��ȑ�i�*J��OȎ�%�]����!9�Xe�
땥�z��B\_��h���;o�sF\[�cλ`�jp�#�����' �V�1��O�w<}^ނ�����٥H�MV���= �1��͝��K�<чOO$����m���y9��5�z|�3"�t���"TgX+�D�VⓄ�!�sr����[����'B���� V�`ƀ70L�fO2�xk:4���/��`@���^��;L��̶��Y�f��x�����x �����Y�]������"y$��\<O?�(@Q�K~D��Me��q2?�l��!����Q�4��b��}�����O1�6]����rX@��U�Rv��Z?43��U����6ok8����̛
�-�Z��cS�
aX���X�SGJ��Ogժ����뙰�s%~�-�d�������y�,�Y���<�U:!p5w�I��6�4��&w?������f�a˼�}�d�J�����U�J������j�����"(�6���2�KH�����4MC;��e!�����?�D߈�`	��klE���=Hw��8�FT��~�BJ���l/+z���3װ��G�}�a�Y��j5�?�{X��-5�B~���*LY�~�����3Y3O�=�зWDņT��J�Y�Vq�t��F�Y�p���eAf�j���d`�"O�B��r52+���Tm����-|�v��=��eU/(�ϕEB�ͼdG\���!]�=!qh�̉ծ�H�o�� 8Y<|���@�53Z����/Iil���a�+b�kw�e}�W� .j�y��٥S�z�ܘ�z�k�w��UR��+�z�Y��[:<�j�pX�h�K���<��~*�H�;����%�G�� ��<�UO�t�������+����L��J����42���ݼ��6��fwLjxC�pxǣ<����Ø�X\<V�y�)���Z�Y�q2���P�J8%��3򹻝��`�/7M3��i賏y�4 �r[�o٘+ӥqc�`���n�d��n㿾Ϣ�B@���"PC��q���gţmZ3�j�yG����d������W^�|�����.�x(�����v1��������g��M��e�&]
��[{緍�����Z.�|W��kH(!�P[}���]L^�j,�q��������YyL_0����V�I�C�Q��R�N�p�8�8\Tŝ�m�����<��ĭ�Sa�m�/J�ΨT�/����*���ܨ� V	S���'7
4W)�Wy����}f�:���'
�Ȭ��� ��K>��O�J�d�)e�c�a�K��	���t�����Ӷ�uX�G�st\��5̶]�k�w����������<A.�oN��fȓ���g���(<�-�~D�b�RTM&Q� /���x�'�8�0���
'R�Ǚ�@�nTI� K~��J�p�DU�"#qan�N�f0����0o�e�,�{")B���4� ���L��
?@�,�.�^�V��^F���`�;�I���^k>�{����|��Ϩ�J#�P��J���<�*�m-�TU��u⊘)�h���<�i�m������ZunH�e�~t��}�8;��-��Z�#�[~�w���ץs�Ŝ�I�Sp����nvJ�=D9r�e��}�W�o�u�A-=�D����E��_��	�c�'	f��tr��r��d�D��#����;�E�b) 6�.�*K"�1D4�dڠ"eSp�6ar5g0^(L��R���q��7����*���4g�'7�h"5��l�����^Ez��{!����%;vsc�a������R>�>��吲e8�\ȝ4���Y�+�|��h~��OR�r�"�e����XO���Pc�3���qcJ"��.P�>�N�g)od��� 6�R�J��H�����ݽ��t�j��75�ԀA˭3�M^.�g3�)�`i��Z�X��(�O#T3��b��v5phjڀ"��w�',�u�]�TQq��y�1�e�-��z3H���ωem��缻�P��ri�6�Q-��s\U����8c,��u4^��\�Ի]c����G�ȳ���&DS��iE��Z���?m��l���\�:_o�{�[�wB.�XHW��Ϯ��k>���{ M~�/Ʒ4vR�m�͌�*�9Eg8~s�h��{|F2�%<��/V�'��b=ߊ�1?�^���uΐ��
b��1Z��+���օ�w�Id���br/�u�/�?�z������~�����*'�N��!ʞ(s䥮�|�����%�_����A-;,C���.hA��w����ܙ�1�;�l�g)=g�ڬsQ_#Y�Wt��tՠ�a)��.��8`�Oe�J�3��D�*� �!Ȫj{y2��?4$W��(��3�E�a�T���F�of�
��ri �r �T��돐���'��j�KF.
J}�f:�@C~8�9?e�6'Z�dtE,C(�`�@Z6��\|��]Z?�{�o�~���^'���Y�}[K S�(K���9�R�2Ur��Z����U��*���F�����}f���F��� wm�k�(3j�O8�ȑ^ZV�W8O�K�Xt2��}��V}���Y9T?h��K�[����8����S.������^��-���8�B<���?�l�D��S�+Ss%bGT=&p�a�Ȅo��|��H���L{���Z\LG1ϜQA-���b�V��s��^:c�C�-�k8!,�d�f�W�B�����:���;����P�e���-��2��s���vq��^����Μ�Ӳd9�YJ�d�
�M!Bq\¡�ۈ5���^8����g)����cb��DP� ��RH+w�=E�����a]JՈHo�]�@�!��m���j_��
W�j[S���}9���|�J�'W#w(���a)����i|YÁ����B�0�ޗ[Z.R�DsGiN��#.,k���m�}�a�ձnd�ڏ�������U�vб��zT_,>��B�bE=�v����Wt���e��ȶ; n����~�g<���q z�&f��"(��H��4��Ma�H�Ӎ�[�cO��?�Q[Lo���.3mN���
���X�st �5V��|�a8(�Uf�T�W�2�}�;��tck
8�jc�2��$G+������lNZӑu���5�LXCv�Y(�\F&���`����M�M��B;�]h�>g��(#ng$��������T[ �S-�ps���ϛ�ZUu͑v0s.�>�tI3KA���yݏ���l�n�?��bGcq`��b{Ud.��e� b/�I�ȥ�HR��=��6�l3�%m������f�T��E%���Y�ڵ��i�p�j�ܕI�BD��իm�\�w���3�5t#�*������;�(����[^�j!7R|�p!����-I�by>d�I�K��ڍs����t
	t�u��)�`�T����p�cF!��\�(P8ŋ��q�τ���Z��X͠�C߻�0e��2�?wC�|k�-���Q�ښx�)��@{���?�y|�?-cw�絢B`s�5_�Rr�U�2��Tq�0�p�~Yj����zТr�ǭ�Q�ㅠ:��*�o��a�_t��r�ξ�F�-�\�J&��5Wǯ5��K�?f`R��}vl�����[�*���3�(�
u�����F��=K���E�3l�޵6�����P�o�t��D��xR �+h�NaQ�1��+L&r��f�eˤh<�]�B�P�nZ�n����h������9�R�k�6*$�āN,I<�hJ[�aF�
�)qk ���4o�%�I���Ĕ3G>�^���d#�����:�=	���y��"/�P�-<yPp_��:s� ^Wa��,h�2��.L���̧#�n��y
�=>�&�Xr��(���L�2ja�rV�-(�a�0�m��f&�u��X��� �e^�3>h4c��!c�H���U����Ո��2�)t�.��pT�<�7lH��d�4-[�x�\v+�u܉8?�u��<O�K@��zu�s���}�~��χ0�3�R��_���7ꁢUmc�B�@O��|x]|e���d�2�Z����&{���O9j��~�E�7Ge�>�;{���D�o\L^g?]��K�Ҍ�>����P�.(�$����H��X��}� �lN�9C��u��T�˺��(�8���}� �۪ڇF���ў�2]�ǰt�晔�F/4\��@� ��W #��4���]$��2�²|�ܣd��l��k�۝Q0��P;& �L$R�5`����Q��*���^�+�B�; ���M�6k�%��o���%���wݰ����-�G�+�3y@�&�0:�y?k�H��-� }&������!ݤ8bK$�P;���c���`���d%���gx#Ⱥ�p�]8����@9��Df�����(�����M;PIV�ۡ��p�]�o7&7�@�0ͤM����}����]���O O�q2��`�������{M��Q_�/�,��7&���An�)�Us�U��ʎ�QZ!� ]�L�B�{'�˙�fA%�@� l�V*���s<��e���?ǒf�_CXW����ٜE��|��2&��rEa�8�ęq�m���P�.h��u��&��H�X[�*�(P����	��Ѽ<��D����J�]c���IL-D
�����-&�s�i'����Wl��3�f��d{]�H�0'��a��Q���˱ny±I �m�P	�ȥ2U���'ֲ�#�� �i��]~R�{�pIj�.�o4hx{{�(�A$qXQ���b����i�7s���$d�o�~�,'��'N@wٗ��Qb�z�x[(��B�n6���Ij�u�^�͌�j2w�A�d�q��&��_��~`i��ؕPgU'���z��6�+�֎�܌��-�k�j�\���;��dG�ٳdp�z:���H���۵�t�O)��9�Q�P���!Uf�$K	�S0s�n��ˬ`c�i5��%�L�`. Po����2���KR֦�|�}�W��6�J3�\�6PFE��{��`x�Pf�'{��I����	���셁�y2�YR�h�u۳�6yA�f'P����$�pn%w�l���` 9�xq^��_Q�ƪ!����'S-���㉦�����aj�v�9$�0/�a`Z�6٭ogC��X�ƻ��^�W��b�47�q� v��m*'65��zÉ�J�90Q������i},|� /������t�x Z;��WU��Е��JG"�����y�d�@b��ӽKwY��)���l�D���#���V�?�$A�
M/�-h�$K�ౣ��H!E�a�:��݀�I�~�ƔR^;\*N�y{���b�Y`�W���U��0�f��{��f7?к��D�n����v[���%˚�s�Ƚ�����7�7��I���'[���Z_H�������yY*b�6�Y�9�hS�lX�`J4˪�A�d/S�
]��G��t���ɀsHS�*x7���8~F� �+)ֳ��k[�pqs%I/�$��ݏ��|簊p��3r�1��ȗjy}�xt��"� ��=g�k�}*!X��R�F���vb	�����w�����[�D8�'�'�	'�,��%�r��(�5����<�Q�@��jjl߽s�������%v�D�e#a6!C���F���-�ҩ0�Q�3ch��܄Y:��p��UV��q�3�O��Q�=��(�Ƽ�Ckm܏��v��h(��V�i��B���goAS�I��,�&_<e5�8 )�êփ9��C̗�~��ܤ���������H�`2�7�K$��2�l`�Ī.������h�f�H%�%xy%0gl�u�͜�G��+9$�M�����QV�)ᷪ�,A�����Ĵ>����։޶���dl��C{�p;�cG-�a�H�?����^�1��v6A󅽒PYtX)%�����;�uV����鏄!�h�
���DӘ=Nu�3���u���5����4`�I���G%�����*kO?i���}�}"��N"C�>o^�1پ���^�p�i�u�\g�-q�G��J9�`�)�5�ڣ��u�E�c�F�I��m���L+�8f "T���������������ʕ�U�"�K��6x�����N����� ���6Aͤ![��_��������F*�`��O��2}���d��gRž=cA�Z]���J�>|�A<�O>2&b��\��ek�Vb	X�n�A4�����U�A��@ǵxp�a�Ҝ�8N������9�d�g�AK��F�8ũ|��K�d>���4�D�����QϗKY�������D����/�,��	�0�@���
�O�@?H<��swWĤOS�u���Iڂ��+X֣y?�0#���ј��v��H?���Y�,���w����k�8J�pe��������S���܈�*h����ώ����q�he�i_�t�p]k��
T��Q|i�.��k�q5qK�\}�)*Y�Q��lE�_<@��ɼ� ��.o�&;f��6�(%ȴ��B�v�,)��X��R�Wh'N�^�'�l t.j��Rc�>k�Sm}V�?��,�/'VVu�LARܹ�+f��!N��Cu;�n�b��(?�D�
�9��8A�;0u�����Wf7 ���5�����.���i�-�|{%�m�����U���:��%�t��U�),����8�+�)3d�X�lC��T0�V�����l Q�~���(��F��Nn�!��� �VB�p2��ez�8�������]uf"��r&7�|�A��9��'��^�>�]<1��]���ב4-X�z^|���E��c�{�x��إ�?*i����`��p�wW���`�����dN(7��2��s��~�A�:�ߣ�"��um.��6n"�_j4��)C���o���u<V먾�.��8)�H�jQKڪ�Y����y��"��<�P��	.fI���̎o�����Y$S��3��h�Sx�k��7l�'�B3�`x�T���X.�r^�ca�Y�a���z��� � ��{��㯑[����K´��gI� �o�y�*�l��`m����6�}Q.#�+�bV�OQ�
Ie!�� ,;{X�����S�} #|���x�L��ۍ�2�����v�qf�+n���g^�Ƒ��I{���b�=���-��z��#�}�?�i��;�E^�/�פu�^o�z�N+���2Ҧ#�2���dXd��������.��n42��]6�+�7�6��n�]{�}"*����g�2a�%^
߅ƨ�����	�t�y� W
�9�v��|����t��5����+:>/LU�3����wL�a�`������2�U��>ܑ���Q4�A�l�D�a�+�ߣP0u�D��&a#�Hnf�]�F�qb����΂�#���H�����C���\?B�.����ǒ�0dz�!q�ʙ�N��
&B�֋���jV<�'�K
r}^U]�!1B�RU%S��`�����;{[�<A�Q]r�%,����[�k�g�8�Vi����m]W�nD�-:�@��)��X�	)�e�?E��l�;��ŉ
]oRZ$pt�.�
�r0����H��A:�^BnN�<.d*|w�9s����d�`�@��^m}6μ5�X�)S��V�/2/�+|֑h��Y��4;�kr�6�ɳ��-�ó��q1��2՚�c �A�݊z�S�Б,Y�{�k�cp��籲R�:�\�� �g����K�e(4�f��`�o����_J��j�H�%�^6'>�8I�!�0w�u��{��j�Fx�SO5��
/��(7̝F�& �&���y���Bx��T�(AJZgZh� ���!{G�8B�D$�m���úR���Z�r�$������󽛨�9;.h��2]2�c}dGMk�.���+���\�mJ�E H�r��6��s'��,�9�7�~)'��,NM3?���/�8���yQ9�(5�Ͱ��?	�J<)H]��㧡��2�`���$6y?.2kȗ���v����������P�r�(;@8���u�K�j����n���f���7�t.]<\���20n�gR�羘���ŻLt`�	��d�q�>�f�W�;"���#*���uW���z3��r�Q�X�7�mu�B�J�SMa	��ܹ>Q�d�t-&�_qpF�F�gn63���$�*of�B���ѶXH�^�(��(��Q(!��i���8� ���B��K�M�w�u�w	���ǫ�c��=���c<��ېjP}���K(�pc �� ���ں���m��Hw=:[�	��yA�l�2񋕰�,8ԑn*^؏��-,���4f���*�UQ�]�@�KH�e��� 9���+*�:�
&�`�zF����M:ܷ�	(�.�9)o �BC�ղ�l��"����I
�����\�	QTB�� ��?�-�Q��Q���kt��E���D�
�m-}��gs[���8	�6$��
~�֚�z�f?%-��2l������I)�-'R��k���	@<e��#���%�����b�R��-&���*�	���r߽�$��t ��r�l7�sE4�cp\TB}.0�������.�bMjܢ�L��܌?�P����5Z�_�Ԧjn��q�c�Q��@�I�7��/�m���^7�-�'�g���o�G����0��v�7q�eA���ü|�i\��,T� �d����� 5���G�'�6h�r�ȍ�Ae>C^E��^[�E�ꈐ''�F(����}$����ѫ�:0G���P%%��2,�9��W�I�dB��o��]�Lk9'�.jBK�}h�t��u�A(�xO�
^m?J@z�q�Ł}R���8��M�5�y�P~�%�pR�����\�Ǳ
f��;�.���,d��{�O/ 4It��6[ gC�g�W���j˭��)�Wz����"չX��l��3�w�[:h2�½+e@����7U���7�����_�I��۩[�N�9Rrk�J�j)՚���М�>y���YM����a���k?����WK�J�Ez���~I�/"Lvt�����W��"�a5	8
M�#sfS��ƆnN�vxHfKL������}�4�.�c�.��5e�?R��3/��H��|V��p�l��e�:�k�ru��~��u�x;�J��C�5`$�f�`��|4�D����m!͍� iK�3����k�Fv
w.���9��_�⻠	�����D�,C�j�(sX�,~"2Py�j���9��,� z��w(�*�R�T�st_�[q�������+���I�eD�G"^г.R��H��r�28�|İy
������T��{B G�����Ϊ���A~��p��;����d y<$
T�H���&,�\�c�F��*����We�z{RCVL
h(�r�WX�Ʌ�:��B��u@�T�5:���ps�B��׸�3�@�E�_C�@׀ ;�4����_'�vi}���ؗ�kU���Z�[�c�G�В�"�>��10�v�5uӫ��5���)����@��	�G���[_�N������� �%���v���h��o�Z������ )�􊀕P!�Q���Լ�����ŔB=e��/,��@q�T�}����z꓆F��q&�<d��K^Tk+H���}�TFn�&N���
���Az�m���.OΙ.F��7���2�ö3��#ěrtW)ǝڪ�\#�!L�׃m�X�(����bu8�)�.1jg���!��&%6D*_��V��hA��U�*�]��8���+N��sO-O?+�ɢ�ׇ���ɢ¬Wnb@�}�n���$�M�ǭ< �Ɋ�YJ����vR3*�n��,(�8'��||4	��p��X9�s';&���?���Q�A�G�}���\�gr�]t5���c: ���|a�4��H򹏱!\_��kH�D����ay1k�:�50���'�0B�Gؗ��Rݠ�M�F%��t	l���=19�&|��SΊ�?���Y+U,)E3�t��T�t�*�!��2fEƆ�N�.�y�2 F�c�ZRy�����>mZ��/ՙ#��u��jP��`D��AT�m񚏺�P��"G~O5u����G�q-���+}�~�>hkg6:�ueZ�WX�Y.E#��èN|�~@T�%�
U���&����>�q°�p��a)�8C��h��K�����u�]ބ�d�'�L��M8�Q�{_�`'ץ�0��F2.��崌-'T�$�邱�'Q�_��4Fn�q5�r���/��qK�t��*FƬs�v�6�- -�r_{?r�S,�t�l��]�����=hkw�w�Bx֝a\���FS:$�>�AW�9�_G0�pp(��5���|�!�}�9r���͢FT�?s�x������
�YX�׆���d��*��z�KFf�+�Mm�BA�m`Q�<�ǫq��81����r%�����
%\�.�˸��\�H+Tх�� ��#C�@>&���NPbg��Î�i��j����m7lŴ3�����ҏhy�Y��nڑ!1�Wj�w%V:�[�8��~ɾF�� �ݱ��*�o"~�1r4�-L}l��L�Q��#�+��\3�����As-;&)��+�<n��B�3����Hݒ�|׾s6^����j��D�:*.1x��PW|��"�� g�����M�|�A�M#��6$�*�|?SQgҷ4�Y�M5�kw��~��t���Hd֧m�h2i�Y#y��uU
�W�s6�`PS��]u���hny�L�����6e�X��̈�M�0�dXw�oQ�U0sK
����� �zm���0yA3?(1���oT��J�-��i4���E�q�X���g�z�#�|�����b��B���%�-"T�dzN�c0���˻� |0B�>��#}d�}$����G���G���m��ox� ��MI��r@��\'����/���1}cD�L��~��b��WD� �,�ӈ����\���	�кG�ͷ9�\pe(L�!����Ƶ%��S[<3�.���:7p^�adqb{����'��ӫ-��(YU��E����F��+&���i����/+��I-�o=�`��Oٖ,��zM����Ku�?�@��O��<��`y��87�ujC
�=�)���DI��<@5#�7���c���SL�#���D�j���h���j������y��*(|Ƭ��%u�rLi����YJ���N��oǒ~ (��T�B�⌷���y�h�.��䋛i��}6
e��~��Y�$�_AJ��%X������;.�[c:�s�I��s�p�c�:�d�a�wu���d�&K4Y��9��F+� ��/xm�S�0C����:������Q>?�d���檨�ݲ�����-(C4=WZ�K��]QA����Ԉ�Y��쵴I္m�>Y�_a�-��.d��6L)d�϶qa��:��.r�څ�c���z�^䗀-D]����h;`Z��!�*t_Z(~��͕&�:,V�'����a %g���F	(���ʶ�R
�ڗ�
U�0}�M�@�G�MǗ��iw����G�V��~H턄��[t�y}I�a�9Q@.v�g��;o���ɠ�h�|;�8ۧ�.6B/W�P}yc0o-���"����vpJ>s=��Z2m!��߅�"lV'ë|;�0&!�b��[Z���۫�-�u�Cǎae	����>:d᬴��d܆e��@FPJ�>p�T�Q/�gmA��/��K�v��K�??�uW�f�7�O�,Kt�(Կ��l���x�hL=��8vx��l#��e�_m�~�
���	����UnUnXV�h�zo�$�ހ��?�FzI݈�h�����DXJ�/�������v/�Q���� �3�����z�L�i|�9�7UqK��)�y�Jui�9H3(3��W���Qjzg{�;�0 �`��4�*���WQ$,A���2Iۅ졈�� ��fKL�����RMQ�-Ȋ�'���a��.��S�,KȋGt�z�k�9Dzr,>�9�F�������"p�E1IT�#V�F���-��a �AW�	ݲ����p$�P���� Ҟ���@��g��N �:�LU��Y+�k�ad��g'�7��6�g],{�s�fHЙ=!׽S��I�/N������c*�_0.�����?��l��-�0��H�V��GP�jC,��zS�8��l�Yu�
�UY*��^����'���3Ҙ�(섃#J
�Ɨ>{�jД���ȁ�/��2&oȧ�����j�P��_���
�"����/��9�.��Q���S�,�V�`�(`�g��Jg��it�^�&���d5NT������r��3�ֈL�q{p�!�f=ᯡ)V���S'�]�Ŧ_@`��ZM��tfC�;N�ϋL[2t��U�_3t"�|��<_����J��� 2}��<��)�T�%�"$�1}�R֖��bX��b$��)�Bx�бfQ���Z����(S�d���F��۰�76��x���UFrR7 
�؝+���HV'K�FS"[�{�"���ݲvw�0<0������;�*>Ý�� k�2����aݏ��7�$5��3�6=�Ē,`��B��Ȉ�~������t��!&-wip'����}����\��m�!9��U��
�"�7wk�ah&�H�.��5j�X��9�G2��V;�n��7�V��u,.�����]�]��m�|�@b�n$Uŝ)����hK�s#��=�8أ{��?)�ɶk6�'�-3��o�G.�������e{.O�aq�;	�[~�J��� Q��J���n;i�qI��O��ִP�`�XbOVg4;����2��|�x*��ӑqk��	�WYc�/�@�%r��j��i,�5%�L	G�| H��<)����H��ق"�� �Œgl�\�g��N�駂B�Qdq{����v�8���s��cK�k�C�Y�	Y�~�� �:�3���r8 ��k?'*a�B�� ��5^{����DY�lm����wE� +�牰PV	�LFMj�:�����}�1�Ȱ��V�i�Ed�^�3Rb�7_��0<Gu׵���}��|$J���kV�
��s�ʱ:��-� �ܵ�"pӐ�:�[!��(_��&�ڱ�ʅ�3���p��[x��땒^���q���b`�V�\sӽ�,���@A�6*�b�p�B�����ߓ�JJLj:ztDgI6��t\������<�b\�;�L�Rz
��"�.�)=��p9rN�p���;�]i{�^
�����B�̷���9�fF�I9�������Z��g��-L���H��cx�cn��jC����T^8���v�U��bl���}m�O���(��`E���`,�ksu����v���z�'���|����*��Ra�jF�e�e�,�d�7&�4��վ��r���p
l���rĊ��T��˒(���6ID��/�r�P�"���/b��	y�'�-q���O3�ˢ0�����Z�ЏʍR������{5L$�M�Y�Ɏm1���DK��P~d��0c��o&;����5z�\�Ijhr[���ʱu�4𑭷�)9k\v�ߌ�BL�_��3��f��rP��v\��I����A'~��Fp��g��� ���#f��b��"��!��%��"i���h��<�-/(�����^K,�\g=;����t�O��8���w`o���JP�X&.eiD�զ�ԣ*i<�;���QJ ��G"��t��Y���8]�W��G�Q˳;��``��J
V�^T�i��*n �Y�/��>���lΦM='�e��_*������9O�6�cq:�����n��������;S�;��$��Q&���d網L6 ���)n��J;���߁�WY(�p�4���q�)��i���8�#7R%�	T�Fߛru�9�����r �@.uD6���w:j7�']h@���r�P�֗�O�l�V+�����m<�U����0���6��O���6U�d��x �h��s}�<���g6���T:d�oE���ER�Xi14ѝ�k���$aJ����_�N!�������!�.��J4w�AA��M,���'�a	T	����-n�>�k����XBf:�x�v�A�� �l)���n �kӬ=M��������UߘX��3�lָj���Ky3f+��v%�#��"Z݋ZKp��ͣ �|�R��;�e��H�(a��iL1���pBhn��i�/Z<�(�S�[:iqD���i����ە����O��QAz��GZ����;���e8NlѶA��^<j�9�;~��(��<��`�.���ɑ≡xFx��W�em�����zIE�6���A��� ��<�
^�o��u��UF7B�-/�H� ew�R6@�P��H=�a�@qύ�S`���6�����i0fg #��X�Lz��[��ɵ����d��Ȋ8����<=䪰;�������^Z�V�0y;�b��B,'�0K�y�j!�`e"n�h,ܬcpeV6�Z��q*}�t�5�{'�#8�V�.`��47�����(��K�=����ߵ@���7��	I�tٔ:�v�'6!�ׁ���N��^:+mS~����C�����Ʃ�v���x@|�p�䲗2���R�����d�֙A\�@k<��vV��
��]P!=Ɓ���c�
���u7h��4j��
o_Pڞ�IpQ��S\CY��s��� ���A��F���5
���s$��ȶ��\eL���[w�����m
2.�W.N+e���_�~�8=V���7�*Y4j�����eP��lAtҸ���ȩ-MKÆnKHq���i�@������i������v�G�˩��w3/1�<�⣗�F���T���N����TO���wU.���bɉ�¡���d��&	rX{������Q��C7�����,K�yt��]�)�K#�4�CǟAu���I��O�MY���*�"LԢ
P\���
"A�}�t����\M��{Ϳ϶�H`��"�_�bF���U0| u3Ǆ9ݝ8����/-L�z8���bo��&{�Uxӎ@�st��e�᪷EL[�4(���<�r� �9?[��Ȅ���1p���-!Uj����&����� �-AՒ�ML����%�6.�^�)G	���V���LϪ8KE��A��ud����?��t�73=/�z�:��6�&�d�*)+�Am�ϥ�!�s�r�瞱8=�`.�:��q�Q�y�jgdH��g�ܞ�=<-��ݫ�S�uGsX�I����㚓+"��ˍz��!]º�M��&SϬ�@�m@��H��a P^J�Xl��
����#)PǄ�V���my�;�ω�>B`a��`�
Q{��.E�����r����}��g�f�#�D�\16ϵ�yE���u.ۺ��[��Dt4!;�O~[�uP�gČv��s�d�f�l���:?���D�;��O��4A0�������3:���AVK��M��|$��uy��7Wu/M���6w���U�j͚�<C�y.�����5�!d�L2htWC<T2�T.�n77��1a�6Qs6Ŋ��+0!�^�uZ�;�m�>�&2"�n3}�\E�����b����ʌK��N�g�]��Π��s�G'������!�,q�x�[f������]9��YݚZ"�|�W�<�hA�M
1A����8^��#����ӱ�f���d��5�2�� k����Q��T��;���?�_NA5D�8��`^���$Κ����at�!~�`�Ԟ�x�	�������߅�T�&�c)p��z1���G�Y�i�����r���D���_������y.�xC��q��|m���轟P��)�*{�Y���'�x ٝNU<���8ho�J<�+V2�d���^fb��F��-j`>�7X	ה��������Ww�-���?��=��T��Μ��#v�!~v�C��l�L�^0�1��h��BŞ�6��a��)�+��d�
�k��\C�M�u��3T����	���"�����cm�<S -}��:������2�s���>�\ye2L ���֤"�~鴣ѵl�{x/����\�J��?P��� �R;�R
���s�>o���e�{����(�\k�{|$e���	��^q�KB��M�%I�tTP�G�9)G��c�C��\|`���]�2W����DZ8�kd�S[2��i�K':�IF�RiB��tA� c~nei��i�F���1gV��$?oz���i�I���=���A�F!R#Ƣ+�6�Wu.����Ɋ��fٴ�p�a��2����J��P� ޿�<D��1�ꈃ�4�n���[���.�b���Ю������z�	LD�y�;��[/�ɧo�i����R���&��(F$�vq�꽱��"]
x�`�ɃS���H"@��e;DI�R50<��LA ܲ��*�Y�����% ���lC���`C �(O�%P�?r�,��������8��� 4���#,��<��s������a�(.�IP	����kJc)X���~C���k�2Ͱh!ȲHz'_�U�.>���Nw����݆�x������ �n��bLG���c�_�W�:�@�ה�R4y��?�+�?���z�Iq6�8|?�Iq���2V�*���IO\Q�� q�n{�������nJڬg��>�����[o��\�S#����A6�WR�^�O��bG+�tsXP�,�@����cI��U�V�pL�YMqD��}ϠzZ�7�Yz�o5��= �a8���*.�H�+��q��|8IX��R֑B�ΫJ8y�V�!����|6� :��3Q���kSD�H.)� �J<e��nH�����y~ؖ��o ���g3��_�9�0��nc���vj�oE�-[w���ǁ��P�b�F�HYG��	Y5�y��Y�Q��9�ͮTB7�c-:��#�"m��4lHٰ�T͛Cfm��b�g�
�9u�+��c�A�ހ3[�	;l �<ղ�R�W��p�r�և�D�v�U���7�g�ZN
�a�i1$��{ܧ*� ñ�J�nٻ7��� �4'�����d��l0��r�@��mx�_/M~B} ��
Yzf�p��I9�%iVЫHО�v�jD������Z�Hm�<�EМ���_�I伭�2���pR�*�W6�FT-�17ی`�$ԾC���\<^���>-k��Q��x�ĝׇ-Bc�e��&t������n1q^����J�1n%k	V�/�*����w!�H��ͦs��1�*s����D_�N���.� ��J"X��?���\� ���9�U��X-	5>�/�Z����y#c���Q-mN_����ͫ�)� V�r,9T)�U5��+zs��n;މ�u�?j`S���G�
�'&EnDhO���������k�HG��;3{%��E��B���_�����w;���7��O*���"�y�+H?2�44T�����=��
Ih�{q�r{/���@�il4�o��p#{����gu�rz�;�Y��
"�,ZB�jQL�j��؉Z V=`0�F�C2�^�< �������ʋ�Ȝ�#�pm������w�w�s!*sh�;E����-17�[�/��pYM��y�m����%o��|�Z��ZGr܀2k�����/ƈN�d  n����E���FF0F��y;��/�=���d����� �ҙi^:	vЌ$��,����#r�2�f�3���>�����RV"�_M�H�T ?�֣�xiheU�\D�숈3(a����.7���1�!�ܑc���?�!�'\ݢꠅj�FO�(��F�v껲�E;D��]�G�,�Tf/���I��b��*��QO<f�MB�|�6�O��KVB�H���� ��Υ2�j����ꔭE�bc3G)8Cß�Б��wh�o�9���n�iR�٘��fAI5�+kD�a�{��6㹅��3��I^�N�~�6����#�y �-B�,��2_��̮�'��#U`�N����F'?�?x�\��>soZ?�	]��}��i���Ur��e�r�7~�סU�8�`����_�x�.��M���9�V�� ��(��)��죐�{���Fx��e�,7�*��n�1F�2�1^������½N���?�oH�;53�C������1�"��_�̝���-K4��,?���^���ze�s(*�I��֤-t��������f!�a���8���$�ztI�	1�~��$!��W-�g2�;R?0Rє�$)���NKp��حR˛.��N9��#ފ���oZ��t몥�q����4��d5���xj�:Tz�B�'��{7�����RC��
�]`OAԳ��[����\�=�N8�	W�����̶��td���i�i��;�&yb������R*A��8������v��[�X]竹�	����t.uy���v�� F+���R{�F!Y1���'P����Y�w�6JI#�-d`��ԯ5m��6��'(ůսͰ����u�A+W��+Bgwfz����}`pR��(�6���[��JW���� ?ih��k��q�<@N��뵂�m�sQ�'ފ%��+H�!QT�/�ӳ�&�����X��&�p�2�1ts�լ�(�e��sX;�r�e���ϋ�\��"$.Vҍ���&WZ���2a;��5��7)m�$�� �1>�2~��x��*l���Dq��x�����1�����LX��	�(h�1OU���^��u�I�c�����s����#��LQv���Z��x�� ��_��[1#ēfh�N��2P���U�5v����Ɗ�9��/�+S,W}�����Y�&���ė�"\.�<�/x�},�fr|�		3l"b&>��.ϋ1�U;��!e[܏�$`Ľn k=郿f;�,�)g�����X����!��߽��r����5g}X�Z���LI��xsy���h�3�܈�r}���fF�{k	���i�:Qn,w�=G��4j��$�U7?��������+
A��3�����5թ��ǽV�˗��l��nn����,�I��iSF�a���D���r_�&F���cY���[�88�++�P��/��a��?@�ä�)v��u	'��@�۵U13-��N��\�MX��Vƕ�1�v=>�nD��3�U �86����,=�y�\�HE��f��J���_�K��]�O{�$�ƪ�ɲ.r�+�09��ol�:"Ơ��}\ka��zޣO��T``hC�Y���b/�!=E\����
v��{m�����]j��TNl)���]$�3yU4�����s�ϫd���kl �q�`"N��E�洅O��l\�`1��8o�=�U .��G�P���������L��I��n��70�ȓ���%*�8G�d=KiV�xw���ހ|-'CT��*?��g���)
�G���P��ǡ�< �ؕ4��lX��F�d`,�Tˌ���Z�)6"r+���a\U��±�Te1'%��i���r�rblh_\�j+�]�����Ca-Vf��_'//0�%�`WWs�Ƶ���^c�'w1�ާ"+��]�Ŵ;���B�+����#�#I��g���&Pe_���c�z����ъK��@��K��$��Y���1�e��˔�g�o�)݂ ��5c��1s�[Ty��#�w)��ޭz��{�Y�v�6����{|5K��{M�2MЀЬ�-�˹��}������
�����bI���&o����"��SA��kp뇉�m�(�O�ON求�3,}�@�#�	�*"� �Tއ������P�n~����;/r��ό\��H�����E���Y��_�8&���80�OTΧ�Qw0/3vl�Y*,�1��Dh�`r�0Ɔ�U;?=��ӗ%�^�U���Qey)��s�DEŏ����f��Ux�~�1������e���5w��X*��Zq7&V^�
TÓ:��G��H���ł��h����)��^g�Q��7����Yk{��!�s�f�$ ���A��_�!�/u����>Y�)�˛�����*��J�>N�M���SƋ����y�pPPݺO��dɒV�����I�f!`�F�d>�~�uP�yg&��K��B� 45����C�зi^��O�{4~wƘ�V1z�ƶ�P�j^ɵ�4�<��Ӳ�S,�����!#��Cg������i�K�cnZ�#�S]o���Oֻ��cx	}-��k�Io�Y?���i�X9J`��G� �9UϿJ��v��CW+�yh�M���2޲��`�w]R;�?z���տ���#�d������]x�ʗ�R�R�ђ>1�S��I\8�|��_�L�L���Rʳ��|�5_#|��2`K�b���m����I�*��S�Օ�s�������Fo˒;'��չE)����NR���_3��&������!�bYe��|�e"�;��xL��2��Ɏ6��sV�����EI��n!&�*J}�1�,2��4��6%W[%֑,�LX4�z�#SZW���iEq��p�3醇���ȯ�}`��fѸІ]op����nH��D� ~k��1?*^���P�gIz g�`�
q���N�z�3�(C���zۈ���4�x��l�v�Gې�k}�1N,&ST�9L�Vk���{g���}i�W�8����$l�K��¦qv24KM�>˂��EMB����ԟ��9ap��:�Y�@��ju����DM�������̜w.��l������c0����O�V�|��=����G��*JY��\�_Cn�ԧ���2�baĐק��{�x�&ᐁr`tV���еe~T���$�S	ށ��ꋲFK6ˠH~���U�63SSq�R���_)�K�#�竼�d����c�Q�.RA���UCGc��4H�!"�A��+���}����Gb`����~]��ŏU�U�F�I7,�by�:n]/����b�@˚�����Sӽllʍ4Kp����b��ه��[jdگ\�^#�U����������,�<,��u�qj^ H��`a@CF�ޱ���R3۔#�M� ��҅s�ӛ���A�p]��"�3�������nqVUY:n��#��:�o�Ẽx|�^�<}��J��H�p�H �>���:��<��t�x�Y-Ę�n��}���S���Q�2��fƸ�� #1��%��9!�i��.Lo9�6�F������f
	e��ş�#��n 1��_}�W,�sW����MD�3��*:�G�s��R[t�זZ��;ۑ��X��jl�Bٞ|8�ڷ�Ər�dR,U�
��%Y�6><i���S	ՠ������#Y��bN��!$�:}�	��6�8�Y�	u��^�Qm��Y*%N�k"�Lob�	�v��M8�놨$�XI�N�/H�����b������]�
�V�G?c}��W#73C ��HF?r�x��|Qץ�!oK��]���dd,8��n�%w�����}UG���wk�*�M��:4�r��2���K�85q���B{K�3�q�V(Ȫ�ҚU�M�����B�{@��-v��8%�����">�JS����ul�Ԟ�.�!%<�5�x�t�w��Ǹ���Y,~V�Z;I�8e=W%1?L͈�Q������� K�zߺ2��T����C��ذ�6��w<<d$,A����f��p #]X�ݮ��`T�mh-�zFfR"�e��|��S��ka,?e`����[#Ss�F�� �Ǳ����1Dy���!
ר9���+��):��|b�����ep�!r;�	(ì�]pUt�D�rEʻ#�`���K��la���P��?4ue�.�_"r��<B}-i��.��k�(/m������xx��RqdFp�3�L���e�:)�*��5s�'	?{��9Ρn��oۨ�
V<��I|�ݨ֊��#�ݢW˾��W��_ʈ� ��e���\H!V��DL�L�] ��5a�٘:P���0��vP;��Yje���i�X�*�٤]M���{�&ܖ������.m��5�;���D�t�E��*��������WH[�H�/��]z�85�6D$z�?�*�:l\*��D�f����A�@�ru{�ѳ�e�Z;��1��<�غ�<?�F@j�șYi��t���A��#�Y1=��m�����bSi�hY!�_g��q�Cѩ�'�7#��w|p���HA=�ȶ�ʢȘt1�`o�Dmƃ;��`P"��o*�4�W e�L�_��`=��~H[s�������DE���(Q@�@Ϋ9�Np�^`��rX~>��DQ܌�6�����(��êsB���|^F3%fj~� �~u���Tc��]�i��#�u�گ.�*� ��p�l��3bV�̃��E�P$�]
�F]���%���w��=n�0-�_��i{G�]�((:.��'�[���_l�3�Xʩf�Z��b�i<����R�5�b0�=l[6�R��(������7�^�G�HX"re��W�d�]B09�W�����*6/��Y�����Mvب��D$ �.��U�"�C�E.�J�wOO2�W��MCk���Ĝ-���w.�~�%
�X��\�p�$ڶ3��tO����*���$T<Q��O�M�Z+��4�boc]��-/_\�RB�v�_a�;��V����D�Y��7��������4�"Y~���������!�H%d�:�iժMr��?ǵ�,j!K$�{P�H�$j�	,�u���r�A!�7i���.}�~�0uލ�C�	&� I�m���vd;��z�D�b	l����cS����JlW�uLlmA�F���]�����'�k��d��)��������v��F�'I@3ݫ6vA��\�`X�X�B�$�Wh&K�~��5}�0�S\�{��=�KW���XW�/����n��F-�#�}�T�n�a?i�<"��Q��1�+E�|�OXD{`Zݜ�j��<�@������af�1�w��)��r8m��%��-�S?H{�G� x������l����zҨF�k�ҝz�
%&�:��E7OХ#/������P�Q���J�o$�mw�aHB2��p�J��V(�P�!�1����Or�:��MMGU����ߠ�XԘ �`�T�9�Vف��}��ш:c�
���q�4��Y�W�ۂ��;}^�e!B�3^�3��KN�H-���1y��S��_r&b�-�>.�f��S�����u~\�����h�w>�Ҷk��v�Ê��w�9u6	��Ff�uj߈��*�����5�Q����^��8z�|u3��s��Y�cS�nC�g��>�<<ط8��_��<��5lU�0a��� �R��f'?�а ܴ�������w,_c/�i*Sc���:U�<���U&jKǢ	\@�c�%`2��K��_��mJjִ�XkF��z%~���ˀ�E��O:����^�u����������?��9G��#[���v�f[n�}f�r�d����o��#�*�./B*�<'3>�!:ڍ�Ye������ ���U����d�!n�Y��`t��71�7�f��}GDJo�ϱpﹺ!�*/��eK�Χ>4��ôLbٚU.�A&К8��PlX,޴&�%ﶞ�8n#"��Ο�|M������Z�n��R�G���<IF���GI�+��Zl�zc��a�
�(0�d��"yx�����؃�E�r������K2��(䆱��}������Qќ�3�\��[bZ�2���]I6^�^@�"x%��v�ƻ�ߗA�G�cg�{� �,8`֟��\}�]�,,d��kC���8`����j��؊N6��ؓ��=�u�%2%�b;~~��Č��l�+?�Ss��~~gw5�Q_��8�DD:[�m�Nڸ����]�O.�j��8O�b�P݂4�$��!��"�^�Ay�i�c�5v��RenԜ#��=c�o%{�ؽ�>���R��Y�L-(2�{�/B����hNDPaPw�	���ϋ�������N��E�Ţ_o?�˸l�D� #�Yަ�^�VdgC��MLP7⁣���3�y��>G����ib&�p�s��yz��ɮ5 ڄW7&��v=nH�)/�m�O"�����ۊ��#S�2h��<�LZ�x�}�Yo,���U���k���Y4No}V"Q¸�������P'%f[�
�s~�1!7�w�T4�hC͌}�g�[4�<�a�?+��k���~�כ-��*3��U�o����fS؀7�̼������T*am�I���]9���UX���a��q�f��p�Ov���Ǥ�$SSӴ��d�|�^S�Jq��h�=�e���Gs�e3u�]���?w��C:X��jb���Zo>�/w��O��F�I�V�pa�� ;W��?�� ��c��F��=�/�EX���|C�sVu�z�U����F�+�XD�瓨!v��_�JU�Dx����)�+��	.�Q��6,E���&�'��1V�Z�!�����A���7�J���ۯ��5�	[�Q=kɄe��L��s貧f���لG�CK �Xy>�A�����]�Қr��loz���e����"Eh}������*A��i�NMp��H��I��~z�HnN��/��٤a�)�(ވ7?���@�H�u�>ʔ�^O�-�C�`6��Z�_�G�6"t��O]��SnA�#����N��=Za%�����KW�Bk��2���s�O���Q���4�$���D�����L�������A�R/N��	[��8^Z�u�E+r�1�� �8=:ߛ��u��8�ʫ�Vl+��e�bBJKqC���	��,�j-�;Rq-�)\��ׄ�N*���DcD���_�
��K��ɟ)���N��_.����٬o�;�f�#1)��z�p:���J�� ��9�^�ԫ҅��LN0�GB�2�����
̩yk	�d��%h�;��p���S&C �-��y��׎������;cb��Ԉq����55vO�L�JW`8hԵ��P<��*AqO/�\�fPR%���,��v?�봷#�����f�F����0GMx����Ϭ%��ԕy(�>d8M^��k@£�?�-a>N��߰����D���@]�F��kc�����{8E�ġ�v��*X���Rz��2 d-�)�NC�)7��떢���a����������\ŝ����.U��O�2�[���*�K�3�g��'=�x�0���գXoʹvM_i���p��vє0f��l9G�je�ݑdw���4i�
�s�����GI��?]�QPa >L��׻�B^��.����s.UR�5l�V�Cǐ7#w��S;���&ߓ��xג�Bb�ހ'��"�0tf����������|�d]����K�@\@х8��2�)��L��ЌZ�ۯ���|�Ջ2��o%|��A썪�(OZ��]$�q���d�Ta�&���+ ���}7��q:/g$���T��Y�h���LmkF�E��m�:����a)�L8�`^ka�Б1!���
�ԛ��c�E�dy���J����>��uuG�QI�Eط����
j�`�-�����ܧ�<C��cd�p}��6$;
s�|�&3�&F���6��V�zS�]-Q��΢0 �+�mΪ�j4���F� _6B��d� �˒pM�s,�f#�-�����t���o�?Th�PV�ų]h��u�͟�Ԃ��.5�)|8�~n�բEl��ǔ����C�mtw�g����Zgô��ԉ�OK)�L�	�R}��Y|yb�j�WP{���>�q��y9�8�i�>	s��	Ϗ˰�X��u�)��3�e0�%����X,���c��*�I1�h���G*z�T��oJ(�Hq��
 �&�7���S���Sd�_����aQ��T%!fx�ؖw+�!f(��:g˿'w;�ä�YU@P�q�@����N�Ͱ{�t<.��E��$���޻��y��Jo��|��3�o�ւI���>���;�}��}~,gHɀ:h@��<%	[�V��A���2���(�!:���������ۀM���b�^lؼ�"UmԽϪ�9ԫ�Ȇ9��F�E��k��{�o�zq��4�,ӌ*�q%R�#T/���׹y��#�﬏�bj�h_�8s���0���*��x_�:��>���gno� �aTue�cM,�v�Gcr�`D� 3��� ���bT�q��a�x�"M��V�G~��-�ي��OWk���d�H�8���B�*��t��ڭ���c4��T[5�R��f��T�˳Kz�y�}�'%���"�Q�j�`�i=�!t���(��d�XC�=Ai^b!�T�����(7���EԿr~�|}0��#Xc��'�TH���`ى�	\�7�)�k���tD��
*����f�%߮�����.P�N?�5�k����?dhM7/�$�����_U83`V�9�U��5�!��� �z�o���d��Ūo�1K5�O�7�*ux�w�����G�3^�l�D\����;S�؝n���V�Y�B)n?[W�0v�%*�,3�A}*��+%V�i�!�R�<D��v�z�@���τ�4@���ۣsD -�������}ns������N����we(��l|���#�չ:=J1��^�Q"s� 􉷶���M���o	���!?��9�Ck�d�c�����_���P0l&�7�z� A��������]K��$wܤ	�'���F���a\��}4},pd�V�:��!n�\|�[���O��`���t�al����҉? k�a�?^��e��'�A�"�l-�`6�]}�'rv8��xx��͵2aAo�� �(C�O1�n�ȥ���.�r��%�i-�F�U��c����3q��gF��Vo���u]�r�h��m8xLH�^4������C�φ�y��/&����'L��p��)3C��7����?bl|b.�t$=�Ŕ�p�#����Ѳ���� ���	yU����~���/2$_X�LY�c�By���T�&a�;��S�� ��Ȑ�{c�H�ʹA��lH��VN��N�FFEϳsS�/?3�d�w�P����������`�����"���ǔp4#�^����n\1<y�05wmhB+�o�X����Hf�dk�>���ހt�s��K�ńym�U��s�ʏX�rfO��q��9�2Y�ɦ�[��X8!�۷ĥ��_6�vl�",D��
A6s��=�v����
�lrs�ͫXOM�R���я�+$A�q����	?w=�ߏ;^D�0Э�d@��8w�a�ܞ�T�JJ��[+?S�a|c��}������1-N��X�6�q��q�+���jop~�Ũ���,a[�zyj��,�eM����5�#>�����������|P�}�3G��=�ev
d3G���EO�'���xjI�"���]}��W���7,�I�2�,ƀ�F[�#�[Qv'�%;�R�zsj���;��=S?2�}� ���K�Uh:Y�s��I�xx�3�N}�D��*�e���6V,���sd>���r@K����à(c��7�P(/�)�*��eA���e��JR��������9�S#����ZZ����%).��3'�W����	ǽ�A/	^�����9ݵ�NH\g}$���L��ĳ�{&7�F��(��v���B� ۩8D?}��@��cf��X.�E`��_ͤ
j�D~�yl7^�Sm���Nrx����]���<6���'}�#���m�R��jU�l�0� ���ݸ���Ya)����E�hA�A̐�л�/1$�A�j�M���ٵR#.u-5S�u8�	R�U��T�߃i�cTa\�b��Lyx�E�����z�_*g23���.���^(�h�|Z�|cȠ��]�L _χ�\��7I�/��A���'�dM	�|��>���|=y�&B��}���)����;5�LaV�wԲ��[$�Hw���6p�����W�)$�h�J ��m���oJ��D!ٿ����u©u�]���r�`<ȼoxo1`�P���#%��ȏq���"l�Ds��հ�SE�h2�����B!���f�^ ���rxAdV7�P�ؕ�"�)-Ɏ��a���p�˘|���q��lM���J�	q�F�������i��[�Xj�
���?�^������qN��#�h��Bv����|�ߕǕs[iO���'�^�}K�BmQܯ�#}į���&��r����+���N���*e�
T16��ނm�nGN�uX!����cp	ɐ�w��d�?ژ���d��%*�No��KG�Yr��ˠ��!�L���j�;(��Zv2�A�/,�c4R�Ad4}�p�Og-��u#���;~E�i��*�h�[�y�pˤ��R�hC����u��x��Y{FI��� ߙ�o5]��K�P�#�ߨ 9tq]@���1��HNE>�iSo�i5��d��ԃ��M�{�D\1�\�J:^����)�����s�ü�>LQ&jE=��
�+�6�:�}���ʒ��r%+���$�զ7q�����(uN|Є�7s` 7�'!�� ���d�{	A��/�ևrA�כ�.��D�e������"��֧W��Mo�y�4\XBQHǷ'Ɋ�rp9f��쥾��H! T����U�zX>Zq��q���)ωRH��dʴ�4�&���6#���N�a{�n�@�^��uqγ�U����3�oA�6�˿�IL?��胾���/%�0O��2�<�|9C�ۜX��.�8��c,Tz��P�<hG]��z�
����Oy���IGr�3���wѪ����hHp�X�VM�(�t��;Ke��k5�^��>GE�+n� ����g8y5��F#�?S~�
~ߙPP�p�2���m�{2����D��ٴ�8�tE���~A�L=�LĸH�)'��u����c�e������'�3�ӗ�ݼ��\�˫������Z��q*@{"�0��"V��A���wO7,�~P�KĜ�F�C1Қ�a���q��Z�#�Rp�N'��<�5�ItSˮI"���bã����
ݙBi�+��a�+.�����a�6�P���Cwb
Xn#o�t�?6�xr��P@�Kt���>C��Hd~)�\HR=�-��k�f��@��pP��}tSܷ�i�8�?;.T�!��t�H�`d�+�
�2�Bt�̴��U�k�-,������M!Y*���0�u{���������ǷK?�͖;�mM{7��������Z ��¼�$:$�a�_�7�XQ�=��!��>مB��k��\�6CDp��-}�
���L%�j������u!�E�2��t���U��>�i���}�N�F�)�c,p��+����v#>4��Ȟ�48�����1��=�Bm�PeZGHz"#N'����&���welZ�O.����C�)�]�@n��_�U�Ǵv�R������S�n\�	�'u�`����uo��VT��f�_�1����h�߶}Wt�Ҽ_�Ya�������Nc����q�@Jp6l���_<�&T�����;M9�|f=�$Q�Y��-�Q��yf5�y<��m� �D�^c���j$pp�F�3��/��b���_�Ou����	�E����<6g,���g�M[��y��ܜ�0*���d�6�(P���Z7x������NQKS���qW��%[�k�U6_x�}7%k���P�ؔ��S����Y�6 �md!�*�]	�`���]`Li�5�k�.!�Q�Ƣ��>I5���%@�6�z���oY\�[��M�j� ��e%@�/�y4�l2sXȗ�x���8=�pWa�Kښ�� ���oSi�*>�隴2֪��L ��Q��u�%�75/����U����P	`����b�nm�a��|��Q(�����&�<�h���B�a�W�M������(���@L�⣬��6vh����g�; @w>�@M���3~��u�Bz�i
r�B��^	�^���d��T"�}ÌA[�!y�X˴���|t�o5lGИ߯$-�����n
�H���;��}`o�;$9k$�T9����Oό���J���uc���1J���:�&K:�|�	�i "eGӴ���Fr�Ѭ��Sb��'!c����:��YW$B%�z+�V��ՅۤZZ=b��V�������`���W�r�vWV9I��N�"%3��K�̮qSz�f�?b�5/��)u������VX���<���́"^�}<��0�p�����V�O�#����Xq���J���:�`a��Z�5j�ֶ�������4�C��ᅁ5�ą��Ľģ��~��Ο�8�ڦkx˂n}�f�g/zϗJd��\�ċp��I���d��:NBx, G��?�TP6�>-I�����~RE6���!G��Ih��1��h�rs������'�r ��R���L�l�������T���)��/J%Q�pZ�{�{��a�L�/-�ɦ�(�uRϴ9＠ �k��Ќ���=�j\����~L�K<1�|�\�q"}g��i{8�X�c�w��`{C,��ۗ�\��*�K!���dE����?�����nV��uHQ�yY\����^^�o�~�$ȯ��Q���J�4hB@N-���� |Yw�
�ae^�^��iE7��f�ɞQ֣ۜ��$�w-d��26ɩ����+�2�d䜤>��C}��L&��BGch+��*��1����R�a�2�
Y�Ԉ߫�Rl�A�3��^�5�#����b�mQ�:#,
�b�b��n�ė�1��#j�I�>-�\�|��z�6!�6ĵ坂�;� ��ǽ�s�뗱�
y�6�$��4�l�7:&f�߸�&�#r��"�b!ⰇN挊L%z�o�EL�B�}-���х��+Ds�$x���g�l8G���k+�XA�� o�6-�K�	��f�#����hi�t;t.v�gC,i�Qy�.�ة���Xe�Q��s�J���G�"i���l�ߡQ��g���0*c���\�q��@��w�$��-�o�4ɸ��T�@�6��f�o(�_�6BN�}�Y����Z�r"��S/:����M�t�9���Y"�ʬ4�6�Ԥ��s2�V8cw�4���� Օ1��[^>��7R���o���"Lֶ�m9�9'����;�̉ ��ӛ`_��o� �[���J_���f�P���	뷟а����}Mh�|c �+e���ͽ�����:�����<������Z�Tz!����4M����,6{��E{,�v9T�oz;��*�i�Ӎ�����I�B�C�X��حZ!c�N�CyP���m�&�zj�C�3�d�.���S�z,ۛ��RX2f,�~V}��l���kj�����֭2!�w��ۉ&eO!����~k�PM��q�!��oMi�z4�,[�<������C�Kb�	T�{!���B��_�Pk��i�*M���B4�Y>���tu����"B���������9:d���쫇��OG��,X�Fk]��)1�����2俊�΄#zk����*�b^7��(i���4������z�֖8��t��qe� �L��?F�.~��O2�Y{0Ku�#[�����&��;}�9AY��&hWղH�Ʋ̈����w����@)���^�����B�W�f"����<�hk�^�=��L<G&��|z"��ҼY*�wɄ�%r�o�w�!�wB8F�L@�c}��g�T�d�5�������,͐-�v�
5}�����G2�;A)��r�]��T�ӇUE魾�GS��RF�vr`x���14�:w�K�nq6 <���d^��m��"��e܂�z.�/Q�U���'j�WU�m�̈́\~2p	&�[�����!e\��3� �ѥ�����k��{�md]ڮ�勰�f�cW��Bai�9Qpњ d�8�[�݉�x5�x2�ۚE�4�QFA�vq�l�$rNF���Nٹ�5����	��2������՞�gf ���py�kx L��N����b�˒s���u���I���qr^[��$$\+��_