��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<�y'�I�z�OB�N��a��M�����`��S| �W��̒KJw6s��	=�H�t�4���`1�3~�aMwI(N�M`�P�t�7���R�Z���nD$�Hг5%tޣ��v�I�9M�k�Uy^����.1�q�跻J�Ww��&��u��g!�U��^�n����S���׊����9��fl����| �Ba�c��)C5����z�e���f�qA�n�ө�2}L���t�)�Ӡ/����ASTu9tI�	�uZ�<eB���%U�v$D�'#|�ھ�V(T)�Y�� p�X�wǗ_%�i-#�N�����^�����>�Կý���5��ؼ8�:��1i���h�� {H���.���0��|uh�ʹ��ܓǹ�a�iGWK�T��˿`��jD|]sx�#��s��~9.�S��j��g���� S��������r�	��_�6c��L���h���&Wl�AuK3#2c����A��"��>.E�Fz���UK�pP�4�k0fB���:� }�F��x윞�j�u��o�5��uR�Ցa#�ˋ���Al�����%^n72�ӡ��R:��Hr-)�I{��&�z�vƖ^T�e5��B�DCǕ:�	����ð~8��K�2P`�s����ދ��?���v�GU��jYjpK��+����/]?�)~	�^��	�pp����������ra
�wB��F�%#|����[z"�%�^쁜k�ӭs�!ӹ�#��!���*�Ąt�IpX?"����~��R��t�ʆ�Z�vyr�a{=��FK� �8�`�X�������Ѥ%�����H�'N�n���S�d]�t�9p�z�e!�ϰY�7"G��f�C�Ѭ�����^/DuąB�2�4���#E�BN�}΁B�7�2�gQκ�d'��1 n�T�^����?�dp(LPN�E�����������s{��� ��xA��x[�E�}�D%I8ɥ�I��W�X붺>��[V�6�Ԍ4x��+Q��g�ZW��`� ����AER�*�H��E��>~�onZ�X�Ǐ4��tՉ�)MM
�jx��f����5����2-� ��$m�-��0��H�}���đ��,$O�t��y,�/[2��	�]&�&��
��'z/��Z����|����z��G������Z�1ͯV
5E�٘�k 0�1R�fEB��o���5�\c sQ��R�!���5��=λ�F;������}���WND���]R����rd�X44��9�u���T-��U�
�FhXz` �I������K�ǎ0L��sjX�/��^>Q�Q�����5�?�c 	'G�vy�����̀,�Ll�՗�<I������3��xn[:�'���r�5/W����Oz�Q�zF3��憪e���ޙw׵��Ov@Ǭ8�"'���͝
E�.~TL�~��*�T?����z~Za��Amd��7���p��'���SF;�
7�}9
���LgY�=���L�6B��D"aȸJ�-{����4a�NbV�� �PŤ�*� S�����Wh(Wm��֩�\������^��c0@&�#.�7�)ZKP[�]� .�w�A���2.���AC״��z\��~�$�a�nda��G�PW���f�^5��MpB�H!��
���TC�ϋ	%�R�#:�2�@��"�,*;�ӂ�zɨ�a섰�ZU���A�Dǒ����i3�-�(vU3��{(��wd�a2�r\QJ_��C�^�Bc��Dq��6qF��@D�Ȓ_����Sk 0���x&���s����r� �s�5�q��>e7����c��
_��5��Ԛ��#Uu8�J����~�%��rJ,O�:mw�,[y�ͽn���.̖*����	O�-=�P��>p������a� &�6�E�)����4�p��a��*8���!���]3�|7S�^�J;�����3�4$(��F��m�0}.��������G�Y���c'��Ѱ�R���L�r~��[ȄL�s*�[�P���,{6�?���y"�1x�����rW��Y�4���P�˃n�M�p��>��Zh%?�^�68m'0����XP=jԑQ��
Ϭ��1HSu�08t9�n�Mv��<�qi�gՋ��:\{�Ipu��!�Z&�! �m	>B��w�w����%��2,��d��2��?j���VҊWt��71:�2� �'�-�'���L����1�5�"yV�X�4
�n�qb�;�ѫ�p]	*dШ�P9lgH�&#Z��'k�$�F�`�YϝU�"Y��ބӸ��益h4���Y��9�ƽ���.���}����0�j���lۃx��+Scn@v�2O�<6P�O�5��Bb	 �ib�2̧jQf�Et��E�Y ��.�TE,�.��f����#q㠍�fd�=B!\���-[X��M���&`�����kk.���������E/SZ�ї7�i�;<8�$���R?�H[D6���"L�:��V��]�'�J�0j��< ��!�󛬭:V�̞]k*c1�1��B�Ze|��#���.����5b��bmE�:�2k�U����g�i��5��Y�($�1T�R��Bi��"�=�p��W_�X� K#%#&�l��0XiM��H8�X*��o�~7���iΊ����v^EBZ&�C��l�"L9���CSf5z�P�}���	<�P?��ܡ"�ء[��&��d
\˟�3��(�i�2;�)�$�v
�X��������B���٥Ma�/%�b���O�huQA�2/�����Y��=�� �Oo�T�:=�[v���@��E��e/�k�6�P�
�b�k�&F���4�*������*̥��5��B����4����l"�� �f���jcD�LClRU��k^˯菿
�#��e�o���;�����P�Ĩl^in<H�h����
�)���
���޵���d{��i(�<�!�#1|���f-ֈd��y]�� ��F����L��Q��9�Ң�^��Z�ǥ/�ҤEw���-�	�RC2@��^Z�C�f��ͫad	�W/����Ibu׉�T�Alr �?�qѬx���	���53\��cn4����C;lf��C夎6E���׊�_9OZsn]{�.
���F,FZ*e�	���R��٘�u��f(��5�  ���Z��e����	KMh�y�`Փ�U�Auk(�i�Fe�;�\C��I��Z$�{�NZå�wBM�X"[���oS~y�N����Fjz�7�W��rom�}�Զ��#o�"�I��[ٗ��N?�����ᢒ~��/��}ӪW��`Wh o�E����ժ��QsH��=ݲ����V�ަ��A�*���7�:��g���ϼ�3��tKC���C���ݞ b�,v��x82{���۝c`:k��
J�j�A�@�a.�`����CF^�o��upF�r�6^�|w��S�3�o@m��D�1F��@F��`K3�P������4��I>��bO���d ٠���V����Y��s���m�蝩(����<R�D�"�̖���O�)���lHL�A�١YR�o�6Fy]cM����D��6=��C����hV��R=���:�k^'�J�YM�9ᆤ1 1Ԕ��T�
~��rDF5A2Z�Y �5l%<snC�Z�p���Lv<X(ޗ�g����R�>�Jn`1�f,�W�{t�k�m��� ���9$-����R,�8̬�*��J��0|������O ����9L�-���!��tO���_�KN��琎F`����5Θ�9���ʩ���tx�8����;}ȟ�0�fY��ER���;����4�������EF���1c!���1���:��=��1�������Nx;U(N�x;�-��Vg����m�Gr���|h�Mr�G���W"7�_�$]E�F���PƝ���^���et贔 x��z�� ��/� J.�R�Чc����{O�E�A����XI =�%Yp��+_��,�h6Rb7!��q�&��_Sr9U�Nޒ4���L��W��~�aц$�3W7�����>�@�=��e��w(���,�]Q�3 !i�Q]QL����҃�zr7���:[��^�7a�ZO����i��I=Y	�a�����M��Y�Y+%���#`JJTmpj�aQ�		"h�e*��ji����b_3_�	�F!"�jS+˲L/����\Y'[��P�{��s�9.�*�L
�ڿV��r{�i�=G�p��WMWH�I��c�	.;�0Hj�չ����T�T7dGtY���a�i��
_8F���O��p�3J���Cy���C{��1�X�saJ��þ���<6p�E���<��WM��)4C@�:�F�>�E�[?�4K���e{�6�%L�%���Zd�^�7+z�|��l��Nj�6��NG��e�%s�9�Q�k���߷
X�7��壓�\1\(�M�j��-����< I��]�PX"?A���XJu9D��X8q�X��ZH�y#<���^k�H�9\E�ޯ^���4��2Oi}�+����R�dzs��T�D��{�w�ϛ���	:P����ˠxg�crA$��Դ�-kJ��H{���-=]ɇx��bݻ����O�)8�w9�wg���{ |�7:���c N �#��*�G��&p��kgiqHU�"W�H7���>Gd�e��������_���jG���=O�|�z_�^�c����9�$a/�MP�٭lg�����B��+Pt^�џ�F�3���++�9M����l����n}K���	�;��4��搶BK�xu^��	�� '��~\%s,��A���l?��n�e�m����s2���`%s����K��F�h�)'��p���;�����Ū���6Df���9�4�c$���E�3ݐVB�&#DX*��;B�5��+E������
dy����f�ٍ���jLJ_�u����V�O�6���$^�0�;�@Y������W˔��Wa�.u����lC�A�Ea:�??��g�|��y�H�<&9	uO|��({�������1^�Ü� ���#[�V���2�J�aϤ_����+Qy�|]-߰�[� K�i�&i�2~� _� �����}�x�k�^�15�F�)/ŧ+X�����D��B��"�e��ف�ob+۸��h�8#㛤j�9�P:��$�
��2;���q4TZ�^�202�*�bD. �<��M����j� s?���`������%���P�t�V�<� 42�HȧC��J�̋�����RS�����=��:1W١�[��;���^�����"6�N��ٳ�IS�_��q��"�l�60�a�Pu��0�~:���e/�wJ|�ph�ۯ!$��c�)x�7S�������b��?��ʮ'�H��R!� e3N��d6[�zy>Nאm���� �m�Jɖuu]���l����i���[�����y���њ{�� YZ���3B�Ѥ�8�I�mB�?# �1��l^�>���\�,���&�J��a�Ñ�ͅ3R��X}�6���:^QI�}�]�F��̳�՘�E����5z��D�`��f�+��@<#Vn��Rߪe�W��u�(��ܱ�U*�mW���ޤ(m\P)b�ӌ�}��
ǵ.C�'*/�g�qd�/x~�K��4ɍ�#�|����w��h�m��Х���4��ݺ��`�ZL0�D��C5uPJ)v�:�pب���5+�ǅ��B�EZ�߯x�)���s����_����{���MHPp7�
��d�>1��b���m�D���dN|u�t*c����l����^�c��/G��G�	3�(t�n�e������^����Ph#�=o���y��P�����Z�|b�JbB)�Ao!�WY?z��[���[��P�\:iHnq2C+�����PNb���`�pM��:�?tՉg��p�+鉘��$�ʎEͺyHW��Ӯ2����c��㍘ѧ�i���H!�_�O�+���(��k�7I&��`� m��f��'�.���Lzb��^z`���`�ц�Z��	��;�5C��;\��sG[ܰ�6��Dy�C�Ӝ���|���h`�7���r�l6�
���u����s~mp�Xb�vv��X�!��eMB/n�c�֨@;ۺ���w����YMj*djy���	�,%�Z����	��ZJZ�8\�3R��8�$pz��� ���CĹI�#��ʼ��	�Mx��	+�بV���A�Q4�QL��~Fm�xI�Y͸��bP2]��B#^VD�?驊k.kJ-��掎_����[1�h�ӿf�L�DK�e�
k�W.��*zA�k5X@N)������S@��3��~��k���k�\f���Y�H�7�,��F�;y(�x +�4�]k�//�g�@x�^�0�F�nť�КAP �'��5nM�))��R�~��Pl-���$L4L�7ȨL�N��\���S��7�d^ N��P�('�xR+��w?�{'3 @˵�R3�7V;��̞���P��8�ߟ��]�l�^�ҎZp%�t=����15Ħò.�{hI"��� ,g��*&�z��E��[2Ņ���a�q��������"�uc��}'Q����9	{�i�	��J�
Cl��	ڀ�۬�"�h��g�HO�2�Oj�ԇ��*|�Յd��Ͳ<;�0�췒���z��23������[7�9<����=��Ѧ�Ql)