��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�8k�)9�k���J�f ۘEN�R��>�Ug:�&�1Z�G��ZnM�X��l���c�g�J��R��x�D�35Z0��%=y�S�$n`af ]�z�pl�4ƈxS�ԉ0+y�H�X-�q���!�R�Hy@�T�ü���ϗ�����T�y������J?�j�=���t�D���X����_�v���h��3��c����`�s�z�й��~�4�����Y�})��Q'QK^�+R`�I����+"4}0���b+���aX�T�1��S?]ߌk��gڵ�Vۋu��c嗒�L�;0]��n�a��(f��s�Q0��⁇>]��$p�QjB:8@�[2������yf��d��c�	��&�ǔH�\l��%���Dً$�:HY�	wm�~��Ot�SR���;�I��̜�K��肊o	FTVNj^v2kee����
�;J�z�l�A�x��"��tFAy�&m�oL`���z���Yl��
T�&�`E�y8���Y�
�T$����W�{���a�Q.L36	�Q����अ$fZ��=��q@����+�hZrkhz߫zʼlTIq�ա�F�э��Go�&�S*�D��
�o?ފ=�i�M�KX.~uF��!��������Q@w��Ջ�q3�x;}R����E-��"��O&c o�6@V��p����%�7���hOg7�nswa��hy���T���u�#r>�1I�[e;|=螈t�4��`"K��V˸��x
�	���y)L�g3��!�*�� �!(kq�/Q���,��̓��n�)+����Z��X�yu2�{PF�O�q�{i^���E��MK�/�Qf<63�*R	��cU�tT=Wa*rBƌ�+�?�\�@�_�z�4��ׁ�ilG�����.M�V�}�W���xd�W_H�u�L|)ֳ, w��p�p|���V.v������0�p;�/L7�z����:��	��0��,n�z^��b"�p�Ҁ�k�Gn4�h����pq5�Y��g
^�@l$�+ �Y��U���QBW�UXo.l�pI
X	jKX�L�~d0~Pe��_�Y��N�l���_�����6�>x7K������v��ÎX��=P#�"�v��&+��(���cH{���}���`'Y!���h躧�Ox�Nl^�{!����[����yN�g�x�������O�cڶ����cv���,�����o
奀WF�Q�p�CbV�v�� =?M
nkM�e�x��o���;���B�����V��*b����u߂��F���y�R��v>w�׎kA|��CŸ�"n�&+�Τ=���;�C��
�xTz�	�UZ>,���s8�(�y��n���B/�Z�b�)�(w&�s�����B�W衑��Y!�H�R�pRUhOc�n��n>�sT'�M�׈��]D��Y5j����sy|ؿN	� �O���>�L��|̮gM��c�Q!.h�"��"��̰�g��A"��� �"��+M8�l1tvzk�2�rO�_��)�"�1��!fyn�1u�E������RxF�KIC

mB�8'����(�9ɨW"9����E������ �� ����$�D����]9n�����g���cBXE����+7@!�C#Ӑ��(����pXo�� FPN)�[�r�P�UNxl	4��V��=�q�=yL�  �x�k)h	���{l���^\1�Ts�Vx�Ok�`��~|��Oϻ��xl���Kc��W�fOϸ�m@�<e:��S�����֋�Vff*�� Ή�}-3RÑE��Ԯ��G���8�,_}P	n%W����%���6+iZ��e���w"*N��d�|}�U��F���XS��Z�� �Cp�jp���ޖ|O<�vW$G�|s�)7,���w/IN��^���u��b�?�V������iи>Ŭ3�	Y��S�`s"��Ů�,��� ������7�tY�N1Uel��H�T����»���cLx6/�ɓ��y�ʖ�J>��ǯ��G� ��YO��In�Pv^N���΃�
D��n��qw��9�P�Rd�bfj���6d_��]�&�ǌػ��{o��h*�-	��!��%w�(,�j*ؤ;n����:�V#������EHqi�c8�����i�3�����K�4@/P�8���CI�߭�9�5.�����CdZW��������3ߗz	[�csn4#N���1f����_�J��瘪sJ��X���i����ļ]����Bw!���n��R)�yf�l��k�ǐ9u=���6W���nE����]��o���ȳ�H��x�� a(C���zgf�:��YNP��^+�*��&cٕF�n㔳�}.�;w��c��f�y6]�=#'��O��uN�P�lˀs���6N��B����Nd�`�~��\���>�Jˮ����;���s]�9�N�7�~�Ti��=���&�F8ԙ�ھ��M�
�QR����;&���r�:!Ā���I�Ũ�����T�2^���ϲ����H5h�]����'�@"C�9��$�W9[����`KM@�)iG�P}�n���0]���b�K�~��l@�ьh������ǂ.G�!���$�t f����v��}k;,E���`F:Ҿc(�V:�d��g�ܶVƒkYĥ!����`-��yg��m�w�0aeIl�0�5�f��fR%e��]i���Pv�<�@W������'��u��1 ����p�� ���c���@��*�ȝ�+2�����P	��6����"�t�W8�z�G$V�zS�� ���1Ō�����5b�X)/��_�^U4���RɅ�Sw�L0k�9�#<;1��(��\��FI� ���k9��g: ��A��L��7�y'����:�/�����|ً�=�����+�WHb�׹\N!�8D�f*�iSsh�`���ݎ2;���[�N��/�X�<Hwn+�C��-�M�Vt�]���j�l��(`A��yC���L��^��%�ɔ�}7�B�X'+�ޅ�
s��O<�/�z�*_mߠ�N��븕iy'�*�������QulQQe�G2���Q�H�$?�� |9��+����s:	�	�6!�ݪ�e��m	R��i{TM	x9�
�1�h�����Zs��=OUGL>?)�{��1ԥL��=���#���.���\�L�� ��z�_c�s��ʚ�*����&O�F��O�B�-��IF���۾*,�'8��G�"�̏�K�޿��M�A�&��{��녈��AΪ�*_*�����hEޑ)� �I����w�e.�Y�w�V�h�n���JqZ;�?�%�L,�EY�N��(,	�v��xMN�ܪ]�U�X좏/��$m=���	�g��zϗ�L�Z=Y��;=
�קB���6e�X��?�~��Y��z�i�#&�4P�+��TZ� ��`��$po�u{vEMZ_�R?�K���k�b>�G�y�q:T�&��;���9��:�<ĉ:t�Oʨ�8�7Rݰ���C`r�k� �so�
��(�ۯVl�P�1�##u����*�V���Ӡ���5��{��P��0�;�n�Q�z���po f � ��еW�W�j���3��=i��o�pLpT��C�|�ն��M �K	�W[+� ������ݕh"�ÇHA�<ћ`�O+�/��u�/e��F����:j��t�������
����c��4��AiO�:2V����+��.�4\���ǼC�`Fh��]�cXP�9�_D��Z�OƢ�X��y��l��m�p�=���	<G��c��}�y��_�Yg�z/���ym�e�ez��	W���
����m���)A3����n��i)zmU�_{�t1
�_��Q0�n~6Z'�����a�3K���8���_bͥm�Q�����CꞘ�O`�b7x�XĂ Ay��>ѡ��G?�	�Q 95"�N<桲&Ll2���� =Q}��I�Ƨ�ܽ�o�[�2�%�����u��(a�y�9yZN�9:�������Lr��V�&����{�[�g!�-LW��Vhf�d5���Z���f}f6�i�9BB|�����F�Ș��G���FE�z���Ǵ�����/Ťu�ȁ����=��W#P���CFu����zM|��>�)U�D�>X-P"��`s�䨂�5�X爘��G,�=-u�_@ZvGw(B�2�T�7KUg*FPÃ{��}wwV�M�tQ�]�PʶKi�9΁��u�5�aC��k�A�����q���F5f��y�Jb8h��6�<1��5���7^[�ڰh�R�80k�R]��_��o� �E�{�s ���JZdM]c����8��9تD�f�<<}�\$��j�؝��4r �3%�?I�]�{����-�RF�Vݥac2?�7�x0xZ�H����`�	�;C�2pcx�cH�R��:"�����Ʃ7�ɵ� ~7���O o�z�2x)߶�P�j�4��r��:��W�O��`�js���߳��#Q7Fφ,��N�΢��?=�����kC�U���rb�l�$C���E�� ��FP?��&���=��7��DN�5����!:�6�%��D����5m�� `�۴�)��54{���"$W����Y�t����?E���Q��@<�..0ͣ��5���79��uq��JV!t� �H�5���b�o��J����&?���\��yT���x�e:r$�O)��vׂKpi��/7B�G�? s9�Ku���d�wQ�wa���W*C�{��ʦޭ氓Z�ڌ�����,��NlʅˠQc�^	��fH���_[���N[�-�m�cki�9_��A䌺tI���]��R2|�*�:�)��V��΁z��?�F�G7�a!��+�_K����|����}�����$�A˞��aG��7͝f��w�U��K��xU���U����
&U�8��@wE�n�LÑhɣ*�N�x�:.�\�E�i>d�2�	F��"��Up��'L�,:��k��Lԃѿ��Wfb�"%6�d����F�9w���9�"	�����y�7�&P(;�%욾�� ��D3lz��T��SB��E����U�=<���N�{RY���ȄC�#�b���k�u��Rno��ͱ�x��o��|09�Ȕ�њ.�$�0j���	�> u��U �Y�xl�q&#֥!e4/^m��z��v�D�Fh�*ZyKPMM�"ڄ,��^4��`[Oaʩvu���YP7�*-��
7_q��ݳ�A��o�?� �Q;�6��п���`_�]��Ss�`���ƙ�X�ء����@�|y�g�GƂ��!���_��u
���!����i���1\����L��^�w1ŝ�����p�MVZ�2%��'{;:�'�a�V[�����X�K��-7[3�.���'��Z��z�F3�~t����֨�j�d�
����o#�S�7���Q���Ƚ�vo�:�.v�h�e��֔+���*�^23�Q���b��i�f�� �K���W}�.y�t88��8:�F�F��O�������J�R>��kt�������.�&g4Z-W@��:sx/N0�i@��2�a�UL��M V B�E{"s�q��(�� �=9���Sw�3)���5�1\"�{ڋu�Y��&�j�jW�Z�Dy�]4��H�d��D#���Rs�+zj��ɚ��=�A��h�����K��y)x���rQ�P#�޶�s���D=��D%J���?�Y��c��7�A^�>|X���
2�]'\,$1ү��� �[.-lU�B+)#�#I�x�`P�C�wȎ޸%�9�JC�4s�WZ��6b8рخ��\�4�e���ݐ�b�@���d!�^z�~�nLd�)l}���U6��z`�lx�V�Ou�f�����N�v؇U7xb�V����L��i���5[���U_�':Uv@�E$Q���X�r�h��^Q5z��bY����9'��1��!&����S�`�Y�����s5=M��(��/6�F7�,�i���`S�O9����4��(�;������������I���k_�e��
��$Sl2��ˉ)q��}w3t�)H3$F��E��Ƕ0���^;������:���1	��E�>��v3�YLi��VZ�Q��T�����6	�@���?�K�6dp��)��Z�93HH�T��ߖ-���
؎��lbp���\J�+�LB���v=��:US��_�mg�z���V5o����p�_���R^<�'�ȡM�z���*�.!Ń�o'�<_���*�.�M�A`}�vGK}x�OB�0�VQ���rG u?;Jؼ�E�fz���M۵C�h��ܮMq<�Y��L��ٰ��P��ێ��^>�"~����s[j�hm܌97��f-v�$ײ!2j���s���w�id/>�}dL��ϝ��["��̋?\F�L_�:�� x���Mb�N'S����O���^�a�,K���D��)����ZbJ��g�OU�$�.�	�u��^I��x��E~�<�"dϖT�db���~E�X�9��i��X��S]:k
�OT���i]�^��2%'� �ĺQ��MهEEF(�y�|���})�z�q��r}dK��(�2�s/'c�d}[K��le%%}�6)�\fWfsɖ���A��a��ǣA���O�'��k������i	� �qBjķ'�@U:�;E�{��۩�v3K: #�t�RN���BI�D��7i��\���y�Q5��5��}�/C�@G��H�7=�����7�����/7u�c��b1Y���.�垵Z�=��{��q�P�o��J�΃q<��9w��^W�A@���A��N�REug�]x�Կ)F�i���Ι^'����[�`%�y��s��i�۪oJ�m��M#Ӫc����2c������&��<s�4<S_�9[�X�VJ�/�R��6���lz������&��e�֭���̤j�Cm�'���}*ȅ�wO��m�E�'�f8�9�����б�Y�LQQZx��Տd��:����e�N�:��DGq��P�80�RF�Z)�:㋲�p�� "����c%J�!��h��Iß�6M�8b�q��L��k�Т)�;Fo�}s��T 76��
�}O5&��ߑ�D��Y��?�맹��!����Q�+ }O��DD/��!uu��=k���V�?^�¾�K�욙GV"`��<J�Q���!��{L�)�/�3�3U���[�M��)�`;k��C���1�r"�w,�)��a��q���N�����?�z<O��?gġ{�^>�(-ak1o~��V�ρ��"W��tSY�\�|Rt���5���f�m�ـ��J��؄5T��e����{̟/�9�E+���`��bk4�o��Gr%�s������d��}��+ӐS��
�d��n��ȰdݘY,o���)2�Ͷ#� �ׇP�I���Cl~SQ�y�oYrn���Ʊ��j���y��2Bt�Rƿ�eNt�M���5al�e�i�ihx'����J�d&+�3�����1z�f_+K��$T��jq�����A��c�� ��P��`�V��3����(���P^�f�z�h�>�v�\����[\��6<c�&;�r\��&B�0I]H-o����h@����U�
B2v�4�9���J����t�����s�YE�y�U2������y�)L:����y���q���J~M�]K��j+]��L��9 �2B�.��:�U�a.���ė�@�`��&o ���ݭ���N> �`s��XR��;�"���#�Zhy���kQls�7����l4�/�)������ր��nn6�|��*���B`��lXq�q��P�Wń4pIu"����H7�� G��u�i$�G�����h�MEy6�U�"����^$�����I�Y!0�aB�ű��-�k�mҙ_���1ȓĪlXϮ���9g� @\�$׳(���/z������q�!�F:=*B�m9V<`�q�7�Gk�J7B�ȇ���%G~] =���y���xأ�����2��5������~�s��˫cQ�;	�5*0��V6�JHJe��(���"b��A++���t��l'�"�쐋ѴS��G�wS��	�����Y��.Ĺ��>B����Kq앋N4�ݾ�sV�RIJ�1n���ez�2�2��H�ê2����;���wR�)�Q��x����[m��{@���3E�|l|u���QX��W�`%�e'��^ر-��C��*��7�D~q�4Q�>����׎��3�Ęla�<zG�3�ʋ&JY��@����.K�7�^��a��C"&�/��c)Ãl�d�M�<��5�Õ���;������5<*�|7��_��<�ypa/���Y��	�d�4*�&�!<��3���.���N��OhS�^����91��<J�i� MZ���^��T����r�݃ 3_^�g��lI���c�':}��犻T�}�1��!�N��+�A�SqѭR�4��¡Zʙpo��T��N	����0�j@3�|�EدO������b�����@��R�BH���c�&���2�-ђ���/u��A2���e�,2F���pXp��.V\e�A�-��H 2�)��\�7���Uuw�Z�
��I��<A(I�u"2�[�X�j?��+���ٴ�>�����Bg����I�}s�L�8,ڹ��C`-���+[�;+�&i�(c)p���D%��,�;�z�m�is�N�n�Zyj��װ���@7����AS�������7��"4+J���E�N�����1s'~��tp�v���on���C�h�g+�I�t�s{Mp��4Q���*9*i�_�\UO�8�� `��Z��c��efB@=�r��P^s�n�!�Qc���c.��\l����!�n"��'�n��y���#eɐ��o�����o񡼝��YJ�+PO0��kp�K���Qg`ʪ<vhP*�VjL��R��yj��&�_�_�VHQ�A5��0MK���$��l�N*�xe��|&֊�K �2(#�2�;�������>�wE�z9����5p4M���-��1�N�+c��.S��F;���[`֤�_P煚�L���z2P�Ɲ��H�r����x��?�B\�=����Ee�a6R|����G("��}ˡ���O��9s;U�e��R�q�#���=*d<ƻ�M�V��X�~y^�xƠ���^ZqA��\�1���Yռ��߁��x�C 8r�grcYH���}Y#����vM�[ <,��l�z���u�ÓS�\���2D�$	��h��AA���������n���<�+�h�&4��pO���BȠ�0��Q�~�ؚ&D��tDګ�┑�����k�pC��s*�%�
=_��"~NdwA.KPk������5��g�����oCgn�pf�G@��)w��F�w��$0���?�;v��
����=Y��䅀���;]�p�Y��.�����C���ʇ�%
 �����W�~jnqgʫ�)�K_g�jK�VV�v�||ƓḪ�����5��U�IA7T�7����o�K�Wl��X�u�r����_g��R��E^8��N�u\s�xq�7o�H�RV����	�r��E��.6\ڞ�a��}q
��`ݦu{2Z�U�Rw3UIK3��o�f+���/T�� 2|j#�o.jL��'��	9Jno �|@!4�y����m���e���t��uԬ��Vp7����}��E���S2�?���(:��H�1��Q-0���6��T�#�?\;!Q
�.��_���aʶrWw���Dj�+6��)m�n��L{�}KG�J ���R�#v��)J��s5*��+E A���-���Ԡ�Ί�;6u@?��Z����^D��� ��Y�=�|R#��Ci��\�;�/�~`Nĵ@�6D�.������cˇ��
=V�0s]F��;Z�w"��K��j�v��! �6����b~b���{��x��V��!��3����?�*xV�����s�0+O�n!��\d�-=l��0�vA�$���!���/,��N@�b�N ^!1���]���Y�6�q��0� �U�<���J�����\�y	�$o��7��Zy���{��+<��6�[�2�ez���kV���Թ'��aY�wH��nx�;���~ V��_.�����\��d�0�x4	�π)��^"���4���	��bb3�05�(��k��5M"$�$��
q�J��a���"��/6�v�Z��ՊX-��7���B4��
��M�5����4�..��������[9�D[C~o��I�o3-8�������R���O��HB�c��}��S���i RN��%���y�����포i�����G��㒛�8	x�o��j�%2�V�\S%<A��ҥ�nF���h��K����}C��ۓ�K1l���5&%f��`����
}�� ߤh���++�<�T�|͗XYEx�}� 73d��D���@�@�� �}Oqv}ԣ˥6G�p�ߑ�pm��	��{�=�w���]��������ľ��w��[����NPÖ�Dd=�zF�Ҏ-u��h�����S�x�o�����O�	���Ƃ�G�{L!�l�Z����%ّ1c��g�~��l.��Z;��Զ�9��v�
�^��Xk��F9`hj�t?J�ұz�+��HB���7�d��01�i<�J��~�ݼ��6!I��.�rD���HS�NM���}7�+R� )3�Ir�j$#�3�:�M�fJx2X�)�#4�.��*2BX�㓕��@�PQ�sEBy���]�O9���nT{��mf7��^]��������� �$\��f~�g�uBC���6�w �1�",Y��{��S��%	�`��G�,4gt_�5t��a��3��8Y�U��W���	a��&C��M���c׎$t���C�B�|�5��߭!���*�!Y�V������P�S����i�P���&vez]:�C0w��ڧ��z�0:�P��p� �ﯩm��y�rؗ)�ԉ����s���p�g|A�l�(��P	��a�_Z�­-u� Q�� .��8��i�Up	�պi��;������%��2� ��®�B:a��W!�$��`A�~g#O����nBs�&"��J�� ���|U��r��B�l.gqy�:�-�Ԗ���3�R�W����y�R?��7У����Mz��FV�N_c��兞Չy2__ͤHgKG���b ����##�����P�q��YR�Z�T��.Aּ�����o^��ߊ=���]�z�3n6�/�];;{�*�Q�4y5��O�,5��ٯ��\�Ґ}����L0s��~2���bǄ4�������?Ė�L��*���6}��<�Tӌy��qÛ����6������[w���W�#��)�P����@��w��=E=
��zA9䏻�ߢ�Tκ?	�RĽ���6Qr{FxY�K�����C��q�.̡���v u���ہ"W$�ͭ�~\M��#x���ʧ��C���1M��KX�>��«KV;5���+g��N2!���@���K���n�7L�#i�rQ��c�>3�԰��
�֜������L����Y����?��$.�gTnR�fc*�(E�`+�?l�Ͷܒ�s�(O���#��+�����@^��=��&�4�bFn���3�$M��-����a�Pg�7�C7�}8u|#Kbm	j̱o��A�������3�'�>���,����:w��@���$��:5�U�����=��e��/���E�=t�0��[�AE�d�d'��I[4�~�0�w_���i�>o����ǫ�a�����<�C�j����Oɓ���ڠA�gR�*���C��$�|@���0�X��2S��Z�i�H�3��4޳$�g����H0]���H�8��6Pі%�U��:�ty��BZ�E�h��dD��ʠ
?P���c�,��V�o���,�]�&������e���Reh��-4ua	����$�����Ը2���3��%DJ�#�u���Z�
$L����ɍ�{���i)�f@Qt�'@�p?K�}���]0�L�X�LBwz&������6�؜�I�T�44��dĨ�?�Hc�����6���_�0g����h+|�`CY��:2�-7�x��Uj߮�HM>�\�<�^M���Qg�8�KXX�:\�B~,��XF��7�mX|u���0�|Q[�G����u���#NI>��㲕�F�99ӡ��ъi>F�>�9��=>iM�'Q���;�浉�!���^$��r4F�"3�J�qpϜ���m[H|�� /�C}=?!�`��f%J-i�{�T��	-������nsĎϸ��#S2��D�l���U�o8�7Q�� n�	��W��c$�x~���0G�M��I��/�ur�v�h��Ig�TԺ{v���2�FtT
s��ǝW�>�Ke(���qI+�) �dM6�7�քܕ.�-�7vSx��n���DT��8e�e6]�&b(����J�I���Ƽ�O~�Zkܙ�ڏ3(\�3��q�F\R�'Z`V�;|� 퐺"�oQM�;�X���O�kb���x�a��!��,V�N2�ߪ�R0�<�@{
!f�,��.S��g�m�/G5a�ev��
˱j���3L�wO+.gl�"[H�*��+��Wc�[V/��ݤ���R�6�{��s/�wG�(��9Ti�6�R9�9j�?��k�c�Kv����V�\)�Щ9T4���
�K��>�)P�Z�����F�r����uQ�M��x1���RÛR!����=`�d��#��񦳇¥-L�j~�i�eTL�:������E$<?wU$�½��ɮbu_����"�Xpd}�:�qsp?�g{�'2�XEs�GGP�ck=�2���n{$^�ÌbJ�g�<��|�L�p�h����)�7���$~�������D�'�����g�Et��ٱo��F���oJ�����n9����?�o�z�3����xRg�i����tM��;e��)��
�Q�#Btm��I��0袼�(�gX��a�W��2��:�����~���+���H'��V�Ad[���Q�bՃ@ih��<���
�l�S]��u������f=Xn�6����i�����.�>���\q�u����h�G���L1����q.8�:�S�D�RaD��P��݃���vS��WT��ĺZ�Q�a�{�9��u���ÒnЧ�����+42��n�� <�E�ڏ�>@q8����%�ӂd'4� �g��`wM�@��9�Z�<�@�����ٛy7Uީ6�h�Z�ŕ5�̶�,,j��%���=j!n�a�C:��.�N�g3xtO�C�޿�t���@(qPr���h�[؇��D��F �����t�j{y~�q8&�Z6C*�,+u���zA�z��C������`JmX�kIx Q�j�v�F�awX �&̋�B����D�6�@!��m�W�����W(�=�j�k.�OCL��Q_����ڨo���y���?A�0���!�;й+ ��+�ֳ�H�� �>@������� S�~8���u�p�)�������0�2|�3���i��M�_Z��l<sv�l�Z8^��9��9�����#�I�$-�����Q4���1���5:_\}i^�7��,�X�ֶ�H$��X�$DW���4l���`]|V��#�R�}+ѭ,(P�~�'FR����@&��x���$��aj*�ȃ�z�`�wpdNQ�q&0l��N�Ywv#���:��?�g։�R8��)��/���u*�?'��Hv2�'ȞsA���ō���wZa��P޼9|(��%�E�@����u�|��F�D��;�81��9�Yib��3\�_A���V$�Z�B�-S!(�Ձb!P��q����!�LG̝���7�,hQ�R"c� *@?��=4:�,o���^��>�*I���n�>��M�Wm��[� P���s�l.��KS���g=h�>4X��O�5y��|�^<�d��}��Li�R��u-�BE����(W&�)Xo��+�X��żߨ�b	Nʼ��I}R�b�y�f����^ݬ*����ZfQB�Zִ��֘�Xu-���J1<�^���l��@q�5��n���ʈ�k)���X�Πut4��n��b���߷^���B�e��4W�:h��_��g4!�r\�F!^Y4j���L�0g��h��f1/<���nߗ�����X�!ե�Դr�7�q���Ν��x���dD'�\55��(��hX�NX�e�R����҉��~��4ܨ�o��UCr�V	�˟��K��ڄs|��'/�)y��;xh����o��r �o��Y"�@0>����:�xW�,�=d��%k8�XQ�_i/����M9�3�<�c�ύ�b�j�D[�)��z�BLLu�}���\���n���E�n�g�%�_q)*ȝ���*�bG줤���ZFIѝ�$��@V#��=h���E�x��*Y��L���=ŏ<A�U�Ǒ��,��E��|&�iO�1�:�l���ԓ�)����1���������G+����7(�%lx�=M]��������G9Z�����p6*.��/�n.�Sp ��?�y�_YB� ���F!����у��<��N���'��G&���'��r`�-.��p�Ì�O��	McX|���9���/�V822�𩘡sa�eW���F�������p'2�P:drR�wzwJ��'c�<����^��jP�{[�U���t�.k.�j���-����7��?�/�ڠ3�uT[{���n�Kݴ�!.֊C�f%C���Q�E�8up��������$�*��a��Ѯ+�겊M��a�4Q�5�@w�����P�4��+�# �܃*��	�}0�<68�?�د�vi[�}�Ǥ��5ZW�w�� ���&ҝ!�+DvF������=b���)�Z��~��i�ː���҃�숓5�RP�	]Κp��gV����;@1K]I�i�pKQ���X��_+��
@���ï?9���N�����?�m;>����̜�_,�n����kk$Y,%���e�^5��ɸ�k�<q�Q�2��$��՚�
�����+Ћ�m���tfM�պ��h����g8�h�	��H.M�T���UE�ɶ�V���Q�I�dH�9��͸�g��;��ꭄ[t7hY�����t�7g&m�p��ҿw�9��~�&��6�2�6�=J��.I�Y���R
k�Oi�o˗H1��W�h)#��T�i�n� ���(�Z��N��&�`��&Zh�6X<@�m��ᢨ_�E����:�1rmI�l9���l�0�~\��>o*)�},<��,�>�ڏ�ƯBO�`�T�}��������������Ѐ�X�~��+�5_�z=��G�fP<�Q���S�92g^Vd?I��d�Ťg[Fw��S��ϲ�\*	r����+i$�w�u>1қ��,��P�u��Ga���F>�et�=��p� 4�;�PA�qW�N1���i������DF�ɳ�ȯ�L�J���;��/�C{�	?�M�� 'V��r3�Xf� �i����A�smS��<���ءwCᰦ>�V��e�F,�5#ՠ层ue���X�w ���Jy(��<k�}���xȅ����뫘/A����@!�㨾:`�V^e�fE.�{)�^lP��e�a��C�1�~�w�c}C�T^W?jl��6��d���J����|��"�!�H�戀ktН���
K�ی���@�������:j;d_|��Ե�P .���	pF$�O�ή��k�l!Ma�H�H�@�۹~��k�g�%`�[0^��d_��₧~�9�IA��\�կ��V��@�҅¡@ؐUD͖����%��UUg|;�����'�i��s}�e�r�Z �" zS���JPy�|	�wP�;�~�o�U'E��C�j����.�7��P�~@z��i�^=���)t����':�� �5k��D��h�~�gĢ�����f7@!ub�Q�_^�sQpZ)K+y��O�<��Y�����!��6���Qp�f��������h���`ƾ��z��u����j�22�VO$Q5:9�a�$�i�c�\r��j�y-wF��K�:�XF����Q�w�^������p��^��e7���UL�kq�hV��8kU-�kX��)=_ￂj�9�	�1�����r=����)&xqA�MHI�ds0�,�8��l�IoDr�"�-%|�;>ٞ�f��l�%�:��ꔅ&J�qg�d�	�)���5��(#�ɌHS 5竹��Њ\H�v'?�̙������_,_��~�ej1�7�)��*�j��'ꒃV�N8�r�^���,R��J6�cP\^�D�?�Ѧ�l7X��]Pw�~u�GBE��8\���˺���5D�l��t���cX$��.�>+:���#���sT��<�������,�������3ڌ��("{RUōf��r�I�`�L�ض�N�
�˛%t�+�z�հ;�CV҅u2rEu�(H��1�%�8��6��=I�b�mg��v�n[�ʌ�<
���C�|�Tsu����C���~��Ƨpw���2K����C�~)U�`�HY�0�{�{y���w)�n��V�U���\�
�W��p�IE��-�����U�%7��o#�d%���$A��Z��/�����2�C��␱%����5�^��.8��HE7�.��4�J(�*�^�N�Tuk�~�s΍�(���a.�U7���4���I���U-��q㓬:S����j��E�8�xʌX��;�΀u-��i�$��H���X���+:si���᝷��p�� ��b=k�!�uj�{��1y\B�L��a�c���n���u0w9�@N�#����A� ˛��;z��qtj�f0�|zXQ�K�F�?�+������T��	�֯nM���2��c�=�,$�>��?�����j��䇳K٨���3u݁R�v*�E�w�r�Wg_��A9�7��5�Z�����7u�� @v�z�.Ƨ� ���F�gq�Y�E���G=�G����9d���R9���Gy㲰L��&��� ��*�Y�"Y�ky�J
�F"}���9R���F#�gc�����*�f�VD�7Wc47
m�����5�(E���;D��U�1�#Ъ�!�0��fZD_��O�|�����F.��)��I��n�e��쾖��'�hM����\��������}�8��(j]߄��oT�U��Y]�.����p|�Ly�'�cp9�̟�PL�k-�{�L���WEf��w���X-/����[��] .�+;je"�MjRΏp-˖x���ą��S�L$���!�u)�Y�n:b�
Ӑ^���a�Be�O>e&�6�Mz�3X��B� ��
W-�h�ʭ<��M* ��'��x2���I�i;:LKm�oa����7��%�V���y׾6��{�z�	Ԇ���Q��>R�	P��]*ؙ�(�_���9��5Ng��#��R�)o\"=e7���@���=��#Zږ�z�h�R��.ENz�$%8��nz�nv@`��}��}DTa���Wp���=��GW��֢>D��Y�,������������gr��P
k�V��z	�"�O����a�f"�o��ٿ�q%�D#�SwhcީBP	0������bF��o�p�^���Pk]x��*I���f3��h��T:r��D�����K�3fܶ͠�x���ʲн^�R�Sٌ \���Tf��ꉫ���+���A@EtX��l��#���fN#@Q��?�-=p.�FuFM�ls/b�5��v�U�<���f�T�3��	�T��8��m��,�-k��c����x\�K<q��W��F*�M���ԝ%��`PDZ�������Lb=�c'Yq������@cb��������_˴n_ Q��'Ō��c��t۲j}�,���ޫQYHDX��X5�n�qU*e�Չ�,XRX�a����x�=k�.!`������b8m�1MeA��_OMDU0�
.�qȅ�Kɺ��Ƴ�V505Z�� �/`KȖ�D!��s�]�V�{4�kX���)����!��9"�'�OPa ĩJ��;��̴�-����l�[~bZbM���7֖kkGSD}�As���KP}@���S���q�z�P���,���ĶHH�-cΒe`	�E�ɭ����o0���pF$�Ii�G[zd����bLP���D��mԄplD��Y�C���q��]���\ �(�{�K�¹��}�ƵQ��(��ք@����)j0L����|y���7�+N;�~R�/��_�Sp��u]+J��G[�IE��d8X������v4̿���'�W��P�p�g{�j4�ڡ��x����ej��cV샩I��ѐ��"�%J��ip�zgU4��'�����_^RQK�ﯰ����K��]�B뗿To�\oB�6�����'ކ4q���p{-тj)�̑���5�oȠb|�@f��qVD7)�=w�
	Հ����l����3^����R�nv�4B�@�< *�}�����Kܷ�c8��uN�3���w�ӡ�����`(c4�ia|��&}.����!>K e5�^�{�*�����O������yS������p�N�R�S��I�VR�f �SmF}���>��?���I�l�}�x@�MD������o�ma'����R�qS^�yN��!&�����i��A�W�&	��m���IY��  Io:�Qe��,t\R5�3�$(GV_� �9����j�����C��_��s��1�f��4���`C��Y�|p�0��?�Ca��G߸�)�i�����<��_�vU�[Ӻj
�%�V������^��>��俢]>���C��4 �/��T~JEDp8��I`�����D11�[%�l^0�΄Oԃ� ɲ�(����"#[~�"Dڨ~ޗg�x�� �,KŎq�'����Yq�~�cq�B��x� �&fbJ�H`MJ�DvGr�2\.CF�^p$��n���x^�I�#�������%փ�I=�B`X��c�{�^5b���,g1S����nM�H� hO�!r	y�p�rɯ"�t�s:�}vb����y��W݉�ڌ��>�e��Q`�^W͚�%��F��X,X����n���������B
�����2�Jss&�]�[{4�Iz��'b��^�u�-��B�ޯ2ֆJy
NY�o|�s��?;7Xiqk3���SFPc�?�G㉼�@z�i��$���C!�\������0��̊��n/=X3qG^�&�T�S �r\�ק��1q��� q���@E���/zw��tE��(�~P����ˌ~oH�x�]��fS�6���C���"�Z&�<������t'�ni�RG,?=v_��u�aA�[���[-�ڞ�m$�#>�cA�mW���1S�M��<T#0X�_�z;�T�/C2�@6�P}+���!���F�hG-{�V�T�p�۴5`t�5͑��1�Q�b3H��O�*Q�	93�y�O���@�=0�7;4����i���Cq��/* "�& vC�?���J�V7 ���>l�(t�r��L��m��i�Z�ӊ�����?v��N�%����4�1Z�#���OE�*��%W%�3]m����t�-گP�����p��1G�pl4��" M?��bG:��C|{�&���K�߇_r�>qÖ�(MR
��Lɣ[��e�-���'�#bս�/O��RÝL�BU�jP�p�}iS�q�,W�C�0'���L�Y����4�O���7����7�0!:��hcl>��r-��â$��Y�2Li?����#H�/�� Y�#�vX���'G�]FSCq}�v]B���z���'��M�3\�^�L�04'Ə�������p��]Q�.QNT�u*�OA�f��������G/R%ܯ���M�dp�$� ����9G�GwH�F`0brY9"=��!5�K�n�r��o֏��������`�^j��][S#��뮾f���"e�!�Uj�/�t��-0K���r��������>���A�mlqQ9�W~�z��21&��beVrDT9�uVP��0
Y�O���U6�6��ȹ����!�ፑ��z:�����6o��1�Z���й�8Y4��XA�U�NoA�����xC�N2Q�
<�2x#��ܚ6"�;ѿ-��vz�w:�=xT�ɦ����Qa�aJ �.�zXL~��Ƌ�z���p�0Ȥ�X��t���:����E��{��6HoA����<bl��W@��"��t�����ͫ(�s�A����y�k�w4�׹��� ��t4w�F�J6���=8[��l��4�f��Od���G���^%a%9��s++��k����D|�_+b�ř�#æd%dn�K㔄MEdP���q% H֌�ο|=6{�0B��<�+�Q:2?�h��V߂[	'�'F5�4��y���F{B\�P��"9���]�ih\���ҐM�[�Л�'���Ѓ��uJ�Z0
���q�_!�R��-��f;��E02�|�.����+\��u'`����d�m٣M�b�GU!��~�;�v��AT�����IP�+q%��j'����?C&l�O��ɂӾCA�r#ԟ�B�p�*��_@�����bL��ߢ�.���i����a�啈��;���L11�t��MDޥ"(C����wx��|�$�퇅E�@ƌ�o�z0R'd<�9'�y�NR-��S��^��9\�w�>v�^�h�'z�♛I^���e�@`�*~�˺%������;��^߾κ��5����ox�Gg�О�A����n���^��RP�'�T˛�ʑA_��1Ĥ���!u�읫���4˸a��,>�,��6�r�CA�sa��6z��T&�ӇN�+u^�{���^�'BJ-O$]����1�D~G�p&�P2��B�`�''�v\���:�^i��ޑ^��ߡve�9�G(�,c�n#�vU	��xd�T� �$`y���7�������,�+��[��ǩ�+\;���߉L�Ja gh9Z�#��MԬK1�2��������P�wVQ1\h��r��W
Z�k:[N�`��E�j�}����h_�O4>v��g�t�d�G���(Pƃ�{���%s%�,冀9Aԇ��+$u�����;|*��{?R�I�R�+�e��Dh���]�.�����䚔,�td���J��6c�w�a>{l��!-a�}����>X.v��	�#���H ��۷Q%]�����| D���֨q��0&�ג���e�8W�Z߀:��[�@8/��P�b���˷bT&r1��#��;�u�z�@�g�F��k�����J�����P����:TG��̗��4G"��j� � sߺ��[��]��W/xJ�qD��1�]u������x�˶w���w�jӷ�;.���@
�YD��=�&M>�U��N������7��#I�����kc�c��� ���)�υ9�ؕU��N��(�:���Ld;e�Vp���*�$xD9P��8�>Fl$Q��	M�Uo��]b����d���詵�A��dޫ7���V��L����g�~� L!X���1ebv�ۃ+22�����v�;�R��!?�"��'��l�nH����o�ۧ*���<���O,�q���Q��f���c�����#�~�k;�ԁ������H\p� v��^���8*��´V���]Bz9�5�V`�n/T]��Q'V��@��l;�#���r����B�֏�c�!�IA'�� �hxSl�xpӬYDh��͔�qǛ�V9�à;��ͯ�G���t�ƵT�_0#��*�ʁ�v]��M�żvS��^���55#D���S�X�����+E]΋4o5CR�v��,S���D[g�[,b�����
(t߫�����k�	�z;L(�����
��A�K�+�If��NE�K��	��8e���[6�����'ZYw���D�gd�M�n��#�8�@MVJZ4ɭi�Ui���,��>���_Ɗ���־����k8K���|��
�Z��<��������1�﹵uuR{.�N��>i�3��$�S���k�l{��|���E_��}�=�ї(X.��1����ʓ�M�cf������6�Ʃ�q.����<�C�q�$��@~���ƾ1މU�>#[���WD8r���rn�$�x9K����)�$؇�j=`Q���U�'�	S���O|����|`$�θk!NS��/�<	{���B��j��Y� {�ł�N�`O7Ǩ䊷��$��0 7��wL���i�i�
2i�U*�zAB=p�Y9�$��I�A��������p/=8Lؼx��\�F �pd�w;9=s���U��r�"�\�0g��أ�/���l���1��/��nܱ�$sK�2�ӮgDN�#�r6��m�ƈVb�S�Ep1�L���_8y!���]�7�({y���P$�q^�~Z5k��x���k����Qs*œ\絷�?}�;��@����-�:�erN����b��)�ar��iX�v�c���e��YM��������$�}�o݉�Z��@�l`���+�K�B2�$-�LDM�UV�0��.�Wco�N�� ӗ�5��h}��Li7�f���! �`I��u�������C4� �jA�T�"2�