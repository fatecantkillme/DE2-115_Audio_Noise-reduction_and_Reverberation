��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@��R"+�"v.�}�A�`"�?�B`�{M-4�΃i�֖8�65ת9�֯�j�[��Z6ܔ��NhK�����/-�� �BO�EE��b^����j�ǹ���^q����l��^�"8qZ�q�����Q ax��y��`�T	"���T�Ѹ����ȁ>T�1-0�Z�h����_��̸Lg9ٲ��CM�8~X��������-R75��\�F�pլ�u���ny�ˋ����Lߩ'ŐQ�����=�וW�}ٳ��� ������]׺�V�o��D����d ��Hɫ�����r���`����lA���V'Ρ��"�!+?�:@v�Ț��v�}j��7�ZD�F�	�R �Mo�&,/��SB�᳔s�ڿx@�U΋s_6U�6>{��#�C>@�;��1�d�����+
��s�A�ۗ�	����l>��H|V�L�8�~�e,��b	���`�!vITA�_��$�O"������qQX@<b��ѵ��d�)�cjJKt�-���bO�-\�e�Z�>Ö3��}1d뛭?�MC
�t�����zr�Z��p��	�D!�S�?K�Wё��~��z�_,���?�f*�������S�����%M�P� $T���:.��̓r�!��o�mk�U�J����Taa.��yZK,
'T����pڃ��'�,ʌ���L��"m�P�ё�T6]�j��xZ��̀�q����\A�����P����:���I�f�Lx1�}���Ɨm�`{��זv y�W��3�6v^���jZ�}5�̞�-R?k.��0�������.�b@�
y�'�P��O҇C.��X��hp����۬�J��孨����D�{�V����s�ۉ��I�KO���g?ݦ�'��;�]�ߟ��Z��W)J,Bޟ$���SK	�x	G�ģ�kx�����{U��Vh���ѧ�g
����zm�'��<vdH���|�J	��y�h�N2qu��ʗ�ڍ#2Qr�Al�_��:m��Kڊ����p)���Ŗ�x�e��}܅�(	H*�s!�D�hK�	��mѝS<v�PB~�Jǧ����7@F�"ִeN��>!%�QH�w@ș�Ҽ��G>9��u��r,�Q%�e̶�H~��u��Hك���x�O1�(�gRQ�<�91�"%T�lA3�����
���䳦��*��`k[��oz���h�K��Cx{���^b>҉�� I��)�?In�d�gA�W-os���Է�c�G�a�Ǧ%6�:,����^�>q�dR��T3�t8�Z� �Id�h�z�Nr�nq
�����w�]_�Ꮝ(���<7kW1ΙŪ,
�0QzH(/��^�����IeE�@��l�*����r9Q�����G�Yp��(>�)tYy�NnE�ߖ�e$��T������;�i�9��$O�WG�Q���DQPK��.-r��z��ߢ��r��>�vM1�G�"�C�o ����K��/ts�5&�vM����*��=Zo�ʉ:��^�z�O�"��A����p�?q��V)UO��a5:ɰ}\��uݗ���?�I~`*��O6"�&��y;���=������l��R������|�=bڜ�=O�s�O�f�b똀����>���X-hO�RA�X蓮fs���WQI� !muFGԃO�H݅�����c�=�)8�:{��{�QS~�r!���K��N���Jg2Ph��*�b�I�:�ΜX>��ϵ�QŻO�lG`р��:.t��o"�Nh���-Ђ_�,GK�aL@��	�ɱ�;���e� �v�ʻu{���)5����5��+�s��t ��H����z��4�=���5�r�0P�8�4Tw\抧�;��v���(��&�u+��ٛP��T
`jP+�p�$v���Et	q:a/l(��ę ���S��*��MLh�����T���[��h&}"rh/.�4�,�U�G�,P� �݊ϼ_';\Xt���֦4�N��y���02�������<���G)�R�'�g����L�X'��;xD(^sS�é��߷�4r1��3���0����8�|�[�\\�2�H�s	yy�N^k׳�v���o����q��]>�Aяf��h2��&Kŀ/ƣ��]�\gjks�:a����Mo]Zʪ]����6�y�ƍ18���m��� `ʁ��W�#gT���2r����7Z�O0}z��t�?ܹE�O��]Y�*��|��C�O}d)�M3#<�����M+C�[�*\���.�Oz�I1n���}}��S�_��6��-�wٸ��9��p��}�][���A�g�4�Q|d{�A5�|��8�F/a9s��F>��h2	L/eE�$���w`_��8������آ��D�	��bօ�K��&v�����&!����Q)?��HJl�M	���-�ev���A��jq/���%mX�/�@��2M�S�1�C�V�K�;d���U�������m���s��t�\ߟ�_��1	�Uw��=Jb������MUвE�p駶��"�V���#}�Xd����3��o���J���Q�jUp^#�f��9��#*�J�ux5��f˙'�1��|y�. \���<4ʐ�,m�w���`�5��%��[��$��[��N�����hM�4h��c<y_�Zq�)�Iso��,0����H�ljv��{s��-�gutb��Sq�4x�
�^�����=[���>��J��C��,��41��Yq����J'�@[� ���V~ek��qK}< h���JR0��O��������E5�s�&I]nO�mQ5rO��e7n�N��V���C��J��`J�P�˴b��귥�'�^�Ů:���R�!�~���M	�͌�Ԭ���P:���K=��XǕ �*G(;�·
b�g��H�G.�@Lw����Ӛ �k�����J���vpq�$&B�M�z���?į<2��v	@��Y}D��p�AG̕"Il	*{�i�C�J��9�v���/ԈU���"����0�b.� �D ���4X�r�ZS�V��J�Ⱥ�T,���>��䴼$�#�[�ϻPs������E�%0p���*�`��;���iS�C�9R!�r�߾�^u�ƨ��/]�Ĩ�rT�Cc��u�{jWe�k��| u�.�m�ƿ@Fb;�ɧ��e�n�?Bv�_􂩦i/l1[���A���Q��%�&�̿���=B�y���:�� ���s�e����[�l� �KMZJ�lC_�؟��6�$��;��m�q�[��V��x��+����@.�gD�K��z���WI`��+�3�`ŀ#������xH�Bb����n�����B-Y-��ʤ��0�xעӗ���z.���j�⿑�z�N��-w��Sؕr�H�U�q&���;@}[�9�^]#�Q%6�L�r��a'��/?Y���j���p-\�,f!BT1x@��''ް�`ē���{���X�P����>v�=�1�˩���q֗����&!�4��i�x��\O��"e=Ȯ��:{�2붐;\��}j��^Ƿ�4��W2윀�y<�7|�ٞ�y�I��8h��������1f^�MN�ffGH[P%����ˀ�W� (J5no��5�&\���^��:�7h�!�K��2��F�=�Z��=�m�F�AU,?ly��2��x�ͦ2bJ�t�1%�b&�a��#^^0�v�
P*4�����qFU9���究�����rJ%�?�VkE�&��w^����\��z+ϲLX�1tI:{�i��8��l�dBb-����9!c�$an7&�
�Bt�r��q?ي^�J���CA��"d��_Λ�qb�M�b����yx,�B�gm��}G�@lj����*�D���q>�+P7?:�H���|�����^�������y�Dh���6���$��m��[D���:�Ko4;m��Ncu����#�0);���_�a�J��PIqX�$Ee���kr��<k����
u���!Z�	�d�jm'��m��l�Z���I�%E��x��t�P��IJ�JY_3��"�ڦ�QD�UJ�����$�/��9�nyJB'��j�����7�>I*nIk�#�I@V-Zx{�c��}KoMg�Q�����V�/8��,���)�m:��h����&�x���o��$��\�ײ,��/�@�a�����z�ڽ(c������K!�i���* Yo=o�Cq�U�K���u�Y�rq����"tÂ��3�Tn�A쒚)�����d�5O߫�2���n⹧��Db;�щRW�"�e��q���
�u�̗sد�}_���,ƨ�}�~���d3��Fk�6���T���D6��)��=!��o�ɲpӚ�ۡcd�]Ʒ��`��}#E�Kt��,�~�A/�e�ycG(R֟�"^���`��7/��t���z�k7w^r�	Z)h�**ե�΍� �\�ov��_���"�P}b���eo��9�(��+ ��v�lN��h6��k���B,�� 1Q��G����h?�%������?Z�qg��v8�bL'&B�$��	������m:,>��o��YX�+Q�
 �'�!�E���{$�9���b7v�7�]�피#�DL����������ޖ�&om�rH&W q�~�I�v�1I���@�S�i���7a#�g��!l�|���:�1�B������/�� ��J�P�Oo i�*UV�7_��Z���7�O���T1]�&?��WVa��{��c�%�����>I�	vc>��u�3��.5�K�C<��(��/DyI�����8K�zū��D�t��h�#~��g�U��9�d�w�oDlUP���Z���,�Zb&!�.#��$�GpJ���x�� �D�|���壔`4��� �K�M]���v+�D�	�iQ��b�ҘHL�仮�({�`�2}�3WV����>K����Ky?�$mb��*BN�	ӵB�"��s�s��駝��N�D�(����/]�5�n	���-E��:���������9�(^=}m���:G#v��0D�$W��*K�/i��8�c~V�mk)�ŜuUF�e��j�oC�����j��<"�^
��/�Y�M�-�$��r;+7���ٽ���c���O��&8.�Ȃ�����O:ӍG�	OQ���v�Yοrs"L;��ht�\9�5�S�dd�5�\�&qN�A���I���� �nwF�d�N�|����*�`��P��6T\����Q�O)O�idi�i��엺y��G�~3;s&��cML��'iB�% %����5}~�vM	�����<����3X]�F�<�X���QC����,<b�V��n6�.��#��pvlR�b�o�ש1Y��I�͹�Q"(��X�ks9��c��S�$���4�#��Ul��b�3k����2����$�)�ٝ˴�K��ɠ���~+ڮV�i�z�qKEr{-�z1��>���2����-�F�&�)�jOU��i��2"�e�BpCWf�.��xr���[Q[$,�4��u�v�{�r��#�=o{0����@!G�I�B|�U7��������'��kd�H^�l��Y��˩(����a��a#�}�Fp�����{2�?}��2���k,2�_V|))s��+��g,��R�
2����V	%X��W��E�Ҕo��w]G���|�3��
@�z�5N��4�1Ww�C�+��R0:7ׯ�ʆ�b|�j�a��VJ����tCV��/�-�P
^��=�$2�v��w����}��|�~?/<���C�0B�c���,��R�~� �����.^OJ�_��"@ͣs���TM`�~���$쮎7έ4����2ӱ���:
`V�x�U ������b�����6Q��̈́͢�[+޴MTG6�[��(� �6�I�uE�9����3plU�(
NS�67:�skpqgib.��|�#&Wm�Z!^��������HE�y5S1���}]/�yʘ���Op�B"��Br%�K�!UHl'#����c��κ4H���[��:�ȦR���K{Vv�[U�v�'��c7�\E���Q��o���^�^��f�׸��
a(�^�)�~���kq�gh���6p �X��*)Ft��i��� f��l'$���e�"����%��������9��^��}�R|���Ϲsa$8�\se�0f��L%��6_�sɺZ7��(Z���I*h�c��Ӭ�麋��KBk����� �i���'@-+{UΌ�����cL�"H���iD�fd�~(Ȁ��T4���j�Qf����B�r�c�`�W+zR���S0}Oڌq&^��)�.��FFSW�������TS�l�Í�7}�Ơ*mvJtP椿�e�\���L�G;���c_ \�[=�$4#�56�@u:nE=�v0�K$DjL�����w�H�W�����hp��֑U��[���D4Cs����M�Z���O)��2,��G��S���c���o�Q,�J8�	��pg�5�e��<S�������j'Vc��T�N�LiP���t�tY��ڨ��)��;)�&P�R��x�3�\j8����Er/s,Ϥ;>3䊪��P`�A�
���x������N���a}���A}RFH������'I��O��%(o=��!i����A�����sAFư@pr׿sv�M����1��Z�7t�u��*<w2�6�.lJp���d%�ޣ�f��ne�Յ��p�m�v���W���jfo��Y-�*���+I&G)�b"Cr�|���m|IVS8�y��@�U�icͺ�)]�^���������-8x?{:Tzr86���9���;&�ev�?Ǚ����vE9�q�]�o��B�]�?����
�0�d��V��ڭ�5��,(y�ч��6��o+�'�m;�h��ГH!`8˗d�R��s�q��7d
K��<��e����pp0��qѣ'�;x��i��`���ڂn��z�R�/É/�\]��� V�QnK���	�U�Lx�+,�v[h��@&iwq���Rz�+}W$�C�n#��W�ɋ0�|XI0�?�~��CHҰ2/��u���Ԁ��&3%_%\(W��)]K���&	�����]��*3248�,�|6ް�(5x|X��P���[;i]�Ã�|u�#���N"i�-�E_��Q-"\9��C'>�@��H_F���ɔ��0�p:���Ƅ� �3���t�h[������u����n�S��.���@
�zF����&F`��ZR��K����(Σs��%R�!�9 �\}y�Uu6ؗ�k�|0�uO��6�v����a,;{��#[�Hۂ�P��i�W�v�9uq�qu�F�y��d�"�F��Kqg��v���L��l���z�a��=L�-Ox�Op�31$�V3��Y T6`�������E`Bl
�d�{�`C4�؇s}ͼ�b� ?�w�J��r03���N�9F�L�MJ*�q 5O���ы�+CJ=�P�
'�C�ڍ`���5\@Ӌ:��|�Ą��Bђw~�Hw���iO �.�I7����Qj�S�?- ��߄�y�:�[���C]�)�b�H�Cm0
�Dؓ��.k���V}�����B��>�n5")���2���U��c��9��&��U���@<�v'��U����K"ƃGk�lLJۢ݉��S�͹����J�Q�'x�����?ֳXq�R/�jqU��#BuO��Ŏ� ��:��VZViB�e1}�D��꣕gʷ&���	F�q����d���1#V���I0�/T�s��gd���>���t�GYMEJ{&d��=%3�C��,R3:E�Β�rh&X!~H��������i1��f�O�f$-R�����	:זb�4#�9�r�rWG,��S�h-$�8�����s��<�; �	B�u�_����Ћ�ҧ���7��%0r4:m�4�`d�QkHQ�/1]��d��U-2�>,�zam�Y؉���:~XG6�S�Ӆ~Jy������j��ZkV�c�z�
�'��X�_*{�֎�h1�-�Lˊ��Q?Uc٨��	B*���i��%֣˼z��h�B° �O~�$Cा�hZzx��~$Ҝ%"}[	|�зϪh����tQv��#'�����~�Y:!-�ʏ:����3{�� �o�}�)�I}h�}4�X������X����]�sP��'3��k�]���i�%��X�mh�
�`����
f���잽�/���9f����Yt)�`e��B2D�"*���X�5�ᾮb��AQ�gK�z�z_u�x"-�C���1E-\���x8/���Q �v����I��m��/cE!�1Lt�rE���J-iq��'y�uM����"�?��t8kQ�"@��|��LzFY7u�e�����0s�8����E����4X��5�x3�<֖�JG�VW�uQ9����K��2	�KD@d%!@���\�O������`-�J��lV�q���^�n���h��#�GK?Ǿ�4��-*��V�@��*b"��ǯ'��r��[���<����e���;���!2������s�%���
�y.�+��R�cA�ۅ���L�>�����S��ݮ���^ً�;��L1`���S���.��P1D\=��@�=�tz3R�PT�}��	 	�ŉ�y��W���#Dq"n�b:�r֙���2��ذl�)�ģ~2z��+��u��{�UB�y:�1�O4�����or�YO��k����w�9	BH���B�S�.��S�?���V��Ȋ��^�|x峏��(V�p�텚#h	��`}�S<pк<��n(��PZM�9�����Z�B��wԃ��4�x��c��aE���Y���.0���)�8�kQͅ��2
����5]�+C��-Q�\4�kt�׺\P.i��xr�Q������a�)x�y��応}�p%��4&؄z�C�C
:���I�������q���jѨ�r}DrO��[�=��OTF=b7�|8�u2�{j�
�;���v�Hg��FI�Y��0j,��v8�����[�-� |v@U�������9~ʺ�Q�5
ù4hU��7����Y7o��y��'���.���f�R��WY�.l0��nڔ��?P���³f��:#$	E*j���񺳛s�"����^x��.�ɒ���$�8�"썡."c!֛{�e0p�凨�2��+���~�)ќ~�?�n>�߽ �TKX��T�#�u+[1C��/Z��L��&�1�^��Z��k������M����˕p{�w�<)yJ$��|��ɭ�PB�2W�7>�����>�6ّ�����%8�́]�%��QR�;]�_��;'�Dʯy�u:�6�D�\Q��%ٷ�ܧf.$�^��2���##g�ތKs��*�y���*�����},���c�*)=ZqoV� D�&��@��IWOa�&^���Eg����*F+�p��%iE����'��d��2�*,�^g�%V۬�[�[ԞR�mQ�����j�ݑ����OX��;�0��V=�T�*:V����Eȓ�l�#!\���y�Qév�ů�	�ړ�E�$u��Y_+?��S�����S��9�B�=�s��}{�$��og��R�"�k�3ݧ�� ��!0��>��₨z�ǢV�Y������L4K�������V/O�Z��a
���:$.�-�a�M�x�OQ�`E�+��q�ɂ���k&�������505�%��4Yb7�"��ٮ�q���~s�x_�<z��i��=kT�nl�Ҳ5�Rlmb^��SuBy��i2��+$�L.����'�
�lH���
v�(��^���d+�Qn��)rκq�'U;���D�d�كY�X��Yh�}db�ٷn�R�:7�R�+����^x�o�Ç��QD��R�_'uK>�x ŷ��e����uo�az�˖;��))=+,#����'{%8�6�����*�5 ��4�sOI��lW��`d���ۋ� �j3�T2k�+q���R����{A>؏�MC�]� E��a��9�ڏ� !w��,5`�T�':C9M����+�!V�o�PE����H=��5�"��Ȳ,�F�_��4��O�b<5w��1ǡ�k����}W�?��C��38��y���ܸ�np��}�ף-�T�S������u�In~���;�h�^tI�Y�3�N��N��L�A�?��O\s���#>����\P�2?�&��E��v�0,�f���@jP6Uaܳk����xX��of�#$ Ɋ���>��Z�,*k�b��O�������N�v	���d��r���@�qty��]6��{�l�~�4��A6�5��_��Y����gf�ޯo�'���L��)^�|��#�װ� �G�ё.m�f%bM�OuA�v/$�p(��R̪�m��om�|��u�j%��SU�fŅ���-P�w�C���S4��O]���=^c<����οH^N	T��
T�������.�8�u�n!���e���	a+Jq��s��P����{�f-E�_\��R�P�
{�®*�N�1�R�8�JU�`��5D�x��ϟ�:�k������}��a�����)�O�����jE��m?�6�����)��ßK�G��s3��MUE�ôW;��Mp)�&Hq+RV4e�a��ܵ�j@ľ~}��뼤��'V�I�-): �'��"�,���Ip@C\�՘�mS�VO� 8Sg%��e��&Y"��(�����,� �Z�[��8i)��?�eo�q�����&Ӝ�p;�ʾom��%]����ܹ��<-����d��x�(F��y;;�M�_��JGK:���A�C�,H-�@F�@i�NiLQ����'��B��CbFLR\���9�;(��m͹�t�ps7�*G�ϵ*<����{ң��ĢY�u�Oo�X@݄{�/G� 6�`��!��Y)9��½�*c��٪ީ��Yl:;��'KY�poKo�uQ���A,���>RKU�����t�j�Q�����%�s�N���OFSXc@�f����8��$�<{����i��s�a���Y�=4O~��/z���z}U���Ë���`�ϻ�U(��S�o>n�C��>Ev ����T��w��	�#�F���T^.ZO"�wl>|8����y	}��b���yb�X�o�	�A�>/�`��n��I��;��兮A֔�/?r�;���@�B+;�|�v��	o݊�Y�T��Ip��H�Y��U]�����$��u��^�sO�y�?K$7�M�-P��F$>{�~��Y�L�������q2AO%"�F��j^z� �K㐔`�����m����������FS-sG��$�ɛ�	����O+QA̛,��U��P�)���=)ł�. J�{R��Eo�������`��@�{?�n���3�M���lwj�,E�g���M�Pj*�ǜk(9�w��h��U��0���&�2lB��y���+��k>=HX�������o��E�զV�\A�$�h���3� �mo����b�x�F;���`3��z��o�2谴����ô��*N�B���[�Jϸ�))��:"0k��qEn�Eu�\��m}\6ޒ�D�ܱ��:�o�5��8e^=b�u�X���I#� �Vy��8#N��A$L��H%/u*�:�v���V'�d�dȷ��8�z����X�mw7`��Jh$�}H�^@��}篏�W��7�	����D�\r�!ؑ�g�z5�e'����1g�]����]
 `Zfߪ��߶9xd$�x�@�g��R��QAb����1��
2�Z$JZ�\h/�S8� �ݝ�P�����bƠ�&��� �#��[rPw#��v��`q��D�o_��� �k��n/�y��S�=�?^x߱�3��c�7�7��>�a�,���F���oo�p͛b2Tn��E�Η�A��P�ǵ��h�.��z���F�*W�=T�h��ߦθi�� 3��	!��$�����]�Lۀ��Vd�"ơ&�TVªء�����s�;v
�ů0�'4���#��͂�ϡ�j5�ewc=����D��)�=~&aPŇ6Z5zh��>�	
hv^bG1#x��NiC�\�&գ��¹�hts�;�5�AH�������`Jn�~i�G��o⢍@ALO��S���*c�\d�1k�"�l�c4hFNq(7|Ӳ�Pst�y&�X��)6o��X��Ɯ#��'��GQ?������V����X$��{{�<�V{U�Nj�@8$�Y�ifhN��|�'�&8G�������t�1�u,u(G�af<���ߞ��F��<wI��Y��p��|؟{s�nW�y`#(�|;���J]>�J}/�]���@D��#g������l1񙟠�teVt��mԔ��b��]���J!��� ;�ŬPf� E��ZG5m�"�X�a�����G����*^�lى[�烒�I����IQՠ�ڢ�|x����B�/?z��a"��u\����h��c܅T���{��F/�y�5�)����\�V� J���PMXX3�L�"�/���brx��ACmv̿(�H��P�J��ҍy�VS����]V!_ә�$` �%�Q�T���=s/���T�4<�V�")azj�ms��hc-?-�d���R.���Ffw�m *��_9�%�?�!&� 07�j�&�gT���zNb�a�(S���%*O��9FV)�|�7L�y~<3( Ɩ3o
�r<&�0�eN���I�ߊa������p&�?��I�*r�:��*�E��g�Q�x�
��Z�� .©ό9��?x(h��p��8��N�mǜ+a��򿙁}�`	��RkL򢛗�6�T�/��j|�,��ǈWF�f���w���3�o���<����0�>|T(���'Ї}�lR�)T1 �\����Hxv���pő0p�hY/��4�J$�²�5����[�)y&�������g��䗖�!Q��1�g�y��O�N���@2c��PO��镅����)�2}����X|��yeŘ�\;a(�DԊ$���(�Z��-�y���{���=��ƴ����w�XO��4�cU:��� �?l��5���	<�y�OM�a"�z��/5i��3���_���qG`d��+�c�Z���N�����/���34u�
����K�E��>�X������[�|�fb>PoC���J���tuFMe`��O�k!�1��vQ�ޞ�G17�0���ŗ+�T�r�U/é�-Z�7�Br��Dsz*��8r�
�\tR
�+D���3J���� ��C��9ݘ8�|W˪���u'4PԨ{���I<)Uc:�܇p�̴i��و�cdw:S]c��IZ"
�I(�o_"���ў���-�I��k2�w�%�-����vu����y�#MQx��hl+�<�g=�\��*^�f\]��໙��>�2�%�1T���vK�`�����N��H���۔��fxw�
ۈBo���Y�S_�ׂ����1��	��c�D� lk��2�sN���ǰ�����cN����_bI�`L�<ܙ�|�2s������Ce� 
;v��`yO=aMϺI��ϻȊ��yWז���h���2�G^d�xK�A`VB���;g�0��0��h$;�����(T
�B��іR��u*j�$$��Os�o�0='҅����+�;�\�^iL���y������?�vbz�#����K`�C/�
s��x8K�}ZX, k(��d��x�>���4rRw&M��E���B*o��Z�.���s �Xx��q&��2<�N<�3�8%D��<�-�{���MFG`n�d_z�.��
b'�4Zh���������:��Q=7��Ʀ�i��s?X�H4͋2����A�~wI)8(�3�Q���4M�P9�Ph��9:8����e��K���|)�)3�|��f\���	E�X(��8�b��ғZ˅�n��g����k�F��%�t��uK`6
���n=�̳�>"u�������j��@��.䇶-��";޼����1�YH��	��?�@c�N�J7�^Jo/�á������Y��z���F� ���J��'���3U����%x��f��:gQ�᜜�
���Ƽ�X���1����"�]n�8�S�+�f[ȏ���,��ȯ�հ��ĆJ/@���Y����$�\������s8�
��.��7
����H'EB��A� ��r%zr>��%�H�e�6�Ny&��>G�*�	��t�Ȧ�r�N��V�5ʪ���@F6�-�<Z��1�<����)�c��J��r;SP`���eP�"彏�~��6i�2�R�_u�a�L9%�r�݄���m�m��1xN�I���(�gee�4!`no\�
�
�1K~s���x  ��jO!��щ�>ٯ�c醃��qNMJ�N�8x��/D��f~w�����4<W���U(N��V�Lsuh^n���k	���������	|`
���	4��AZ9�T�{�#m�r��[�:l&������Kף�]��}�Ys9R��#�f�T]��8��^Ɵi��@,�����Y ��|%�͙���c�W�u��"�PN�d�$�<� "5�o�\94/A��4�D�%%<�W�Eb�F�b4��]@�`f����qF濨Њ���F�����y�cn���N"^{��*Vt���p���GL�e#�t�we.`.�ٙ�9�� �l��(�tL:��Fw{/��֧^�Q�-���Z6|܌�L0~)�)�
7��I�$4��p��r�!k�J��-��;ü��_%���D�e9	�?i���0 �T8�CL.�(0��)x��ճk(ı�Y�<��dӪ��,\�5B�-a;�-�/�w�P5�v�3>���"�XPoV����EڙG�� �(~^��\��������Aq��Z�AB���i�ϩ֕�Uqz4����SS�Us��5�Rӟ���� V���U�Ò}��|*��fIY���E�������H�ñ����K�b���I�04Y��<H���o]�j��PXi{�u|В��i�D�%E�_��If�/���X&�<���I����œ�t_���ĞX�Q~���6�L��}�.&z���3���v^xJqG*e=��7���D(@8�0e���n��,�3\'�ب����N^JFyu��m�o$�nM�-�ę�/ߓ�����a]����u��}��
�Y��}�o޿T��)����?_{
��`m��(�ja��d�*�`�_S�W���)ꓝj�d�V[}��$st��6�i2ta~ڐ[�n\�L!�[G��VJsh2������V0��r�8���o��9�ūY.��J��þ]�.�%5�y�u.+He{ê��А�m%M��ޞ��9Z�)�R����9.)��]��I����c��!s���"��K
��D�	�;�����7h��@��V����ï�=Ȟ�i�-ka���U)��\�8x�m�r�M<�k'R�T��>�B �=�������.� ���fj��6��a'{��Yo��EJ>XS�7�pp���*[ �Ŕ9��0JٴC����'����e3)���V�����O�x*��A���H&�G[Qt�4��T>�s��a$2�h�'�3Dј'�����c��l%#�y��Wߍ�Տ�N&z>��&t_viSh�n�&��_�SqE���c�_����l�<o^��M}ޟ��<{�:U���	}¹Q���?�/��T�[N��V ��$�Y͆���6�W%^
b���ߋ,�������Gk͸ *���p�j�g�����HAݼ<)~'f��5,�'�@�l\�ʕ��Ư}�5�y�l(�}�=j��nvK��N��M����*>QK��s�-�Eto��1�J@�-�'
�{@j��.�^!��QG��\{���Z͝#}�2���U潆�N���!rb�C�d8���D:Q�����������a�>-��9*�Cc-���+@�*�f�&nn�,�L��~3=�=��Qi8����5�,�Lȗ^#h5�6����^�n�J!qP!�[EsK��>`F���Ryad��ʽ+=�Ɵ=P�Ô�"�_>|3����.@@?�ĥ�6G�]+�e�-}/k�JH��C,��,}A\����Ja��k��ﯲ�i�>b���� ��VG�Sn�uR�M:PD%��mO?<�G��6(��Ţ�#����0 �Q{���B���47���[�.~�~�H��e	�Y�(�t:5��P\�e�A\K�נ?QУ����H����}:�Z@��?�k�*���u�G80�F��X�O_A���lv����LZz��p(�B�N�}�������0n�|����sC��[�� � �E�mPu$������2W�y����V�:��ܰ_TR�<wOKX	N䱳�Ƹ`����d��m4&5K@s�bF���*� � �n��L�|�J��u$��`л3O�)��3)%��k~.��}�Ysr�3���|�>��E�f����W�]��٬���F��1��u���x�8V�ka�1���`�Pleg;�Mr�R�	*}g�KQ�����M�P����2�F8~���6Fx���p�%�rqs7���R��&��O��h�7"-�h(o2��Ì���+�� ���é'p^��k8�%�X���
�sP��7
.E���t�I���.�]�^�&��y�(c�b0����myȇF��2&�;D:c6d�c!�r84Z)�2Xba���4s��p��$bk���1�_@�+�f%t�7"�J&��w��uqO��">o��6�,4ݢ�s ��sf_X9���	�龚ֶ��%���~�jG鳱%�|\�P9�'�%��C?�ߤ_��b)ժv�7R���j��w�wmm���D�� o�P�f��"
�;�Re��������,�����c��\?��d��� yۉ��^��4����蘮�n��d�ѕ��ݐ����-1���|�w�+N�T�eA�~;�ϏT�����)�\��^�����t�3e��o�����Q����X5l�Z�	�N)�E��Y_�k��
���麬c����i[�t��~�Є��ǻ	C���R������Y/w�Ѣ��6��%��K�5�"}���k���e6����߯ߚ���L���[/���h5ok�CJ[X���F`���9�Y��i�.⽷6�ށ�P��I�O�E��|]�K],���_���b�°���Ҍy�qd��9�)��c��In��� ���1F���s�.P#=��N���`�Vg�;�O��g°�_.�� f� ��V[�&͋Fs}�W'�ȇw���6��o��C\���3���3�����hsZI�9�g/�{Q�R[5Եm���>7����Vڦ@�SZQ�Vw~\���)�i0�꽑�u>�  �*�x�4�׋��V|����/�z��/�"c��b����l|��="P9̍�\�����7��J�o`�yfj�-tz��L�o�M����R�#���y���J$gQ��S���u��3P���C����J́K����ɇK5�`����5��(U��[�)u��슬f��u������wܬ�o��A�Ieì���mP��3��>k��Т���p�δֆϦ\1��L��Ͷ�Q�"��ofW^KM���`���X����%S�q�Ǆ�:�W�9�%��c�?�����n��J�[��C��Y5�5x����%l��j�qwa��5��)zD~�g�6�V�o1J��lkK��f�d=9�
Sv�/ �W'����6�D^�^��fԋ5�X M35��݌�s1 kK�����V?!�bj�4�ο�1�+N<p�5J6o��$�k(��ȴm��w�^�&y����d���*����ȫ��>�{�KW��QB�˂c�IA���@V��,9H�G�́M�#������*��vy��1R���y榚+)�8���"�b`,�<%�<�PMI�Q�K-�o������T�������J�����I���m��O%��3Ǻ�W7��Jw�M��](�Ha�v�E�d��z���:����՝�ԏ�>��̋ie�y�(&��?�*�`C�1y.)�D�(�s�3z����e�S!J��[{ν�"J0�%���j��-	P�4t��1F5k�^H3�h�U�щ�@q��c�C-��x��'�;j�2o�Y��y��ê�NP�����Ϥ�eI�lﱜ��/��%P����/Á��;�SȥLC=0��$Axs�A:P���9�F?�x]�0�����7�*�����W�^��,Pk;�*��a�2�5�c����m�Q5-L玘�"��Q{�Ӌx�}[�	��=2-�y[�ҙ��9°y׭���dbre����~Ǌ��*�v*��Ƹ���᪁<
 ���C���Èd&��ᏍvU~�ݦ�a�������&��Dd�/�\���ض�Ic	�s��뾆Q��-v�?��r�xvͭ�;�p��{4��1+e�O���"�68�:�ea !B����K��WKs?�C�J� �Х�oF�j.9���5E�!*�D<+�I!�l"�M��ʿ��:UHˍ|�.gX���ςz��t��@��FO�Ht����o_�_o�H6�|;����B�h��j?��p偸��O*�|ҁ���Q�z��L'���2�d3a�Ԃ*�5��X�rRL���;� A��n�A9��H����,�*�jԾ/��=�h=���E�׸s�1񂾐}ޖCB��:u���?3+��|��$��9� ���F�
���nV��D��0�`U	'+:�A�����W�q�476U�O��P�0� Y!�+����7����s�6�pzlSٲ拡�P�{IL(g��;�RYf[U[x�9��O�q���-e�x^C�[�5k1\���Bm���k;�z�~^�F�|�N��ۨpSl8����Cu��d�/��Gܚ!K� ?wX��#�\v��6����.C�����f4�+��Ô"���kB`ԓ%4�������L�41R��É�gP��v.k�I� [HŌ)�I�]�@�Q�ѾX�I�o���G���썡�Χ�+� �&�-����n�ȧp�3�?�1�D���־��.�-+,=�#>!\:�l��X7<�;��Ha���gٯB�?j��C��C�_����ؠ��u�ep�-×l�z��M��ܷkң���Ϳ�V�IM��kHT�Q���"�����j�B1�ܻ�P �趯VKOx;~�Z�m�I���8~~�L��ilF��U߅��&²(l�����M�C��n 7�������n�q&AlU����7���.A�I�7��D�����O�$rHQ�y����v�П�?���5�b:ܯ�f�}B<��h�ߕF��5�[�0>d<�R.h]�9�ˣ��H��5�f,�� ����5���bXz�U��`b 1*�}�0���r;�wYw��%��&��U~2:���A�N�KF��TU���)T���k��� s�@Z���g��#�[lp.ER��(�_�^[c�7���.:�9�*�� �<���I8���ן� a�\���8.�U�5q���_\l�z�T���#��[�DO���[����!7᭯dޯk���=���@������"+��Y�##�����c�$�@���vF4�5����P�9�h��]U��R7$hFR�pn鸷z�DmE1_d�N����7f��o��vΡA�P+�CNS`=�c|����y���4�T�<EuT�"NJ�a��.<�tU%F�>�qG�����a4��6�o���b�a��<�xפ�_�U�)ߜl�X��h������	%�����������iNn�!n�ی??�=۝P�¨|Dcu��x���S6{��� �䐃>5�fi#�f�to�H�"*1�2˽@��<�9���|F��"�>kcǇ������.]q��Xܪ���������77h�3L��C<���Tn�4lh;eә~����='�N�S��=�S�P�Ƕ��Z��Yg|K^�FI��'F�~vY��N�F�r��W�H�.,�-o�,r��t_�K�jx(���Aeg���F$e�+�-j��ҹz��1�By�b���%��~�j��M���}b|΅�[5ùAz�z��쌬"m�r����$���ܧ�NW\�N� «�5ke��Ͷ��Cpt:#�"�A+A�V|_U���q���)4;=�&#Wb��:	r�ن���S�N��.�BhF"�E�`���dm��$��0l�*�0U�t��ĺ�������=�1^)4�>��o���|���"��3 �Y�H������P���� ;x���F�T֭����&cd��+�,��X�f�	('IQ�؎�_�U$��>`68��n�7���\�4�X��E6z3~-lD�������Π�����1����l�\��OT	�����s�Z8oQ��Dd�����]���ڛsT�(9<�޵6.�N���E�@x�$�����1k��j��0�rQ]�_�V���煭�pN���i����D�X���nx��yϤ���+v-�ƛ��h�s	&7�j�uJ�,��#ޱ��F\�*3�y&Xu+w�k���Kq�ﵚ�FJ�l�V��#o�W���8��e����Zb��b�* ;c4O�S�>�,�CPKC��wЁ�`��7��g��(�c]�µ�?�qs�Lk�s�EѺh�{E�a�e�ZL+.�Ï915�(�pӑ��JM)3�²�rm��t!b^��=��̮Į��g���9��@Dz:b5+����!���E4��gfjbi�'�3y�RZ�k�C�b9.1��9ZigOtGA_Jz��bI+�&���s�%=%
oe�2 
1����A��57�X��~�:T�p�˺����V-Y�@-��mDAF�)@���R��&��_�'�;fE.T���\�V�Ϧ����O�*����8�>�e �{��H��镟�GF����;c��;R��u$���&�&��2��:�)�����$>�S��="'���ǟ�&zZ�r�����rF�&���e�a �e�,���&c�Dz��;H�E�G�$����� B�
��^�7���������?��bк�i��ΓC+Cq�顖�pT�M�P;��S���}�Z�j����M�����E\����?�$�$��ML�p[�eS��B��y�K�<�P6�����lI</,��Ԓ��drE>{(�A��݉Ft;�S�W4�'/{g�B1��Br���Q_�����n`�s><�%����ܵxn��Z<p&L�v��>�b�G��&҂�]���	NV��fH*�aH._%9��]o��x�Q�b�4��)��!��XvT�'��?�袵��})f������C��{,���n�v����u~u�z�*yp�'�q��Q=m�P�̉:�]�ܪr*��zV1!V�YB�s![�GX��������R��ס�0�C�0�]� &��&�Ғ�ań�0١��t�kƕ&�UՀ&M�>YR9��]���i�W���X&��}����bC��5���6�}�r����0������KA]�q��T�����q���Z�kyÉF� �5��6�BTX�d���v}�p����C����d�w������r��م_4Uk���M���ҡc��MϞ:<k �f!Q�pc������
j�0`���3.�f#���¦εI����W���[k[�1�#��.n'�Y���9@�M�炐�}gQ(��$�*��͂�M�KK	�C����G���zL5�{�v|�~h�޾l����d�+�4_
=�s$'G��"?��{t�Y�H#�؊3���YG3��"�1Y����7�x�+���ry�وOX,(/懌�f�E���>��Q̷�n v����(���H�)�_'��8v�8UN��睄��h�lo3���ɽϛ)��'_b���7U��m\�����1y	B��t0�)�.����Gr��B��"@7L1ʛP�g�D�q���YF֥~	�����h<��&�����07�3�D�����`8��vm&�6���H����-�I��~�f��5el.��"��[�1������9˙��k�XcZA�?[IH�l�.���o�M�$Y�P�~1���~�0.�^D�aT��5D����� ��)����8[Vv>/�;�A1��~H_�'�e�(DQ�˺�~f�,b�[n �w�ͨW��5j>����-)�0#�E<�K�������k����HF$=����v��0�C�����<#)?w�#�f�«�U&�Dm�in!9��}���u�X����L<Y��R���۪o�.>V���w<O}����$�J��P��z�5�֟����"��\ �_�Y3��	2��'��������#���ޫ�n!���vd�~7 �Q�f�<��ϺmNB��hJ[U�\��p��!hQ���"���O5����љ���^�%VpZvW�����[e�X���o��LL������Z�'�&�$�̕$kٸ��9��~�S�6����f�2��';�ȣ�����]7�=@�/�XO�l�o�Thۣ|�p��<m�^{F�<"�5k/Woҩ`���*���������o;��=�{C7��$d����S[��j��.N�G?��!��<N�_�ޡx���ĸ0i.c�_j/h�m�9�!��S#�za<�i��'W�[����L�|2X���!]s�����d	��M�=X
 s�n�b���MW�#��K��������gg^ �/8�va���#)?_��y"�z�Y�t��J����s��*
�K5���P��;��B�� ��P�����.As�%ƒ!���XV�_W�%��N��:�p��UJ3�%N-���\ �)M����(���.f�M��,Ɂ��ip{sp��mEY\
�?��<�%�E��뉖���#��qb\��0��v�7�=:��T3/๕���}�?(7cuX\J , CM��.��v5p �ځ�H*J�|<���9�vJ�Ta�y0p���Uf;1<�h��Q� Y_LZ-#ui��4H�P��L�U+\�B�W��KJ��8�Ϗ����$�Zn��(�*5P�����˄�2��F�/=u9�N?LZ��\���|�>�oQ��M��Tݎ�_N��a�׷���ױ�G���>�Z�Bw����(�(���Pj&^Lk���Y�ȴQ���������Bp\Qq����&}�c�'�
R��;P��%�!݌%(�3�gK6I�ǌ�����E�Qe&}�2� "�
����+�DsS��@��J�Ʃ/�}#6<9������썎5K�����,����x�,��m�~��4�0ve�nk$عd�{�Ï:;5��44�nzLV�^��?�#�'����#$2��hF��"���c���a�`�^֎7� |J΄N�GBkY9lK���NU]b��s� ���eh�`�����bY�:g��-�#��k5�?(G|sM$�.q�k!j��Y��>�B�{���ǜ�����.h�p���;pF)��9�"3W
�E�6x����$��b������J7�aiP�����\.��	���7=Q�7��;��s)P�`p���A�R턇KkT�����d��y��s���j	�h�'�eʎf��IKI�����s�>�]�����BS2j�>d��=h�	N�i42��jmX{����s�qJ|�k����Tk���Q�`�w5�?a��-�&����|0���,Pp曽4e+��2S��P�-��ؤ�

��j��!aö��J�y�g{��U��Y�ƫP1G�g �W���p��AX��M�R�"a4^�W��_g�Y=f���ʩ��&.f���;Ǹ%{P�!2]����C�aT6Q��5���$�&�dW�>9b�qz0R-����R�/oF[�b�a�ō6��~���}��(��i1�t�\�<S�+0\߸�Mzj�(�?=r�4�] ��:���Y������i����p�9�r��Z��7�j�a�(+~/�T�����Yq�$n ��}��wqOy����WDc�h�#9*���K�R�sA�&"w�D
vC��0��I��H(8��i�)��S�#���b=�d���PBݲ�����$� �3%�r�WwN��S��3pk��֢�+�_k�Rՙ�hϡ(�W���c�а���RN����*��P˲�����@�˶>oJ��f�ڞE���o�DFq�HL׫���tx�֤�k�~�33T�f��o �gP�'M3���Ɖ��H��O,�������[��J@F$>I]T]ׯ�6Clc��Q�u�P�#[������VM�N Z����Ӕ����YEf�į3�W����W�n�J�\{��O��}��X���ܟ(�a=3n�ّ$�"�.i(WZ�,�[���"��1�(�>|R�B�}][�쉾�U�V�ߓ�Js�P��k�M����t���y�������.��H!����4q��iX�ь�ֆ�C��=�
;������ρ�M{�j������;�6��̇:��5�[;-� o�7��c�)6��)9{%"��1�0��ѯD o���s�7Z�W�(�tm�L�E��gd�1)���ˮ{Qŀ}���d�	�}���/L�~\�(�
�TeZ�Ao��\�v�b�~���P�HD�+�ÂpE�
=q�=�m�D�!V�Wz�h	�˭Q�����\;
��D�^HX6��{��}I3�sX{'ű(�g�]k�;����a���l��yp�6����.-���֑�cГ���j��ٺ�{ j�hy;\�����O��ׯ�0@e���%hW�k�}١��H�	�.w;��\O���JuXn�9��+��|Y��]�[*8�W�׋Vi�1\>�mik����{�-Q6=��q&A�> �?��--7�Bv��=rR��s����@YD+߈a����ˍ���l}�ZƦ�bY�n�&�oI�2ҿiK��V��L>3S������$B�����3W/��N^�H�4�Ͱ���w�RV"-���7������V�Nx �*��9;Poj��y[Xt�m�;8W��Qb��#��Rt�0Am4�&j���?߄d���k�s�dz5�C���!���bo�=4��7e�Úzڐ��pa�#�7��L"� >7�2	�qi�ʻ��>��mi	Z��8&�x[7u�v< �Q?�4_Pd��\��ZX/c=(��]jES����>���|w4VǄ�w�a0�E�et('].����ө��:�%�b�{Ai \�+�@
�9`����,F��o��;|>Pe!��*�^f5��)�r4�#�����Q�PpP.�2S���.���&��;�W�Ҫ �)���������"��-[���^V:���7��@ncl��X��4���2Կ�]L�hyU�v_I�՜��DN�᝖r�&2�n��iH����L­9�n�+��J3N>���_�N⑶·��/�JW^oC^��-Z�1�v};����^\�2�%������"�;�X���o
F2>�ozd��GD[L�koI�%��U����G��x^e��*V�d��?�1�kO�/���Z�ڷ�P���Uk���+�˩6:�0�ML0�BZ�2rI��DbYnw���sD���l�y	�pa���>`�UD�� RT6H������pCO¡��W��V{oMHA���⏗��K��?��5�9ɧ���I�0Y��s��u��M�A<x&\�WB��*��Ӯ�Ur��%�P�|^S�dN>��-���۪Yh��}Rڎ�a�|V,A���͇<Fd�ַ�E�;��O�-í�R8���r��M��L"����
�_^� �N�&`n�w�[�j�nI�K ��{;��8��F����D鰠\�X���8�O`�d��E�@{�҆�*��&6����wT@rv�)h/e>xF~ �р�Uԕ�_���%�6]�g�ɤ
95U�$d�bۣ��k�{6���F�63��)����Ir0��Y������:�ܡ�`ia*�]��[�H��<�݈�ȶ����z�5	!�[����e�*y���g�M r�?P>x�l�J�sM������y���8]�!ӥP7��^(�%����
�7����gi��oZ-�䤩��y/6�w�,�����d�g1�5���Px����Q���b� ��r��5�!� ;)��(��`�h�@<K!i��J�_e���,�����D���D��<"�7<s���2v�~��.��`��AH1,���V�0EZ[���=uJҪ/Ʊ�,������[('�s�e˝����?��ґ馭��o��PR	���t�(��n@�6�v�>�.D_;%�
Ef�� )9O�J�N�Ľ>���!o���op%����(\��rP�9�?ɟ�@��Xo��Z�|�/�|�I�x��V�C��OJ*�����!�Ċ�~�v�n$���|�պ�ǳ+_�aN,ό�8iiv�t	�y���� ف���B��T�A0�����Z�go�d	F�3�[+!x��І��Pę,�;Yӆ����8�U#-ˑ������\�}�}�ͤ�Uz�*��-�S9��	�jܴ�*#k޽T�ˠOf�p�1�H�:D�}���A����D����S6ԍ� ǒsd������}S4��S��:a
!N���į��`�]���J'iCR��NR $b�����%��|�"Q�i�V;��Xn�z��h?Uy����ADY���<�E�����L����uE���)Yk��e�X����U��W���4(����U�L+�X�~�ڗ��wc���J�Ҡ�>qbZ`�_p�)�4/#n��?	ѺՊc�2�Q���5��b���u5%���I̴ӢiC0�Ԕ���P�lN7i���~f<��.����¾.)����T��c:�VQ����,��Et�g��R��pE��Jؚ�7�7UB��PnyC!g�awp�oA��U8�k!��N�~���6�B��h�C)m��)��?�J�]j|��¦a;e�����2��B�釬��A���k�ĶC���:��D�D,2|.����7��}���[��fj	���طI�.e�s�</M���U��n�K'1Z!"����������xBl7��2���1K\���H�v��/)��^�@cgϸ53ު�j�b�nA���ɼI�Q�c>hjDN�dQ/���ٲRo�Os�m���\$���]Ȏu$^O�.i��*�J�Ⱦ��f8�&��F	�)2S8Q����mRi�Ȯ�"�F8JFy�k?hc��T'�k�lyx�ؘ5fA���*w-:c�݁*Ne��8f��M�L@<I5�k�AJ�G��7@�R�}b���"3�)���r���		b�q�0'p���A^s�t��Q"u:�!<��1;��S9��/|7摅�}�!Jx1MSIY��������]E�Ce�pF�����?!�al�iX�S�=�٨��0��ҕ�W{��=�9�ߘ�oa~��~���~ő�H��+�����s����;�����Np�COL2��i�d�BkrlC� Ѷr��cb
,>DR��3۸�y�.*��yl��$�	 �V�x����-_�*\y	�� ��L�9���>Jb�X�"�Z!a]VE׾+�mL\wL>c�ɮq����E7��P�+H��v�y=K*
����e��SY�W��3ꌎ�:��B�b2�^:TY|Z�PU~��;��$2Olg-?q�̻���L������.� �T�Y�`�iCF|�'��p��Ň��
��0B݌!��Ͷr�ҍǟ��A��x������ƻ�D��D��"��3���jD���0����q���[uz
̔�H;�1��v�0�ݰ�<I,Ќ.ޛ��,�T�2"��a ���IU5=X��n�6l^d��MǦ�غ"ltN��7�V:�^ %]k㷶=J�ǓS��E~­�20.C^�C��;M�ۧ|]Ȭ�m)7X0Bli�wţ�k.�����|�Ʌ�c���l<��1�}�vқ��f축�������<5^�S%>f?�-f�i&���PՑ(�
<�E�hu���Fe}�D)�A#����ӗ�W��3H>�i��:C��P{"N���9;%�k��B�$bs\.��r�Z�G��E�]�ܘ{�.@���g
���j=
5�-����6(D�9v�U��M��q�`�i:׽w�q�;
M'*�Ɩ�������us�d;1f�77S }��nd�x��͍���F��'CH�5�í�t�W�UG�ԉ#�7�[�]����_1��Q:�W���U7���A�3�b.��d����&�G2;Ff�1�SY��ʴt�LY�e#�e��HF` ec�1�����F-���(����H6ʽ����V������؀p5��҉zat�둪���t���^��%�-�k&CR�8�'-b��G}F+(���|�U���Ɉ6��~��U:�f�+��t[�j�TAx����PQ���-B�I�&Z�OҤiI�����,���鳡3����8>؅^m�q�y�ydz_@E/=zHk�<�S�׎�`���|3Çו��(]��?��e`�L���HgK�*n6�y��|�EE�����-ۑx�����)"���#�M�j�0�RDU� �	�V�����:�CEO�����FE�)���Z�[����۠�bj��XpmJ����\`S!��)}�����T��B[��Sk�l9�����e9zY�� d�ȩ���.�G���l��P�	�y7	׳�E+pE��"ş�ΐ:��ol�D�
���_���q�fkga�n�'q5z��o�y1�?���/�<Z�wKrx�i*��ݱ���}|���o��=��k� �.2ҰkTt/��������U.-Ùg�)�1�*�h�p�uT75�l���60�ĂI+,<g�Mթ��fu"�`��_��x�Z^̙��l:�M�%�l��d$��>�RG�����өT�N)�C�Op���(R�ۯ/I_����$��Ul��E}F{!�M�a�I��oh[�����7aP��h�m��iK%�?��/��m�J��K+�AݪW�E;�A��t�\gj1��%)�}G~�8S��bi:$].\o(+"�3�2zX�QI�Ja��x��ɷǫ�u�׮�
f��^EQ�$7a+0���Z��03S_�a�9�-�çĚ�j�͹X��]ЭSf����@�B]d�����k��]ae�3���U�p�})c�d�b=Z����3v$|�5��-PC�4�8dVp(��+�(���Y�5̑ޤ�TW�!�>��:�N�K�ՈLT�5Qm&��.���z����.Dۥ��+p+c��|��� ��g{���H]v�1��ح�|D��q�\096F���H���v_����W!�Ψ�}�q�yn�%�'�I������p��1��2��U`h����2x��U��LS@a�Ž��R1����f]i�������B�%>�ȸ���C������]wǢ�AM��1���!mZB�+�]���9���H̝S��O�5Ԛ~�h@��-�s�x��8è�Q$
�ne=D��Dy7�,WL,��^���@o-������X�� 
�a.�i��SM��w�a3a�wN������tw�<��n�,t��pňsdj}��qw��"��`^O���,�Q,(�WF�C����kO��3fތh�>T�������y���W#)r�$O,�6.θ/����S7$���d[!禤��y�7�rZ������m��Y�tVh��C� 4a����(�o��>���/�f�e@��=�6o*/��'Z;�К3|0���{�{��%$�KqŮ�����9�Hb�9�^��"2�_�@�7/q׼�������L��Z�ơp_bPO�+�2�2���S�&�� O;��^@��e���;��l�g�2>���R���J�}.#
#^��\���N�`� ,�n͖"9�l�?����Gg��=s���W��������C��C�L���M�c4hGk#y}4���\7�����f��=V�g�T��^J��ާ�O��ԗZ��2��[b#��Ϸ����Ҏ��I����˜os�Y�4b�/� ��G6��|iy��*�FK��vB�v��i��m��
yխgr^a�UV�Ƿ��߳�kɑ��+�%>h��n�#ڏ��C����Ω3�HaA�nI��6ܳ�_.:sz��ӌ��L&�<�A�M\���v�8��i*x���vYL�n(#�ã�e�z�ps�;9��=�De_��:����ǥԗ:jǶ(����5�N6��ib�f����5嶟H��6,z%+�
��4�� ,N��"��R��@����*��,�h�z ���Va^)x��c��8
�4���*�~�;�s$�������N��/�c��I��^���&�5Lg���C'\����`�6��r,�_�� i�"9��-��SԮ��+�쫣��T���2Q��?��~���%Hu@�r]�K�bp��U�s��:��u����t�����f���[{ϗO2<���\F���W}�j���d4F�7
m�!�0 ��2��C �r�M>Jxz+�S6�s�\�?�fS�Z� SҞ}���n){��#V�l�f��K�u���X�������v��]��y���f���s��`}3Y�3UH�g�1x�S���vJ��nc4ݲ�F��I��M�ʺO��	�E���b8V�����gG����]�C���r1wrU���(�|�7Ǩ�E���<ݫym:�^��4�m����z3:��Rه��p���ꎐz�1M$>J��Q<��jG-]J��� 鎅��D�6μe	������r��I޲��H��^���c�d��p�ӎ����|�z���Ϗ�䤣�����k]�[t��:�]�u�i�&�X��ڼ�&(���R�����^oX1���uE��3O���-�\XK��ua,,~VERQy���$���+1C�sz�2O_L��Ķ�K��[<�D*�l(�B����o�V{�Ѣ����E��A�z��������R�?�ՈYrWZ��ܨ���.�G��jѼ�����Ց��J�,Xɥ6?�	6����B���=_���@�t�����Ezv1�i���W�+���?�2F[Y�Y]��a�7��T�
�GYH��Iװs��F���q4�O�q"��=�Q��9�L�;�c����XF�p���sÑ�[��ϱ�r0�&컇ωN	W�`y�ĭ��Jf�;w-
qJ� ��	,1��5�ʆ��(uw���\^\%M{�{׳[ e]���'Y?�C��ɭ!���U�j�M�!A$��#l�6; �MܩO�fw#�N+$��~vd*�w�D�6z����\��i���8��v���*�������#$��t�]���r}:;�%D�9w\wcD��R�[�`$=��y�`
����Q��ض��',����3����EW�uw�·h�=0���jO��c�UpNBW�bΣ�:p\���+�)��!�m�p��:����2�t�x��"���:L!R0�!��r���=�C��g�M�C���/�ـ��SAJ��9Cx}��
��ܴ1�@Jɧ����q(���7P4Y�@f��rݚ�y��X �`[K�T�O��]~��ߜ��6+�~�^��'BΤX����w���R���	�;�e�7Lz8���Jm��.��Z)�)bpO�m��'l����[���
���<��x�'�u)��]}�vt|��'�|�iF`�=��F\�tɥ��i�7�9��?����$���2�w��7r��(	�l�G�$�+�_E�8i���kS�7������w�����'�#��H�$�� 9�?s�����]R>�(imD��R��$��lR՛pHje�Q�LT��{9Π����y�.�ɓ�5�Ǝ��2��L��6FU0SU/�3a@wF���1�r4�W���ɧ"U5�CN�P�D��%ʒ�;�j݋���3��m.��G��Io7u�>e~|� �u�=���
��G���C�yz*8=3��u1W�(�~���>�.��x��]��_�	tӄ>S��}O!Ϭ����ŭ:w�٨�/�g3���J�D����l�oE�1d9�wl���"
��A�����S<*�:�d�^�����JX)�Ƿ�;�S�1�!b��y�nn��z��[碍6�:�ؐ'�rE�Oq@6�i:�Bvu3&�+U�����x�Ӯ��Zb�~���̔"�k��Ȧ�����d��b�l>L�ɽ����!=�
��j�$ ä��+��%�&95Dy�f�49'X�m'd� ��m��Jۑ���qM�4J������Vxsf�"�0 y(�7��N�,+]�۔��ή�srC�:MX·��{NR�23\F��ȡ�MI���h�	$��7k��.]^�\�Mz��J4E�d��p�{Jh\+gY�������0�]���a�$ǀ$
i,�ˣ�I��8�j�$���4֤�9��(��e>��J�#���fP�!OӨ2���G���'H��0hN���J��c�{4x��9���V��e��0�m�C��`���û�o���GѶr@S ƿ��'���U����Z�o+�}Z��vw�/Z"U����4�!l��d)-����ސ۱��E�ǌwOy�"��V�o�W��c�.�Q,"��̸-�?����}ĢK�ۅ�^�������Eo����5�X�D!�Z?���-��N�(wa����L|-ݨ���m��f��Ң����,&݂)�-�G"��^�9.p76�A���Vc�ն�d��Y*�c�u��Y�ǭ�C?y��i�#�v6B��ų��� �5�r@(���
M�/X��]�]c�!�~�����YpE�'��T:0��	�%��{�~ηa��/�s��'�3���e����F��ҕ���ed�&·oj,Ҍ�#m�����`���m$��^���޵k��?�{Ґ���8��ɟ!������(�����8���)��=�T#�?�1�8v��rp!�G�;�8���fΝ����!Ծ��6ގ}�'�d_��c�c#|��YfH�ٯ�n�}8�R��p���-�W�e�y�)ZJ���N=��>�U�V�t �θ�`ٔ#������	�H�c� �.E��P���*�?�R�S ��]��� g�ܤ0ω'��p�u����eX�N���� �.7y�e�M��ڿb��A���e�y{8r��3V��.\� 3ޏ)6���Z�a�kT�j*���R��5/��CT���M�ϳ����7�p�R[�v��y�J�HU����a�`� ?�nS��C]\��q��֦��Жx�=5F�Ф���.Mhz6X�)T	万ד�X����E�ؽ��=5@O��c��<�à�mz���V�Gԓ廃C�^��bȔ0ιc_�u�~�������Z�cR��x�N6�8NwG�5��pP��m��ާAd0�������'"�9a(vT�ϥoR�������,ʜP(@��h��qG�L��o��J,q��p!��eYz.��)��ި0�:���g�3���)x�WZtʜ�o/���T��t�w���M��
.�U�� �J���1^s�� �ٻu��f>�b5�x_�gYΊz���HK[�?�a�C�����G#�3�v1"��;dE.��a��8�xBJ�����ކ�Ա`�^�x��u��\HoA�w�q��6�%�yq��vΆ.�Ӿ�L�+��6�=ƥO^=�
s��y�΍�g���a�9��� lr�X�{�O���@NJ/W��r�n�����6{U�;	�U�|3i��߳ا�w�K_RZ��&x����	�M��zV�'#��4-z�*\B�Γv���ji�1���5�}�# APvO��e]�֯�>��0��ܓq���RJ�3{՜��"=_��e#�]�"nDI��W��~=$d��CPfL�\���Q��X ڏ��ũV�Ʒ�l!LE��/��}y7كե���M�"\��*��\mǚ�� |�����Z"<WhMx.lz^u���Vw��>�Y$=T����X�Iʃ �8s�D�����~�npO��@: �r��N@G��}X�������<�V"�V@r�|B�h��3��*�F;�;��4l��4Lͭj��cCm>
�*��J����ԺE0\�vƀ�pݕb�J5#�|���C��iS`�y��	�O�7�a
��v�j�[�8nW+(S'�ߖ�X����E=`�4%�%��p����|��<��&TiA�tQ���e,C nU�d����Gx"饘M��
�э�3�T�2vwhȞ�ُ!s�-�S��/$F�ئ������͋m�~���w6�Tnn-f��E��޳	�� Ҽ^�ZTQ�y��1��o�RIv-�,�<�.5�.н",׋����.~`�)D���hVu�١�{<�Q$0z��Ɂ��F��Qm'}��̇�Or����N(��A[�����B�#���C�J��\e�KK`?���F��C?��e���*vz������R��5X8Cʐ{��s���H��Ӷ��$�H�՝N8@�^ܺ-k1n2"M��Su�Ȧ�H��)�uI��n�{�	����ۄFp`�(v��a��o���<�O��UZ�V�V�57v$H��c}����@+����i��92�����s�������r# �3f�zV�>.���'>'��^�y!|�h�L�h�	K='� �ul�JIp��x��F���R)�U~iA�����[F��X�2���7i�{<%��� �^YDs�1h�lS�}� �)Rm�y3�Wb��̮���d�������<Mĸ�UrւǛ� �@�=�]���HR7�4Sr��'û=��Vdެ�P4�j��jN��}��%�Y=d'�,P��Cv~��Ďm��M��3��Z��B�no*���k5'���(�ʌ�du��
��^W�+��0�D�F^��mݿ�I�dҧIr/"w�r
݆��*ܛ=�ȨXB(�h��B���iH��� &*�ϧ��PA�b7x������	Y��6 *6��$�,L�e�q�9`|a�Y�\d�4�rȍ�٧���u����Ƕ2~�IY��:�襣�˹�(���V0�_�ɕ~��]O3����V�d����.ט�/�Zk��;~���k����5U���.�a�����`�N���̵��ֆ\���F����%��~� ��Q'���k��Z��&�®p姛�RW�l�2ȖN�Jg�S��{�!v|�l�u��x�9�<���N��ãKx7*ւ��5�����t�ZDAd� O݉�)��vT1`�H-��9��B,�]��85B������@���ɣ�e}�"��s��y�E���ILC�ꈄ�y[3gB~;T�n�w�<(��X3!��;8�[iG'n1F��N��9=�;*�?��!²���� axD-��u��.Y#eY^�F��
f��,B� �_�>>������E��a�,.V>��ׂG!p��Go���,V����H�?����������(Rl4���1 6�����~t��L��s��8v4R�ۓ�k�����m���h�%o���c�Z}�M�Dgşo=E(D0�W�.=BG��L��ߙ��
!�,�D� �bm���;���k���S���t��db��wX�5`��_f���֋����U7p�@kdb����W/#u$���,#U }΋m�yJ����a=^
� ��?���D��n��%�S�����M|��I���#�x���{�)}�p�������od���;>��t�{%�c�xf��z}0���.�I����|j��n7����̂i��D����T>�?�rT�˾H"ɱ+�����\��z��;J��ꄹ�P@A�0��σ�� ��4���vx�E7���1��9�����Zl%ґ�n;�Η��$�+k<��X�e��O��N|���&�MWIĜM�vA�(�N��6�̄��iCŃe.�\�K���w�I)cj��O���1�%Y�����'���i�R��R�{��7�����Tm=���>�Fm;7=�$�\�i&�x_Ӡ�6�Ti�
`��M�&��N8]�F�-�OՈ� ��4�dO.�˲N�V�y!�l?���G�i�U�Zj��:.������N��0�/})��M�l6��#��0�S1�v����8Lr���y��H��]f��]0�s��ỉ?��/�N�,�6�B�u�}j���tK��ߛ��m��%��k�瘥�-L?���x�>���T�S��?�i�p�f ����B��>UE�{��|	�f�e��p��I�d`�F�i�!J�6���P��SH����iR��ckP�Xhd���<%��l=�2�O^�d�6�҆IZ��E�m�~���Suu�,	�}�
����++^���
��b���+E���D�Ox*ҡR�G�#mK��
��7ƒܧ��6�,]�z���v���-��vM�>�݉��7X�4�ꁌ��3�b�_����!D�R��lѪ�!��A�����p9���&g��<\�����(��������m�	��z�}R�}<��V���"(�d�4�kI*Wn�Yth7iz�2��D� ������Ƒ�ŕ�Q`S����O�[���`y���.pV'��n��+�k�L/��ͻ�b��� '��`�0w�����	F�=��X�DY��� |Ҧ`6\"���x"l7ض���8Ch��j����=����l+�T3mt2�'Le�b?��e�3�򗯨u�B��H��sq<	�Or��a��g@U���o�\~!�ogۗR�'E��/dp�(aU}H�c����G�G���x>O����)e�a/�/w�^���Y�"��N�J(n�!���<D\�# �Ǽ�?�6�	���3�	ۥ�뽇x�(6e�z3�sx�a��K�_�����g�����;��N�ߍ���K���zXnqr|�e:ȜQ�
ʠ7���m��@�e����� ��͈��H��H(���x�"w��=�	(����$S�s^�����w��ۙ���T\�A�΀C4X���Ǖ��z�l�Ѳu��+ל�Kl]=��Ou�:L� V�v*�f0��fIο��sL�J:>.2��J��_6:r�����x�`�ר����z\G��i����a�9�*�T��tR~3t��dҮ�h`U4b-
�:�=��Ug@�]�pWJ�I#,�(uW�y���Q)[ɆV��Oٳ��f�,��J{j��5�j,���������_����ʨ������aKۃ֐�v��!o�.�"�Q�%3믾j�6a�`c��a6o%�F8���� $Sr'�(�ʋ1�����mH�����F���2��s5���B�"i��-���*n�r����=�gep@�`W�'��l:�5��&<��Y�4�]�m�ޙrj� ����k��ّ�0{� F��x�SJ����p�����6&eOSV�!��+n x5{���]�슇��A�,�/�J��\��g�;CƶTG�����&�������~X0g��+���7i��3OϓO��2���x��2���ŋ��A���ُl�'"���6����<݅h;z��)r���UOպ`�rӘ�����*�6��Z� j+�o"I�tw<�ڵ���6S9�@q�=ˑ�V�y~��߰d����+�9�z����%�aN'`�,ӡ�����)?��՛X��65�=rC�Iʶ����9n5����k�A[�![k�|�s����v�����@� �U�f���y�9��P����9�0F^@Y>Ԏ����Z՜b�p1<�xel���Xj.X�q�3���e�}�ƑH� &vѵ��$��]�jG^S$_�I�>2�O���OpG\j����C'���_�9�,�q�1���A8	}�Ϳ)�����I����Tw����rA��_����\8�&�DI��
�6����h!�<U�����}�PyA�E�t���@��F���-C�g�|�`�<H�i[�v��G��?L�#S8s{g<�
9���@�c�>�jX(ǻ;��E�!�^Q'�L�<��K�_�6�c�+�g�m�U�~�9��Ϛ���Nj}:>����Uk�ib֞�9�$E)�8s!��C��9o��Ae#�c��^���%�5���Yyh��"S>MG+��;� ��iiȖL @Q�J��`	�bW�Xo-�9w��l]N9V��٫P/�K��VG���<�F0}��'�Xu_� �l���헉�r6q�J43Z��|���ʟ��J�$�� ��D��4��b#^ӳ���^�$AZ�C�-�pƢlm׽Gr�_��W��|�@h7�_�����_$U��&<�1��'��Wuz��c��5x�j�������*۱_[��/G�
��Y"��h^�a�D+�1����,�� ���sg(��Q�C5ـ~o�#j���!��U���I��X�yugA:4&���#��W!Xr������F��denE�i��]��)�˴���}?�v�b@mӨ�d�T~%�7�C¤PS8K{>��8�t���@�&�5Ji���x�K��)%���oRpT#��fh�jW^ϣ��tt�Bb*�r��O�S��(��"���8��9�D�*Q"��g-��������K�=��Fdf��iO�>�d��t,�&8��t}Āx� �vI_��(W�Z���>��E�-�x���:g�Pzcj�l�ĕ��^�ކ��4*1��e4������j^��2]�+�7/~�)�2-���^B�>d����y�zz���&3�ޅAFP!�#�26��[f��LQ"�(4����jP7������Xi�{O%��v�Je�f�����ª��q�~r�?!��
n�v�g�����T�j��X'x͆B]֗ь���q�,�.��Σ1<SC8����7��f$GJ3�[(<�c6}�	��\k_Y��'x�c��F��������_R�ۈ�b�zٶQ��^���8�!7#nwA��<ܞKBE�Z��*\���D�|�o��w�^��^%��7��hZ2������4��.VE4���W6!8�
?/�7��f<4�����q�+7F�vL�� �!(�5�����Ui����6��w����\�ɂ,` 0h�/�(MU�Ћ�CX��{xB�����s�4��e?�>����K O�8�ָ��	/��6��@�5��t���N�ˊ~�K@@�J&�d�T�^��Ǎ?�&Y�.q�;|Bx�O�C�E����uB�@nU����o�|7Ϣ{��$^W��l#mbK�n��μJt��T�;����i�F�TX/�6���
��v���ߛ�}��t���w��ɫo�ǜ�[���I<t�h�tҲ�����O����ؗ5\�� /��~����|�͙ӳ������v0�]ۘD�?�l�����"�L��_�ﺂ!��j/S�e��t5����*)<���
J��É\T��v1}���0���S�����U�q�ʱXюҩ��P�5��YK��M%)�OT�%K��o�E�݃S�ߢ�
� ��y#�JV8G�*g�N���������t�S��@���0�?����k��9��eUw��k��+r��	��B9x'S���m�Wh#�M��L��Gs9^,�I�^%�+��J�p���J��c.� ���  jI�z�1�0��z��}fP�'��R�7p�IU��_N
�/�Wh�	�'ڿ�+q��u�)���e�E5BT������r�]�q\z�$h�[�8�XP?J�giɴ�t��
r�-C,�ؘlw��?���&`,�>��<�����~��tFb��NMY�Z��̄�M�X�=��g�R6@��g�jB�TRR�U�ZM���
΢���/������X����3��=1%8+_����Vfw��g��OE�Fv��� r��0Dz���R���Z�s�[򍸁���SB�vO�˚�$Z�;�Z��Y;��K+p����RAu3��]/��{!a���(�ٔl��W.����!�!�+ʥ���=�.�l��_&�VI�#z����U��]�ǀ5%dF�M�	�{��NB�EVC�n�n�?�����]���H�, 1�^���{�l��HaUp፡�7Z����w������A(��§w�R����I��É��ZA]�{H��$��0\�T���$Ue�ai�O^0(�p�Wi�3���>o53ۙ�*�F*�5h%m�e��oZ�up�ܪ:�k�u�=:��f�����A��3<&p�a)�˺��E
�6�4٩ǫQ5�x�!9='2�yQ�l ^��)��|�~.$;�IA���-[�7���'���4���~��Q��k����M��;�g�Š&�W�F hT��4�(	w���$��-�4�!��CO���
W��͜�jZs �zV�jy�oh!��%{�"_���[��-w�YF�/.��T�q���+}�'����l�V߸���[Ue'KK�ֶ�_�ڒ^���3���uZ�\:�SY�LYߢ�b��aM�!�C�j�{d��e����H�?�)_|Z�;�{-���VW�i�������Lx�5���^ =$Q�\_�j��j�Y�����p��Ҹ��"p9!��4M'ˆ��4?���ʨ\�G�(��gtq��$�1xF��m�U��5"������M���<��A��pH��� Fa2NW�R�؛�	����")䧞�����������P�o����fI��A���M^7���_`�)�A�ݗ͔G������(d�x�e�����y���d�Q�\#%4��}�+m��3�Kf�����b�� ����?\����|�@
v.�ku�iHߟg��8s�3P��c��+R?;1?{%5�����k�#�?'��א��8�.�� P��>U�%���
Nh�*Liǀh��X&ҝm�/J�a�|�ӃY����x�[ǻR�J�.��`��p��_�R�o2<�&��|o�5%��=F��8�Vەm��ǍȻ����=,t���Rn����y�O?J�6Z.Y�:��+N��z��1:[e�l��uz�"<:���~)�j>��VƬ���)�}����k��'��E������4R�����������a2�a�	J����}�
bJ���)7`�q;�I������zV��í��D`�ڇ��d΀IH凅�:�y�<��@��UPI�F��y�nu������LԆ�
����&\�Gd��ݸ�7�%�:No��@aP6�,��D?�X�D'|�J��\���g	�4��b*�1����!:�*�:	���Fv��}ix�<���
o #鐛���P��cȟq��	�bb�Ԙl�v9D}�`CQ�Ym�h{��D��\#ܘ��^+��R��c��:�u.��a[��b���	��o�pA��;�eo�gl�(��	�#Wmp�!a�R!��騫]O«��XI�f,�"q�b�$��p;�.b�V��{��tö��ʠ�Ni��6&I>�K��M�m�a%׿�*������p������y'r�E���#wXf���B�8Ҁ��f���8��,�����4�;�p�B��:w�}�HQ��e�����R�o���E���R|ܞˢb�תA&���e7��0w.Aۗj?�x6gsXLM�~�n� l�$T�O.	g ���xJ�
��ؠ��]w~P��ۗ�����Ga��-M@�m���mK�!�44�)z��t�p`�U�wŢ����W���<�BF>��9���<����6�[R`�r=���v�������5��ͱ��U�ٔE��d�y�4�A g��D�O)COڠ�^\{ё�*�Bd��M��ަa�9p���P�E#p���c"t��\Z%��P�d����Y��:׷,�g�wR�`c�>��Je����kV�Ú�d��v&gf��F4�b`r5,E�2�����Q��#���M��X֧�3̇����
/�&���Ay�U;F�%�2���6��Y��hT��ߗ�OK�k��w�A�g0��0���	��P��@݂t�,�8��8�o���c����~+:)C�\����-���I�n!��G�{���+u�gB�ڸA��U�)�͏e����ڣ2zbҍ#��b�hY�+:��g��Ɗ@����L�%�'�U1k�4I�g�P���Z��ki�>Y��"�0���	�i��Ӟ\ݖ\���w�EZ���%�/��M��T%j�U��=���%�A�]�{ 7�F��#�2����A����*�/�h��0��B)N!4"�0��<D{å�5,-�-��%-���obꭉ
q�5�S��k2�M�%�L�~� $��W"?�:a���Y��EC��&��n7�hQO � �Q��Bl*a���G��@5q��}쨘�|4 O�1
q����16��N�F��߾���}Q�_�T�Nͻ7�8��+8FN��=i�j0ym��lޜD &��T���<~��Z��kz�a�;t�U	*� 4��dB�Np�`x+	�B��S
s�nd��Lh�{��fL��f;�)pY}.��r~�l��0_��yL� ���z���V\E�"�)5r�Ǵ�k?�+�8��'�39�>�5� �v35��70�3(
�8�nR��q���Dtx�� X!�����U���T�"b��0�X#��;�I����dډ �k��;�S�iu���\,�྆���;̛Y`ϟ(ݗbA��s[*T>�����磍�l'�$;cbx��tEOm��J���3��D�r��&C��G���m�s[̣ڎ|+_���>K��ҽl��O�?�66�w�d�[��J��ܗ˒Z]����b�qvA�^���ՑT"���7;9�����c~F2�n/0]��̷F��J}�L=��=�8��{K��ϙ	���s�O���T�z���{�;�
��+�V�O��Ndv`�4��{}�*�M��D�0��lW1��dj8���������DN�2>�*P4َ��g�H���pr�7��H�}�_��r� p{���>�[������I�3�uxv}G�ND�y�oz"5��e9`�O
w�p�@�d�:�2*��SS�Y��UWFя���c�����kGȫ�6��2��9oc��9>Q����]!����)[�&uY5�[�E����"��Si}�]W�l܈:��n�.�u+1Q |H��jN�ȯ�N�D�䫅^]kt���a��H	�B�vrr�Ã�׬��"�5��o;�~��^7S���" eH޻Q��`X����knEs�L��R��� ���B�?��l�e�1u�&6��O7�'�-����Q�+㇡s�o.���6j̩ŏ�i��]8)�VDglk�\
�n>=z�1S!����nxk�сc�Q/�X�Y1&
ݸJ�I�EWT@�����/x���-%�l��.$R��8B��ᶆ�<����vU����y�m�d�G�Biº�����{b�pL���s lO�c�^�Y��qB�ni3#T���i(���$�l�� �ǸnLh�Szhj���_�����Vn��� o/��_	5kU ��U3V�Ŧ��,T�&)n�0�mu!�V6r�/<%���S��:V'���<D?v����M&����J�Hz��KcL\#Fn��[��%"'d�i�~���kN���^����TU������@��V*�/y���+u;�����ڋ�p�ַښj�O�k7�j�z���>�p_�V���c�aG�[�Q璂� jh���p�]B��
� HW��O��)}�y�3fٖ�7��
���iX�,���fT`eso�����qag�l�c��s��(�U��#fCJ�5���(Y�X�V��*<�mw�E$��o��BG�$"j��	�k4�E_�#k ��9;F�.�����(��	��R9�����0�4�`� �|�j�[�a�2u���ʦ�� �o�$�V!`Ň#[?�<��[���)���'~�����������ܰh�O�a��l7��{�)�����~f �%�.��/��s�Vhn� ρ(̼bl����[/��Xo���$��8�΀γ�
Ŵךz2'��$�#t�1�ce���![��8��2]kT��w�'��\v����0�=�s(��̴Xy.�N� �q�X)#�������<s|�����e1�QZ�<pdL8�S7��5���b2%NFjdw��y6x�C�Y��6Ռ�m����*׽�~��F����B����=��zaH��E������xG��B��I�uˉ���k�IG$k��)*��~ B��I�&Zƛ�ڒ��&9D�����2d�]��6u�!Α��O�@(�R�$��U�2�ib���ʹ��J��{:1�,
�O4@�K�`2U���uA��H��y�(�v̧�cvv��^HL�H4��5��ȋ4K��w1%[k�K���H�k�H�F�����?~]1y��@�2[�`L�9|���=���׹Y�.�5����ā�_i3|�H���I��3[�W���ㅽg� {�@�ET�cp뗴njFR�p���;\���8��&?���$<2���v/ $�c^�CD�d����1Ɣ_��ȗj�4�="=����+������PH������\
@��Z��1)XVcW;}f��X%�\��{)ʡ�;����J�H��c[��v�W�C�'
�G��/*թ���c�#�V�N��B2^4Ǟ/�P$r��6ZR��mp?h3��ZmIJ�0X�K:��6�	��Y�L�5X-������mF����pt%�}����1B�G�����Z����S���E�:�i_b������-o@���w��!ԙ���Y����`c���{�����H#X⮳ɕfKB�* ���K�|�O��0���T�EL��VF�ԅ��ZM�;Ԥ�@���Ń�J�O\��Q�Wi��Z~�u�����V���\!N`~��v��<��@A{k����J f�j'޸���6^&��Q��/�ѻw��F��]�DoK�[7�O.>��S�Z�ݥ��Q���;:U���|��< �ನ�[I��M��	_�����۾�F�_@�$[-x��f����Y��*��y�0��E�|�N7��}2�;КF�iJ3���z(���
~p��^~0��<��w_���ځ�vʄ�̜�b���?�b�:����7M�x�CS��ڹ�r)�y^�]�"�g����a#d@�er�	�������-?����E��E7�j��(��ap�QF$������4�T��(���L�~�_�T~�����&݁6��R`.3���m#���mh�$0��5,�h�\�q���n�L%�O�}�yѲ�����n\)G��*~��0�:�ւ0"���?2�Oy:�=�La+����+C���|E��,�/y����F���:IXA��x�S���k���,@n:k�Z�%��z��4���L�݇�s>����-���!W�nqs��s;K�6l!�_�\�?7|������0�GB������TDz�j��P� �c2���Iվ�>�	��e�o�me���6������1��L^�$�����%��s5I�(Cf�T���u:�ei&p8j*/�e���`ظ�^��I*�a8C�A��������LI�+�'�Vz����KBS�P��)>��WP�CU�g,�]xg$6�0Hf����pe���-��C�̶~5!�6�v��6�F����5����y��]��5k��"S% Q���훔�$�X��&ŭ��%�ӎm]�j�[�cu�f�9[g�\�'/qI��>�eo��܄�����]�syX�r/�jT��f,%\)3�F}E.�cN�u���&(�+���M��7A����;�|d���0���"n_2�O��)ݙ��!]j\��M�Y(Oй7�B��׌)�[4��<|�6[2�	=!�aY��3G&d���$^g��-E o)$2�O��d��v;���MnLׇB��*��NK��c�8�U���Z���o�X��"J�t�Pq���NM�a6�BK�lf�Y<�N:��t׿��BO\�!�0�*i�n	҈_�Zq'IPo�����@3z��헆���G��!�P�v���	e�F��R$�j}�� �BM8��{���h�F�-T���h�C�nm�|U	zQ!`���|w�2�Cm��	O�Z���81��ڷ��u�.��(	�F�U'�Pυ�F���������'��ƐH�J<�S>����kok>�9u�W Qx��CMZ����)o������`$%	�ea��-|��g�^�U:���e9�,w��Q���PΏ�<�Idݪ�:�y7+�+t��)�J��F⃟�s��K{�p���#r�,SU��9 �}��1��ש��8�1�,�6��˛�~G��oq6eDx�7Vb���EEq)šF�}K�[+� N�	�f���1���d	`Z��-#=��K|!Ȥ��d�_B[f�Oi4=�z̪��Q+>ܧ3a6�~E�7�%��j;��-�����ҹ��6�����
���.nO�u���Â<8�<�����Fd�V��NI�v����;ru
�`+[����oćledbE����g/���b�ŷ�\�7��4�͠�wb���u~ֲ�����Ο:�Q~���TZ"(G�.lN�W�����P��h��*����������3T�tB"�7G^c_�L�>z����\t�� �OGM'�9�)H�\�A��`	:ms�~��:�卨 p���8�r]'0�s��a�"Cw	��>g��aet�t��})E�:gSs(�#�~�μ
WV�O:c����HА�o�S�yk��D�n��7XOK�ŧ���dP�bk��A�A�f�	-���(���?�U8���+�Ku���j	J�i`I@�L1� aJ���3��!�����F��m)hm��L����,7��Y�!��6��M�t4�c�^��(�G�܌	��n�1��Z�1~S�,
)�g�o�Ѯ��Mx�F�߇Ҽ��T�q�e�:uu�o�&	�.���6_��5�*���}��u�3���U���/�o!�0c�Ϋ�Tʶ�b��oL���L�(_�s�/��m߄���8�P� `E����zDȝ&���@���l:�k�>��[��z,���������G�t'n�?��Ն�U颌���/��͇u̰��B2)M�9̫{ S<&Y��|�Ky��G�<�0��M�TPύ�L�oV���u
��k4�b,�5u���4���a ��ͩ�b�h�Fje��e+�{�S�ˑb(%Ce�v��P�-E�L�M+���H>Ӷ"r���[d�^���/ �k~M�;���H-Tc?��hl��#B�z!��ʇ�[���L����M刘I���P�U��M<]�@z��dd�,��"P�F7�۳TF)���:�3Z���yޏ���HQ��뛲�oS������O�e'��u�h��!�g~E��G �AI�3���>a��-���N��y���!���@��0���^)J��:8R�D$9ϙ����nC_����,ѹ�g�f�#!Vp��4�h��=�j�?�I�;.��}�*�QtN��p�V�Ԍ��I`��ހ��s/��x�����HS�>*´�O��4�`J�_C��b��[��Ϫ.3n��`1.qG7!�穣����Ӑ��qԁ�����L<�p�'S<=�n?ݚQn�r�$h@��M�Y�ϯc�xO���,08b�� .�o�Oh���:g�v��җ��o1}*�Ϊ���.��[�>���`�i~h���ŽX����(I�
�(C�Hd{q���"��*�Z���w2މ9%�h?��G1Z�C4$m-��#�A|x̚j��#7�9�.�r����օ��'�t��R;�v���K��D��G@;�dZ�n/�|��ū���ǽ	��:N�����ݣ�t=�����TR�/$��O��X˕�1Y�P3�b�d�y���bi����9�Q�$�7���#u� ���Bf-���wF�˴/�p�Sx��[JH[���?��ja����p�w��.�/��� ����ޙ"zd�Ұ< ��}vk��.&���+���<n/��\�İ�$�+��~./�5�Yk��9� ��O���l�~WN�����O�UC�B�*c��җc�Tm������$��@z{���}�
ˆ��}A�&���!�{ıj8�58ts��`�����?_ۘ����(���T���;�D��=��g��SP�M� ����m�3�c�K�t�.
�q��/~=��t7U�PH���Pл�s�Y��#�Z8K���I=V�S��%��'�X3}Cj�֛D!9g�194�ܵ�A��7~�"3k���(8��B��I�D��?T���RWR�h�V�o6�Eq�8ޫ��C8\�A�lC{VH�^�D�B���ʿsp�w��@a��:s�`�����#�5i.��n�rǲw������䯿C��%ew�=����"Z(j��c�{u�)?���,����.�NV���"r�}��I�0n.�yW�M0?��� M �q�k�LBFYjü���)����� ��X��EOش��2��!�^�Q̣��m�X�D�L'"㍯�5��)�����ێ_��w�������� \����-qy��#����H`Qº� �	��~RO���H�K�����z9?4��3|�� {��G�J����e����o���f^BBI$�kU,��0mU<:.1:V�j�k�<A)���i=%?t�Jh�q]�v�u��״����Y�DZ<�{�I����n]ŝb�iZ �f��$�㲣��J�(������n�o�0�R)K+��/|^z�Aɖ�{i��� �u�����2�з�g�P���#醧M�0l)9^:EN&hXI=�c5Ɋ���6]�ќm�������̸z�Ϙ�W4#ض��C���6vج?F����y�<Ђ�Da^��52�eC���U�bހ�%&G���W��{���Iq��U�s1nv˽,����E�����s�{ RcE��V�ߌ����-�,�&�;aY�<؎y	f�7���W�}c���5�%����5�� �3e��x��gp��|��LŨ�j���6�}��xB�K��߬��.K20�>����u�S���I��p
���-+dZ�қ;��R�?���
�s`r<Ʈ��n)���پ�������S�*��s��뙉�I�Ge��a��"˸�)����3��%�Y��l�0o�wml����ЦM�hYG�,�\�,Zh���v��8H��Y�g@�Gώ&�)t:�>���V�6,�C4�e�N���W:1�q)*iB��x���Q��Dh6o�?C�c��_��Sw^�� ���/�#p�n�����#��(q2m���(!��EGx����Y�K�^��H������S�p�Hd"_\=����S�XԘy�m�S���2�.�����g6���$��2%쟿6}O�X��PY��[J�4}�$\D$�������.t�c�Bm�s}�_����=лm$x?�}�C1s�^�9R
�m㽞�B�v<��Q��!����ѕ��.Kr�i|-ݭP
��F~{MB@�ץ5}�����4�jNi�"|j#��W q�1�̲m1gs>mA��S���o�Q�}����K�t�M?�܈#��J!0����*�Ak픈Q�mR�`+����۩����s=����-T��_�Fw��l�=Z`}~�wV�f'�62���M�[��m4��S��<���p�=Uw�I�|7�ѵ���Tx}��Ľv�z|x�J��VjD�4�t�0�N��
���se��҆e&��Ax�"��	�j0L)�6�I!F8�tc2��﮺REFg��|��p�!а�:�ȝfUQ(�o�K��=V��Bc�~t�m@f�'a!�Ó��_E\ ;��}$.h`�;��_�+�̔�/IMm'R�W�	7Y3����M�;�����)yF1���΍�0$���C�:�qr��2?��H�I��ԑ�co
�u���0Q�A,��ж���Y�lݖhI�#��=��?Z��k"���R��F�*'v�ot��u��ض�{Xt/��c�e�P��:�z�"B*nkV]}���{F�<�v����#A&!�N)L�P���d�U���p,�"�n7�)�7ó]��u*��A�w�o[g�����݁5�WD��=��o咑~���񞲋�X봉�ߧ��7�t���	����
����K�9�!�3a�x^�u$�f�\9T.'XXs�h�{X?HX=w:�W���_D4�!1K�@3M^0G����瓮�<.f�#z��I��'����Z��b�C	����mޘ}�CE��J�A
§P����n��/cW+����b���I��N�ύ�32��=HJ@��m����xN���oh�!�6'�+�>��>v���[U��6aF���	9�<�3�G�^�Cl-�ۤ���v��R �r���F�Vb@X�򕑎��jd6�~١V��&s��@��Bb;hm�E���M�_��)"��Iw~�ԕ�Z��ag��V�XB�3?i��ɜH���4ׇ6Cq�� ]6�._�uI`��G"��d��?,�읝r���)��;��	8��}`f���Q���md.A"�A+Ƕ�{�qv(te��&�7ӳ��� ��[3��U��Ҳ�X��x�?YUw�+7�*����U�+�(��B:uǏ���S��lHw��O#n	4,��.% pӑ��	�f��"�Dv�|8�p�f�(��i{�_���	�{����\5P�s�m��H6'z#Tlo�$\.׸�t��ɷ�ٻ���YC��x��wa��X�%�	c�Pn��O+��N̜��!�l��Y2%�c�M�~a���D�m']WRm����o�J����M�6%W���dO ��v� TQ� DI��{A4��ᝡ�P�2˼��[;De�3��*�h@��:,�@ޙ��
'�^�w5���&��B�c�y��Dh�-Q�l��Ra#6��Low�,⁏l΃���7Q ے"v%���L�.�*ݏ?�s�VᙾqS� 
�-)L�P�U�l,�wRN?��/�_�:�]#��(��c犘)�ݵU�S�{o`;��I~!���A���O���f���3eĝ���lϼ4J�/mڼm�#,��!T\ܣ0̹��-���\s;o"�X���<����v��`3ۍ�����>����y�HC�F��ObF$��3�2�Gλ9*fHq�h�٨d��q����b������z��B�Vj~ ���_/6�ܝSu���(Ӊ��[���OI�7e5��&&>03AI�x�^�����o�*���m�2P��q���r�48���5�y�=��_���%*���8l����' UL@NE�`{�A0X �8�������fjwV�&l�G̨���J�oeO��4[����Υ��fK���]��k��}�!�L�V�[�_,���׫PL��Г\ �1�5���yc/�oi���4Fg�u��Y��)w$� ��K�7�D��5I�{Z0?���Bne�Ո��F�+Ac��Zp,�sw�
�]��zC�v����+>�} �> UC\d��?U?=���P�~��k聆n|�����)�K�J':P�����{Ʃ�<�ږ,�/T�
���e�9�[E�K�5���P��T|�
�,��C0d����G��(�ޜ��k(y�8wˎpד~�U��J�'T�<=@�"��IR G�������a�U�Cc1N��7L���I�Ɗ�[�%gF^H��و�,z��	u@Eǥ�oWf]9�On�|X��]��e�b�����ןh9���ni��-�W����Q=��f�FGۃ����[��?��x������4��(�
�s��,�� JR�Y����@C���].n�[p�0���[��w��'ov��Ivҫ��42��Z8��#kW�hȭ/��,�g�L�!}<q'aC�6�l�<<ǰ����̵���w\`��TJ�j*-��7� ��9U�:9x��t��F�
�[��N�0]�Gm��� ���;B�dw�З��)3g�L����i�xTl� �������	�6��c�j%�
~zE‚[[��4�6����W��R��F��'�l�%��4���י�θk��SO�D=�N��8���_�];�������L�� o�C=����%&�]����$p�s@3��h��q�|�r��A��֬.��6�S|�Ei��A~����Vm�I�Pc��H�4	E�Pu:Pjd���u|�`{s�<V�I��jv�~����/�x�V3Z�
b�J�� �e۽��iIm|���ԛc��ֳ��aLwn�7������hY�%s@���c-jӥ*�|ks�X��>^ya�վ�m]y�JVE^~�l��|����x�r�,������0�#�����/J���j��^��e�a���f'��s4ޫ��2z��Sɓ�Fp;=y����|94&cV&��_{��]>�,WĜN�yκ�h�d�u)���@�U~�ܸ8EN��!c�&~���=�� {�u����h&���g�y�!���Z��!
��:NP�c�� xh���$8�Fa��יgC��!�k;�(?b[��$��hKVɴ�6�vס��6��[%Ɍŝ�$J4�X�~��&�2��6�Gm���N2��"�c���?fZ��7�
��W�����m����og f+���CH �owG�zq��~���l�}�oG(b��r��>UE��~�����^c����?d��d3��˰���ˡ1�7�Q��8 4/��*����D��&n��!��tD����6T��c��1�5�S����j%c�z������0,���҆�-�z�vHR�چs�C9�IsRy	��IT���+?SL/x��x�	-�����&x�[c{���&q�Q�廩
j<�ٮ'xC�n� J��?��uRf<01a�p+�9�i�����$֬��Mɹ��WB{";���Rb�t�E�"�e�~6*K��z>�yi��φ�&s��l���Z+��d!��v�m��6_�x~Cc*ަV��R�e�=~u����P[�����\W?��Ы����=��,5��P[��E�CM�i�r�f�+���V��sn}f�j���Y������-���2jי�B���M�K�\䇿�Y�a�T ;�����="��|K%�g����Zp������Ym?��wvWU@E�� 1�|�$v�Á�HKưDYI�:W�g-�ף���]������xX�P$�s�зX@NdP��۬O�k��6��4��D'�O��W��@������f�&cR:05y��Rr�3>������^ĝ�"=����ko����1P�2�[���2W*~W�[��*�5���v��>=�n]7��B&~���1�İ�&W���/�}G���2l�B�#�7�?��0���_�Kژ�e�-��/�D�
a���I=|L����UB�߳\�V����q6�f���A�;�X���������F� S[+�� ��"b��&�t��\,u�#'p��`"�6�i.�#f.�
�Bj`�q7��"�����	t(%M�`��^��埕b��>��?��������U����L\Z��z a;H2�w�$������A�����c0��j
�%:s��@e&�d���ͣU:�͗��y���X���աr4�n+�3t�����.q��G!x�w<<9���b�3m
�P�`�����-k�X��x3�M'��"S�E5�o����s�c^e?J���T��� yX(8<�`��?�~��R�����?=�h�P������E�`
eg�d���l��-���mM�FGK\>��"�պ9��y5[� �de�����>�3 Y�w-P	�e�U`��j�˔����bqx9����/��5�Q_���GT�0�(N�E5����(U���n��]�E,?A������
	��5�Ha��=ף�
�ς��e4���.U�,�tg<Jn^D�SL?�� ��̞)�9���ks_'z�Y����D���0�����b]}��p�4h�g�x��ʦ�u�07��o�G(+�*�/�Nw�5�UM�!�㺧���lK�;-�^�m������I�J���խ�b����}�cta���Ra����G^',�Ak���磧����MATLp��[,��1醋a6Uu���tq�n'��tc��sn�4��$�(
|�[�=����]���s$��0�(�#Ȣ� #��\��KIb��2�������l{��#l�f���k� ��L��ؕ��0F�#sv
i1pCW����rw�v�A?<�\*Rk-]�Nd9S��Mѽ������x��'�`d�t���VW��	�^K�&�j|�����)J�3���u~�⓻��5��=�*v�����%�xY����Y7�T���I�8t�?��U4,@���<�*�� ��M&�M�J�6�l�9pÎ���sTϷ��|�9����4c����y�B?����.z9�6���k�����9ڣͬ\@�М�Ė{���p��a�Ӎ��}�Š�2��,�����Ǘ��.�K{S��a�&*\Ĭ.�Z�(r4��v���W�%5ѧ(�����Z�- ��0(���&�۹UW���͓ta)���C�0�*�����K��eYb���Uьn#x��95/ �ix[��H�^�oI���zi 艓�X�@%u
{�њ�1}�)`���PB�B�n�%`Q^��AA�R� ��G�q2��4���1������Fh˫^����]���?�������I��9f%l[<�?$���ṝ����'>�S0�Worf�1��0k�Ռ���� ��p8J�+.k� šxB�:��MM�����0ލ\4H�7{\�1��|�H#�뒝':�'9G�㑺�B��h#7l�b<�I����"M�z�B�Kh�G����jZg%!��>�[FL6���-�1�O��YGg[ْ��+�lG�n���&�G�7C8��]�����?����y/��3[�'["�X$}*x�g�u�]n4<�Rs�'��!��]2qs���3�G��|��.�/���Wo]������)U��`Rj}���X�k�D�@��,�ѝbC�o q�hX�e*M�6C�T�����x<���{��#=���F���2/{)�.��7_�5�dȁ�2@
B��I�g'A��9c�>���w��(���P���vEs,►�� �Wɦ)ǝXg��fU���q��fË����|,_{Pvx�(�_��HH\+8][��>���*��	Vھ���|.Mk�I�$g���#@����sy��eI.�Գ�ݜЩt�(�)"��j�MjO1�%�7��\8��܅�a�Q~o�%�։_��_.>�/��0�-���B �����F!u����I�WZ_��)[�Ѳ2Y�|�4P���?���&{�����T"���hh�7`)~��?�dK��ʈdʳ���Hk|�yR<��Pq:��� 3�v����L��SM�[0�Un����;e�`FF9(�S��]�&�֠%����0gC��4�ι�Ӑ��9r��̇f�H��x����HT5i5�)q�m%��ڨ��7�/�I�ֶXD�;�^gYA��f�H��}JncZ1)G~��j�,�&B�����'Č)�%����'�P�e��|��:U��i�.>����.C��]=Ǡ'EO�O �i�|H�d�Y�|�(}�&C�y������ ��G��nN�"��d���,�͟,oK�мE�i��Ӽ3�B�N�Ɵ�IR����9�.���T��o�&���R�sdZǇ��2�~s��/��+���\���Ӷb��� ���9ӣwÐ���~Jӄ���h\�m����(��-����V�L���\0����d{Q�<e�0A�K���3j�|��t�@Q.� �����ҥ~��W�v��D
��5��$����]X��z�ן�u��R�7%��J��k`��� j0٦�R�Y�"L�Ӵũ�
V�!�!��q	$I�پquIA�m��l�p��9�Tf@뭩xHL9 ��{r�5����L�7n��ry7���E���S�&�u9���+���[)ģk�-
�,ب�G#�����YÄ�3vw���{܌eL���T�J�[$�����^��&�Cd$E�蝭 �C!@�����ҭ�ȥ�Ķ�"��u��2��ch:Y�9n[��-[p��W�^�ӣ�����Փ}X�s����z�o���0���2k�>� �`�f@�;����������%H;����[U�v'Z�)�;tDH�A���>����t�^?�;Ϡ�Z9Z��&]q�N(�+�2�g:�¸7�+�w�-�r��nn��h�2F�Zj�XI��b�:-���u�T���J�҈�����0<f�iQ��%"l��{��]N#�L4Na��\4)53�W���oq�WL��)�B��r�#�W����G�<��+)ZO�(t'�-��L�����}])��r�WD�YӶ�:%���s�8t�Q�ا��kx>��&y�����EOP��`���Fxr�lfD���ea�d =�:q�!::E��e���^���굊�"#����͟�
�_ΟA��0��taz�q[���N��������n�#\UW�F�8#��	��\��y)Ｄ]�'�m=��壨�ۃ����d���Ҥ#�RT��x&W����Nf��6cw�zukj
$�����7o�WK�'ư(��Zb��f&fӏEV�#�.�{!��{쪃�/녃�۝S:�6����6#~��s*���l5bbt!3�Ҥ�\@�b��$L�j,Z)���C�o0�}<9I��; �$��}��r�ٱWI'�u
��]m	�#�D�%�7�%۠9#�
o�u�q4
��vw$v�N{Wn]ۉ6�3���c}8���i��欫B@~$���Y��3�u&�e�`����x��Q�$JnE��6_y	������b~��>���1�{5=@��l(�q�=����j���4o�H�e�>�5�9��V��Y�eOYIZ)mU�<w��b���Xw{@�С�Ԋ_��-:����z =uD,d�Q�	�%ѥ�%/�F��h�N��(%*��0jC��q4הX�q�ٷ����V��3-��o�^��y�K�3n��j�Ź��� �i��Z�3s��#c�D�+�+KN�x��Q�#��;�XY5��M\S��"�S���u�n2[�n��X��7�����9�6��G���I�&h���eU[�g1�U~�sC��탰��>� �S5p���G�pK��X��QC���[������|Q�& 'Ǚ�կ('��&��N��	��%�Ae����d0rڴ^c�-�D�ڒ�i����P�9Oƈ���lux���~��Q���ԊiS[����� �lZ�����n��
�b�Z�'�ٸc/J)�+�i�1���%�#��P��:'`u��wTa�#���l����-�`��k*�PN�}h����~Ww.`FAbծ��ﯝ'�{t�1;uq�̕$w��RI��r�m#�,�H%G���ɘ@ct��t�;�ΰy�'�u�!������߅�K��m���u���EA��H�s ;�J|X�H@JZ]�DH�&���R����%I��ij��n��A� @C�ZI��ȿ/j�*�F���Ex,���DS�]Kr��l���h JP�2Be�M���My��oRǌz� �*b�<s|^Q^����Y��.8k�4��)$B��=��淫Z��c̤�S�R�r���1&L(Q'��6���#�K�W�=�	F�EQ$2�%p�����]�slI����foÕ(�`',�/`�иw<w���!{7�ߛS����I�YV�%���9n��m��C��e/y_���e�>�&<Rk�5Y���KW�MV�<�~��\�ښ���׹W�7jF����̒���B�9�v�ZsY�TE��W��z�9ޓĖw�QJ�&�1x�JYId;=�ƿ���8�)�}Ҧ�q7�<�c0�(���U�hA��4�s�V9��R��ex~��x��XqKd�Tk[��s�/ ؜�o��:�c��(��/-%��b?�+��&���H��WY,�=����.�,:Ƚ�>�@����Dn4j
���H>�%�����=����>�le4t��J�v���V���5[����ȣIr���h���a�Ύ����ؽCeH��5���ђU�x�>�0mi�R�7Ќ���#"m�ߊ�+���Rt�����@fm?���!���/U��9��1)��{4~}z�Fh��"�yf������Nݒ���B�'��:�z���ߖH�!��1R>Z%�$�~�D�v�U��Ti��U�@i1��a�K�"l�C�W��������k�n�@$�d;��D�N��G��m�?M�з|�ҷ�ܖ����@Y*t������I���35�]�Ȫ�!�A�Vr,	���]�ї罅ĪP}|i��W��k�w�KǾ�t�m�G
Dc1�S3����'��υ �d�8�!�Y��<|��/!!�W�В��d��C����`&"������ =E�x9o?�4_`�����=�ML�<��J�>wmnu�!X\ �����!�U!<�h#/�1T�7�p��Ĵ��:���Ǜ����)uM�*ab���h��7���R�e�����#�H�h�����鳪J+-˸�ew����_d
$��#�v�E����`vH3����z��Yk�>������j�D|Էp����F��R"f	z�`�=;�F�h�F��nq0�?��4j	^6@���p�>	m^��#��oN�u0�E@� ��A��n�=6��a:$Ў �K�qy&|ߥ��������r�ؖ*���?og;DcN�'GԂ]=Q0ߴ`�+_׈1Y��D��%���Á�({b�����|�����=0<���~��C:��E�d���CَV�U�$�x�?|Z���rkWnf��g�niY싋�e���{`�F��k�G�I�)1�k	�,jh ��e8��>�Ș���[����ɄZ�V�ʺK��Gt�5��[����ӻ1`Q"���I{���_���'��ӵP ڋ5��'T�'���@c5�)�d�)��q�W�4$�_>ǳ���oL
�ӱY�tUWT$+53�������0.n�=TyQ_�B��T\��Y�7�}lt7H���������/���{��N��?���Y_I]N�!�Q����V~-�s;\Kg���4��eRf�C�`G9Ww}�
|�Y��1��l���DsK���J��Ǭ��v��l�Dq<?5�c�MJT�j�+y�$ɧ�j��P� �)�W|r� ��0r���Qݪ�T`al�
���
�G��&\�Z�\T��&�g�ܭ3硅k��	8SI|��
�Kh��y�� fl����2�G�'������*�	�aN�cW��|v*�t0[E�E�>p�?)�ll,�[[�d4��E���A\��zm/4&�� h3B+��?ۮo��1ϭ5zS$|t%u>a"㈞�Ċ�U�?�xj����e����vŵ�ˢi����2�7o��n�l};K�S��eѝ�׽eG�Zn���~���R�k���/4�sn�7��QT�I�3x�x�x���(`w9QRz�`@�M��<���[	T��t�@"7�
�$��2^z3�ũO��Hn�_D16Jve���|��X��VlYuI�#�����(D�+[�*P3f`���޷\0�N_Bw,l� �F/�ȖVv3�+*(�"���v�=�.�,.;(0Bw��+�u�븶u�1�?)P0~�!������t���6h�w3^���V���"�ǭ��bmPD�<q�]N˲.���έ"L�y�QU�3���\yl���X�c ����f½j�:��&	<h��3F��T��T��T]ޝ�z$�t+ĎV �_��n4�!D�D儴f܎�Ul�=ԍ��j
8P��Sy�l���~�=�}�cFŨZ�<�>6�-��l�����&����%�u2�{j���䅷�N����{��θ�c
S\/~�^HN)Q�^�?OC`}W˧|#�� #r�LuL�W)��8�^l�����*�B|�Sk��>rp��a�xj����j�}�t�!�����ًZ����j#{CU
�d���)$����ULL���IFe�}�^�3][lF��&y7�4j��O%�&6`F�����"A���,(���� %��*|c�O=hY��'7���3������@�;K�J���v,Y�4���ZX&m����1�4�@r)��{�K��,؇Ԗ��� q��7��d�r�m��Mݲ5�<�
���P��|�Ύ�eW.io��M�J��#y�lK��m����}�2�gɏ�w7��;��y���$�q�g�e T�y�2�� N���%����E\R��Qǻn��6�|�3�#���e����J7�kTJЍR��t,��<	�$�>�rO�6��e�Y�t�����Yr�c�LAJ����&�c�U��@%�ڷ�H~�@{O�̏ǻ�������ZDVz@Ϋ��s���L� հ��2��[R��\��޹�6�BY��v$#��U!���U��n�<��$Oj�T;�N�re� x.�}�b��G�`�܎��.�v֧�A��?AN��b�<�z���˲��W�BPZ��*x�X�ф���i����1�I��K�,M�x�$���
��Kp�W/�Z���Z��'�Y��?��
���|��Y�rʯ:�$��_�4��q�5{h��>6��)J�`Sy�`AX��~+`��>=��l>�$�+jX�(���%�ׯ�������0T+��/z�'������_�'�E����HIu;��E��m}�s�*����Ap��U~�fv��#�3�z���A s�׊��՚݄u���&zP�Ո�M�9�Ra~�L�:L�H� ���Eb�?A�?[Ú���k��`��SY-N���_�?���)P>�܃�����n\�s��6�ވ/.�;@y/v��ݵ&0ls�v�/M+y%��)��h�8]�pnĄ	�ɋ6M	ϼ��,?>p�F�tk�E =��FP�V���?|�-T�618<T]�8*� �c�[��w�&���g�8�l@�t/p0�*#uՌ�&E��"�!7�E�|��,j�p��˞�K�גr��3CmVt��~����X�L=��`l˒�q�6�$m��IF�Ps�j]"�=ۢ~��&]����������#D�ϰ�qwc�]�s�9��f��R��������&�@ko�Us.O��:����_.ϭ��&Tl�/ϔ�`�nى�.�s�.}E�'T9�!�F��)�p~p������>f�%���5T�4�~*���H�fq�߮?�2��3L	�v�_���6���1��;��C~G��c�W!�#ƨ����@�_�n+�^��A��Dr�a<O5}l< ���#V�����0ս?��W�����/��?��m,ϋ�L����cp�s��Xb��p�����{Ah��r/����3�}����Qv$i"n��W��k�xv�b�%�2Z�%{�X~�o�Zu��r�"���w�n�a d�}���0,��^ܬ��<#RЖ@ٷ��ZH˭�?�����?���B�0���$U���p�˅5�1/)��:�f^�lO���)N�����[q�K�N�Nu��p�#��%� �8�M9"/ ����^�R�F�a$&Y�Z�l�s��B=i��A�3@��-EM�����rl���F�h�n�JY`!�;���IwS��j�l!T$�����2P#�N3?}e���Q+���(o������Qy'O�|�Hy���%4��H������Na�՘�6N1U_@=*o�]�Wv8�S���_�S�ad���vX}c���[[�����H ����D�7f�?k�;�-�z��>B��}*kI���0�vj�V����S�vF<��q7���M���B��Z��$�f*�ʚ�h����Z+�4<�^���
e��qONbY���~��Ƙ������GQQ��wW������>����Sd��L�]��Q(8Xg�;���<6�Pd� A��s
!~yK/2��T΋ODK����X�g���c��W��XDg��g^��Of���,����
e���E�-9��m�z�a�%��L.S�{���1:�q���,c�n�%J�M������|�l�q��
*�����zT&Vp�f�	�J�Ӂ��W6]ƭ��<����ƏF>�%��^P5Xa&�㺚��Q�g\(�L��_�4���0�'P^%�Q5�f�k0u�����nln���������I�=�����y���7!����N�:��#"�풺���׎�s·��&��*C1�f���=9灙`�$/,������e`*��]������Gu]7�4Up�-�o�v�X�x� �Xq-�|���e{����$K���I��@�ڊ� Q3���j�C�g>$��#o{r�d/�n��E�Y����	����)��䂟�䮐�6�%@���{������}�;�Y�S���2�\��k���s��5a�� j#��ݣ��8E��3m|���ݴ�\%_}+��d��n�,�Q��v��9r�c�]y)7�8�(�b0�� 7n�/#%����q�j�� ޽T�揔zi���(��|e�N�Z$�h9�G�,�1 �8S���/��%���U�)^�״�LMˀ��B���=���D�e��y����a��x�&a0z_��a���z�ao@�	�՚�䳺S�O���ek"/��M�2�z��N���G*dQ2S�>�zr����Ԟ�9Q��ڔ�+n[��#����ibܴc�1��[#������_956�%S��Y�mQOL����}�&c.�'if����̛흟<��6#@�`)�i���j�@�0O9�e&�9��(s���;$3k��c�w���{����m�3� ��D8�1���:��x���_���N>��bwi?�r6���X\ͺ�Y~4����C
�gŕC�c�q�l|�HwXxa�9C#�a�a�3S��fǜ1��liyv����m���U��5x=�:��E�]��}����l��Q��5hAY�1�=<vu`��|H�	���v�P�.��0H�x�n<pk[#�׷a��B��mzT-��y�$&�yx��\���R�&ª�+８�������- �?�3.�>?Ɉ U�g�����B������V���� 4έOĩq��4��G>�*$��Ci�a�V�X-o ��m{!��h�N�a�T���t}�Tgsqe3�կ$塨) I:�U����_����#��=�y�m]�/Y�2=<�<�yjl�`%\��"���J[�Pr+�w�PK�h�P���Щ2�z�
�\%=�Y=S�T��C<	b�����:"�ɃTf�r�`c=zQ��!�U+�6{%g�����i�"��T��^������Qb����,���Ӯ;V������'���l��T<�Ϊ"�ZyO�v0��|�QZ�	����&��rt��]T��<��0cY��$%��X�����q��۝�H���![eS��'Ŗ:̻+����#~����Z��pT�/�L�b֭��
_�3���zZ�#&���'��~UyX5.d�����=}dA�1֩~:wT'��/�ti�ڱ����0���|G	��^����!�a&�b�!I#��(U�Uw���O��nJ_����o�&��A���-QE%�o��:��Z�}SjI�Ҭ���-��#}��f��}� `��m�[��y�ĺf�,���G�,
��9U �m#MX;������Ӥ(밟��w�E����b��_Ya�1cmN<Ǧ�ΰ�F(k������CW��S��;6���h�ƞ�,�?<���FQ��ZH���ڮ����M�_%^�	��byC�l*N�N?���v{�m]��5�e������U/Y`��\���P�%q�{ <KtG}���nW��m�(��C ���9��*�M��8���ͫW��6 5@\*0U����A"�;nQҚ�����E��ҍ�����|=��wlʱ��J�P�CC+Ş���P%����d���� uT��!#}U%`������E �"�0LJ_,��Y�0�EuY^�g���t�S�;��|m�)�P�d��h���][~Ίw������_'D[��k����0����%���m	��f>�m��w/��N�n5{�����R��"���u�����X�'�����&?�aM���;w��c��!9"�4D�RfG\���Yx
��kX@��9^
�+�'����
3�$�AbI1
p4GI��w�SeKa�(X���Dc4����"^YH'���q�qn������gV�����4S�P���F�(�]"6�$hk�S����S�Tb���ڣ���Z�ͱ�7���	���D[�M���8����05Ѥ�%v'P4�.Wz���x#��r{�Ȫ5=�����V�Ve�׺�"�b�CI\ ���{��w�r7:�r�FE�*q�m����KVnin�{)@��+��,��̒��}:R���<R_�m �4�����L@*���Ww@��'����l�i�ձ��B��"B�@������%ߑ�-�2�:���=%��wB�> ?����e�d6�3����V}��[�[�p6��SD��o����q�DIt���ɕɭl�s:��(��:��Q!�mZ��-cx4QU�FHf�����ORx|�`��C�������?�K6�Z;�`x��Rs0��)���o��3�#3Ӹ���%F���BrN|��',�@�ȓ�L�@��Ū��E3�(�P�by�oM7�p���!�Z_`����	m���$�N4�\����̳�7N�rq�~5���U;�f�hvC�:��!b�}a� ث��uf���z���+�Y8�^ZF�om_�~��C��=����p&Uz�@M�fc�]�;��9F�Q�����5.���(5��"�5����U���^3��P̞ٙv݉��D���&�I�9�
X1�::Qs!t(I�����y�P�o��7�)	�AqU���+��h�._�'�Q�N*�?E[�7Sm�Sa�坰�-�9�w��O����AZN�>k$c�b�*�R��a��S�VW�}�f�!2/���Aaԛ�`�$��e������=)�1�����Oh�>̿R0��Es�Ee����,o�����7�qZ��S���3&1X92���B�8�^���h�aju[�i�2�_�У��n�s��8𝩌��FȵV��z�9������s]�G��|�9̀~�iRCa�N��]������θ
�v9��K���u���%g�����.Wl9���wlc��r���e!5|�"i�=Uy��T�����"Uo��s6 ��2�r�S�&Rnжm1�o�LrJ+%�Yr����/f"�2x�Æg0��Q�gd�<�O����I��;֟���;�5�)f�j,�U�AX�[k8\:�4n�u�Z7�4�	'Kt�d���m@tla1��3s�}����dC�9�Ӣ/���`��$�6Yxu��o��d�ן�6K�&��V����dO�5�ݵ��l�v�{B�1���gv5/��9�#�+����A[������M`�`c=R���Ce�y�1�
�bd�_�'l�;77U��6�|�c�b�f�Y�3�w���%$H1u�Y�-�ӓB���I/��l��Bg���I?��y��F.�3�Z�Q��O�'���Vd�h��91�$6�L�S[Y�����6wOH��7�c�c5V#��`>6�0�0O��q3��?���@oy��2�M��M�����4��b�F����	H��j��1���4R�J�U	
��[�|���� �6b۫�~tuP�h$��[�3L�c����:Ǽw��Ճ�������e�8-@��3��}��wao�ؾE�m����&H�0x�m3S�u�D�;��
-��B)g�N���1I^Hَo k3���\����q=ɮe�P.I����� ����te{Ѫɺc/P΅^|ZA
zU ����xv��=X�F���R�=��p���Ѡ/�Ų���xc#���?}�_2��c�M9 ז��T�*r�Q�=�
�b����;�3����?��j�SfL���ŋ;L�@�i��5hH���V@A���䅡q^���\�<��V��گ{�<7�we��x�tMb��鴰כ�PM;m�gx��xlܙ�!EsN���D���N�P�������=�ۖN�
���-La�F�إB	7��H����V��0��o[�b���lxj�u�F7y_kF�s��Z��i���O!lg�<�g�����J���m^8�ؙ���	���YT�=^3G��e@�� F5+��ۛ�9$�'s���¡��A�����i� &7/�S�=���\G�ǰP����^�--2�S��y����ʟ*�������7��nQ����l_t��D2bhN F
�9�zdA�Ɉ���6WH݇@!�H�Hg�.������#SB��U|��m��^w����cފ���OQ�����6F�,�F�͙�1�b��|�ON�/�pG/R��58�ֱ�ڟ�rB��(�_"wjY�J�����'���-陝di;��ز�S%���1;���3�l�*��';'�Xv�Y�J	�p��%JR@DWmVbJ���o�%&��C��1�f�|q��SҘ���s�ždo�1���*�wBl�P-����h�����I�������]�ظ׀��/h3����(����Id"�����8#��ʡA�p�}����/�O�z������9E�\SH)n�^s�u#�=��#vq�4J�Q��iY>[�J<;��W3+9Jܹ�!���A���{�2��8{q=�ޔ�By�+B��>���?�8�J+���(e��F�N��(�6��R�/@=�Ē���&py�GU�+��P}s|�Ԋv䳞Y�cr�y�~���T��	ᬐ-k-D5�r$ˉ��s�zWᢳ�V2����P�y G��A~xG�bŀR�̂hϡ�2�e��ǟ 7� �6�'Yy@��7�Oo,&���?�-��ڡ�f�o8 A��M��J}���5f�ӏ���\�CaRZ�@�_����|�0��L�BG��k���:J�e6�]�l���6�E	�f�
�4=W��)PJ�s��$��f��/��Y5~.���88��3��晝n٧�x��T��U9-���I�E����@�q���헂PA)MNyf�j=���S�p7��R�g����������8�xC��-���X�y��i��c8 �vU��A%�>�뢌��@��v�>���u�.4�rs�����'(��ӳ8�K�P��2V|E?|P��-UݏVk�-x荞fHS�CA�]���]J���I�VE�d�ɔ�û"!E��t�閶C�U��n�g�=@���d�K69����?��%���������� ~eqp�¸�IT�� ~�d�����\�g�>������W�P�,D{V�+^�a�I�;���y�Eצa{�~���m��4ښ��	[���s*Qi�͵�r�	 �GN 1�kN`��,���c�m�!�f���g��=j�ȎQ�'��VZ��[`dpAy��i'��@�I���n�Ȓ����)HS��t���4�+¶�G[����^""�rϭ:mnP#uH�@��
i���0���%�ڷ��m���ՆN���s-�C1 ���	%q��I.?C���EC�����0,��^�
�Z�����P���Ւ]� ��E�t�06[�$r��}� ��o��|���������F��|�hS��t�B����:�N6�m�\�������6K�b���4@YᷬE :33iki׾�C��/p$U�T�ο��-�i|�Ժ�ʜ?��]��<b����1bv!�ɓ>؅vش�7��k�E`ڒ�i��"����E�X�<|4�ީF��&]�C7D��Z&��/I�g��ye{�ƪ�^}��&,I^����gLM�����V���Ab�Ϸ'Z�I�,�0������T?�OKꍲ�b̶{�$���.��\�-4��/�]Iw&_�z���7��I�"�`m�x�Ǩ�#-�y��oɤ�0��W��ϋ?C���Q���J�Et�A���r�Y�{�����H�CU�6lኯJvB%�|ۦ�ck�w��c��'�{����5pиC�]���O�����*�Ig pvt��H���_QXip�9�@�.�ɶ��.i2��h=T1�@�J&%z��/"�o^�E]�^7o3_�K���m�ly�#��̩�9��pIWd�I�ݎn���y��J��i�sV$�V�
'�m��@!��g2i�Q���6 6�g�sG�Iu1�.Ӎ:Ȯ�EP���B�@H|W�v;���8�[;�u.xE��p�c�ǃ� ]��<�Qa�d+�~�����Z}��h����"[���G�r�(Fa	Q�u������PkL������(��p��{㝽Y�by�)A�f'�7rPQ���o��	^H-��d\��3T�d�v@u(��t/�O&s���������
�X��t�xo����g��38��/�a7��A%��'f��\o�Q%[� *Ot��lȳ����w�Q�x�a��rx�96������0M@ؖ3����ǷY�9�����6�3* �
������ժ�(�b�Zu*H�;�y(��L� ۧ����L.��{�]HU�Ԣ$v���H�0�A����4�VZ@���G��#c�"��2Z�c��a�[������]"t	/���0v�TP�Ch�uBL�,�����`N�������q'Q�о}��;| h�W&�����M)�3-MP���������p�;�e-�)����Tf�8~�,�/���	���ʝУ�9s`(�G���R	����y��J��:����I��{�DG�U���G�� ���^�U����;P�r[��b3{-�%�¿&3�{�g�%�Z�k)l�l��(Sѥ�|�0xaDA�� ���)D��G9��YP1fN'�*��®�^>����\M~��d�ׅ���bC�S��LU�)���g��An�X������A���wF�zثϴ=�x�Hȿ���:��;V= 'd4�&���p��CbH��0�yc��s��>Q�+$)Yh���������WBM�ѡ�49,�c��_K�čZ�FWe;c>�ch�F.�_�d����PU5xNfF�4n�dr�֣�;�7�&3A~>����cM,J�<����54�5I"�ݙ�2Z��4g�����p�.�D�%⃻��7=��Y�s��(�t�Y:6Rd���A�r,��ϙ�V�1���k��K�ҟ�h�8[hR�X� ����L5�-�M�_����ʩ��ԓ?�2�_����cU�7کz�ê�,�r[��9���]��>=n��NP.Z��ߪF�&� P�'�,���3����RX���%�xh�?ej�A��E�U����Ј��%�����3��Õ��8�6�^������zZ���{��f���T���^�.*&��\?����@��BO��P�[��Hi
���^�Í�aê���+��5_�2��:��3�H�$�U%}�Wc�v�H��X4�<@��h$�8{�������1&A���ѿy������k���&���8�����"�c�f�2��g��|qL'o��02Wdez�|���{�J
������V���>Naզ�WEx��ε�� Z}��g&��z��uT���8˟� r&}��tx�٢ŧ0Ή������;�58,n :i�f�>�D��Q��4���L���_�ѿ<W5D�����7��1'Q�����i����d�w/gas����a�M�`�lA���� /��:1؉��N)�s��.���9���ĦY����A`#�6h�}��Z���m%�U�(����!������T�$�()��Q��W~f��w�O��S<ޒ��WO:�%>�^�Z<Q�!c�܇��ѥ>Jd��?0�P!�|��f��x��Q�� ���B�:F����3�P��c��#�3ӯ�c`B�ؕ�6/��Ǭ9B4�kނ3��Q,3�N
�)��+�#�f��/��4�<���� ��z�╩�Ȯz~~�G���z�p�E�(�}U�φJ�m��@�
��"�����1�78�VZ�g�ǄEۀjK7��wu�>M��濷8y�(�y�S��x��i����'��r��:
�����b1)���d�[tLrN<�ϬN��=B� ��:�T�����V؆�3�J�΄��wƲڑhl��,�����zq�g�;�F\2\��C�r���hǡ(�U�"�x��x^�i��:�~+<�/�C?.=׍E��ڛA�Z���+J�I�6J- �������4�%~��^G��H�[�Ǘ�]G���V�W$3n=� I�SEXr����J�N|t�|G��i6L��@��.�W7ML.�GpaB�K!Dz� .RǢ	�U��p�V��Z��L�����?�^m7�P����W��G����%���|�Ȑ�vV3y�Q����K����x
z�@��{�z^,��Y��|�~�kp{�DD�P�ԛ3hxÕ��mr�q��~
\i�2�V�ѝ�Y@a���H�<���_��X���\m�Y������j�+��t�>Wԗ �CVe+�1q�g�U�f��L�%��{���$��(��#�l���f��}���
0�F�#�a�6Pp��̐����H2f}@�'� �*	�Gwg�z����
Ï	2�c�c�ܱJ�[:Z�%�YB�]��^��M��%w�N�y+��K����D4��8�iG:��]�� ���G�MƄ����X��Iz�ug�^+��=҂�� B�����Bs���C��Ko�}r�kqP`3�
���'ǆm�Ơ����y���`��⋩�����ؕS�vV�()NhI�(��9�ʈH����a� �_�y×���v=k}�%�a� �<}���C�w�&�m��D��Ð�%�g�!�_��:�㭡P���k!�F���=.��Ϙ��۔T?���χ�i_Ռ���Z8e=Y?+�I� �f��W<��T�sr��Ϋ�[��4zh�/��E� ��3/�|W�)��|c��2�&��A.��5.�_�
d��N(<�`W�V��9^D4�I^�YWh}�a�߸Nj��hҟmN[�Q�,��^1��J��S
�[�����C�h��HE������g1�����|��a����Rv9�UԹY��dnqn�X����y�BM+Vj�՚ou)�W����5?:+Vz��DU�H̉ �B�A6���F�=��&���YC���[8w�&Y�p�%�7�Y�� �a�逐ya5)Z{�v!Q�.%
Vy�����<�W�k�b!j�-�#|�:L����Gyƛ�1(�s6q"o�J�F��$���3�`׻wr�H�P���^�2���җ	�u���g}�iNԤ���:z۳U�����0IiA;O��q����v2�x��r��v۩Jf���o���n`�p�r�5�ΒH�����}���M7H*�w�ំ��nK��ך�UZ,+)O��WI4�߱���#�U���RI��V���~.��h���>�o�\|{��e�C�-��s6��NR�fE���;'º��
 g�)ND�W�̸��!o$A�u�����r��i�R��lsA�\������ n�F��Cc�Lz�k�$f��$�;5�.�(��x��@� ��c��X'�~L��+�[��	\���m�9�}���3�, $x��!� �B�N8ؔC�W֩t�����u/ sE��d���� ||�b��_>͖b�VA��ݕ�!�9tn�X�vf"*�#U�	R���>�=�-H�N��i�����*Jg��_�>ʈ�;J�n���;��Dz�/�z/��jrݑ�N�`���ۘpv7�I�T]���
H��F>�g�7y�B?�A.˩U-�Ӭ�� HV�{��.���G���)ۋ7�w��J(
�ʂ�� ��V�(�R]�gK�-���&�a�2�\� ׺��T��mq!$�������?�,�TNyrXb^j���D2e��m^tr,�aָ�0��Q�P	�t��zvx�oJc,7�����S|"�{��h���|6��8����������eYp
��L��'4L�opF�/�@H�Y���c����/_Zy�L�gs z>[M�����E�b���C6GY�pf񾇈8L�+1�H8�%c��/�����w'W�A��RE[kZ����s�Q�+WMn�J}8��4�y��j#�`Ud�pܛ��s�[��l�[���BNv8C�-X���2*��D��v�O R������%.5��Ɠ��lZT�$�`K���&1�]�QhrY���I 4Gt�Ic����H�!e-���7��9@���	���2��.��aS�-�����=��'9;��
J�i��kY������	�I����;�մ��Ӓ7MM^f��������Ǫ"$oq��w���A43��-�5��a^{��� G/��D����~�׎a3��iP��1�) y�@��Vh��9W��&6�(>�*� 0�];P��@�Ͷ{�Xx�k�ij��%��Q�3y��y�F-L���f�P3V���������)�¦��'��a�5ˌq{�&_�[c��Z�
N���D}t��L�!���������7h�A��=��ak��ƝI�5jZ	�}��p+��j�=���5�bs�bv�!��8�񈤭k�&¨:�7N�F���Q���Cr��/���&%A�	���R�Z73Q��{@���C��9
t�sЫ�H=�&��%r�ب��:lC���c�u��^�s�'�-z�[ �\� ���m:�R�u��i�r��C�T3�)>�M/�VHmZHF������P.����WW5���5�[�z���4&���s�@'Wb��N'{���*��������u�^�h׻�X�b`��m).�3:d���˂N�o�L�E!'��]� ��I���[�i^2��d�sI*�b��5P^�]��T�r��ڞ�׌�Qh#P�iVL��9���
,��2�i��P�9�� $�:-�){dˁ����.K$d
��/�����`��zX3��;CX�E��P��iCW����k�e��O@M,�s������`/���s��b��$�Qہ�2���F�>DU�~�a�O�#��C��$�9������ω��B��&d̈�3s�kT<���iB����^~����y����_�Ř��OD��� A�R�@���x��&��}&"�ΕX���6�v>��ڝ�a�������B�N��ud�z�sn,Ļa��,�F�8��
�ۑj�8�>M����$8�=<FMq �ݹ�}�E�R��Zf������.
���� �d9�lTX� ? ��ٵc�r���%O�;�pH"q�$ ����3A܎�ˆ�'�l�f��/��a��x�� !��Ov\��,`#so.5��x�M|�������X�R Y�R��`Tf��@<�t^�٩QLJ��G^1��I��]�
R#����q#����U�-��M�U �p6Ă�s�L!z��"�zXA) R6.������z��d���4�썥���/=:t�B:8,��.��~`��	\�g���-'k�7��9n�������A:�������/�����t�w�e}�h ���E1�B�_uz�8� 2�j:�78���nj�@�8bf�>i��l�:�g1��Uw$f��Տ��..�[������!k����-_�1=@��n
\SЙ�#=z���LQ4v���/� 㩬9��a50��C��j�(9H%� �б�]���O"�rM���QV:tz�&�ǡ�v7�����י�`o��2X-���/{L�'�:"
C�52ħiX��77����M��'Z��� �a�+\߄��Hsk�<ݏZ̓�s��y;F���Lɓro��[�3W��Kʕ#�ԡ�ӕ'|��a'��۩Rşg��Fl��杨�b�{�����UkzK�[U�����~ը)��`��9P�n��.-,z&�匎���'�1ƿ��#r)ȩ���+�DMQ��o�@!ۭ5d�^6v�j��B�	4�l&̃���'�`[��(le�,��	���]۞�<�}��HM�R�~�j;D��9"��zE�mkqY���h�v�65�Q�#j�v��S���I�ۿ��)ꌩ��Oi�XZYf�(�:����S�� �+",��%;G�m���P�>���s��F�NgbF�/Ҩ�_Hg�5@Ý)��}|����E�F��Nh2��a�S5���L�;�Ĺv5�)�b��8��2WZ��AEk\-�N�Y�� w�D�-�+"o�!�¤�bG����n��[�.�O��5���;@XR�pg�!V�m�a�S�d���
�j[//T_�@��0���xYg��"M:��?���ؗ��a��*���b��.Ug]��]�Ph��H&Y��bK���c8 3�袝���:�-z�lvՓ����Sm�:f���~a���Å#6�Q��K ڛ0U���[�}F��_4�Ǽ�/���bw���5 �x� J�
�A����g����7`T%�E�#�
�/)\t�"��׏*F���]-���cۘ���2��T�
w��P�c|A��t����߆�A`��T�2���h��}�l�q�J�j@��J�
�aav�d :�
 ���%�f@4�S���O�HĒhlh��w9�
j����_��n`�#Z5�����{ >cY0O̶��\�*�\~�!�.��A^>W[����c�}#;���r9��3Ĺv[�0o.�=r�}�������=}SpC��\wn����IA�`y#�ڞ��G�d��z�e!o(��l���Ē>;���u��"��i��C��fL1���������� SB�� -b�j(�c��j@m��=c����0����;M>��g��t��Ԧ�O�zCB��OL@z�&�R�����Y{��;�s0O̽�j�)b|�r߾3*h��騟ؐhgMu;>T�T�L������bK��?��%=��O{t��;$_7�d�$���a�\��<Fq-�8�d:��
5�u! �퍸�Q��uf���X_�k;��gm�b��q�.l��D�-�S-����,t����{t(�=�{E�QD�a�y�,��+���5&��6����cV��2~D���:��Ob,�=��b��-(p�G�T��h�-/X�g�\����AQ=p������:�$x����1.4�`�|hø��"1��ta�Ñ��D���]�:u�� �(�
-�`J��ߎ��TgӪ�]T�y��^���W/��լ���t�M�*����bȣ\ ����yӥ��m{���`�����JߧG-���P�4S��$�&�Y9��9�P�{��C���*��X�����`YCU�j^���>��V�)�tM�
Xp��������������>s�{ҫ�#��\w��ot�Ew�~��"��#M֠��U��\��hʷ��Ko�V�hIz��w���I�y���xa_��Q�� ��v�j����,��̾�e'8Q�Qo	d��
Ob�wfx�oh"w:b錼�y*؟7a�5�E���(3��k�N�4�j�r���x��ld�İ����fТ��D"��)��9�>�q�F��e7�2�IP�	��'g��Q+�]!�5��2�uHOm��]��r����Fu�2�g��u�:�R����Y�=��l$T��xo�TN��QN!Ԋí␪o�@��6�$B�S=��%{՚f�܃_|u�&D��C�ش�ٸ��X��[��((�z�{�2��ӫ�8�XE��PG�vGؒw0�#�9�>CtS�<ei:���*�9�5�@`}�j^�%V�0u�|���]���e!�I`�6����<�����<�����@�M�56I�<��.&��1�Qn3P���+t%���=
["��~
�KX����|��(FQ���6������1P<*����'=qԂ���VEs�$C�r��ЭZ�z�I(M�f� {��=ѝ�NC�}�:E�� ���i�λ5t$z#_E�<��|�'����V?��6���������I����v�&H�I���X�ط��:��Xc�j7�X�$;�LD�R�H-�MnJ�`�z��Z�?���)�̐P�H��'y���Go��������suJ��@�<����ק3��;`�C@/��%�f�6Ns�A1J�u?��,:����-~�x�Xk�YF��"�\����-Li��� �\篤Z�$= ���`���d�*h� ��\D����]�Z��^^O���^�)��~|﮾��jvӗ�\'u��Y䶟��#Cq�K���O`��C�9%'�_�F*C�}�|��`u���+�u��FrD�)��ڿ�L/�Z��T0�M��(�'���A�`�of],D��N�%\���*���X:貿h��ў6wGH!_�����!X�K�"OL�e�&f���)�*8i�R-q����8"8�}� �#E�J�!o�^�H�M�dY�8�mH��ә󱽂2Q"��)�8���S��-���;Ƒ���ӠNkz�dW�	#�0v������'���Η��\�ڸO'1�!:l����t�C�����^5CO���e}��w*��ȇr�-�^6T�2�������-�\ǽU3�{��g�D����#�@=�S�'rX�[Ԟ�TON���K�v�Q�wR}9֓����B�Nxjλn]E�E�sc���@/��S�ʐ��/�<$44��^"3��D�D��1�q����{t���s4��[U]Gu*0�؏��P�>EyU[&bۨ� ��",��\�_w����"ˈ7B��J�;��Nib5ek�c&��7Z*��\t�0�>��0�wc!��Rc��,�3����QQ��t���U`o뤕P/rG�����XJx���q�?[)�c��&�F`�)8˲������7"��Ѽ+��%��}��2\˓ki��i9"��A}������(t:~�&D���邋����fE�q�l�}$���#�6. ��l�Y����#*9�ZJ���=�)��‧ �)��ݡTpEal)�1���B�`G�O%1X�&a=���֯�?��%���z}��v3G}�����}?e �^{\}oH�ߔ.�{���R�����9�����D�tu��ne�Z�b`J�9����X0�{fi�%O�9�¶��#�8���:v0d]���ۍ$��<�Kk�5�3�sV�Δ�Z��m��Q���N�B�j�p^�zK?D�K����"Z�1��A�;͖�LnJ��f@T�a��Ԟ�$6�\�^M2%[.��H	b'#��a�8���nJ�t!9�*x4
�Es5�X�}�H���J)�R�]a����O`� �Ɵ����;�I�ͣO���)�qe�~8�լ��D;k�l�Te�d�懧TG�A��h�����")";�(,�D���i����L�6Y�tx��7����RI�[ٝGٻz�,Tڎ*�<[�gL����6���<�B���*UX#�-#e���k�lqt#��Ͼ�����#�Z�f�?/�ض&zj|����m�:)B�9��'�t��NZ5��/b˹,ly=���g�L�$�O?u��^o����\?���I=��?�E`�>/L9�&;r��������!t�+X�vGQ�3b���h��τAk�p��5�e���s�O������K�R�C�/�5�'m_Oį|Y�ZD��5GG������zv�������\$J��/�����jr��y�N����l1��W�6�tՏh?9���NF��&g��Q�g�{6�����{��m�mJ��(X�*������rz��0!2 m�+3cPy��T �6@ 5�;,2N�~\��{,��ֿ��?�����D1��~V�F�F�����'C��Sʚ;5?�m��n����jKl�Y�Y�h\�;M7֮��[.�K"��NY}��@{wI齂�w���5[�n��b[���}�M�QE��D��[�1�{`F�O�pQ��N'�'���=�!�2(>����a��w��kN��<I<_crlex��b�Q=�ܣ�b,:�۩"�@N���SmNpqbݰu��ƠB�+in�ְ�C!$1�*c��
��/M�O����8�L�h�xT����t/2��k���Q��WZ���a946jY�	DNy#�/���>�T�j�5�O��a�-�B$Y���Uk��l^)�
׏�S�Z���"a/�" Wf@�g��H�~��X�Jq�)Y�*b�a�%���"��꥽v��6>c����bw�9gwY� c,磼��zǕ!���ɗ)�&��Ǝy���-���.��V� ʿGO�?	�!uE�ȢBv�'C�!�<e4Gshn�n?���8�Pom�?�W���yb���if�`�\X���v=�-eNC�)�x˷�S�:��p��UP���=�t���r Q�Uo;���Q�|W��E�b�{�:��^ܦ��
���N�~�d��v#����$ؙ��"�@:���a��s���%�0TX�y6&��m��$�eL�ne;xݞ�OH^���󒳆����?�oxp���[9����-�X��m��]�ȝ��)�k/���e��)�.�{�X*ԞKq�TZ
O�B�0NH{ӡz��#�1�*�i���1�(Mmo4Bs-�l)��v�t�ӄÌԬ�dE.��+j�N��C�zأ5;�bR�ϱ��:)�b����oMnU���hfk�j���X%���R��9!��ϟ�О�հ*|m�	3$>v��B� 3��ɜ����qe?�>)�CmGdZ�����n-����M{��-� �8�@�y>�i�O��5�
�����]��Ul*���2���(�e����A��*�>o�	G);"~��|�䰜٢�@�Q��ŷ�&�@��5F���0�%f��2�,���&xC4�iNa	��Z�:�7����W���<��qMi�!�DTa!%�V�h�����v����j�l�R�p�46�ٚ )Z���tA��)�|��f?0E�ၩ���ȝ����ə�ϖU/RiVZuf��5���5�>Z�f���P	���18.}uMej"�n�d��D��h���IR(;�s�d鱳!h����C�\��#$��[�o|��&2(�;�ZR�]�T�;]$�Od�M�xv0��?D���y!Ǿr�m8G�4($D�,.���f5�����y��1cǇ:��)ͭ?"�C&l��$4��3�)�|<g�J?�FS/�Zp\� �+~�KU*_%DǓ#�+�Bo+ݢ�]j{�t��V^�O%&2�K��x�;O���sѵ��n�6�q�/��W��|a�	\��Ƶ�h�&��(�q.��A�l�LJ�+O �J�g��Y��3�1�^�U=�1/LȊpt�4X+Q��-��:���O�@!�3�qH��GF�/��6sr���[�ߕlO�-K�d��;�]����d]�#-I6|y� ��"7`,k�Q�0�v�HXDP���^~Ⱥ]�t���O���%ĝ|�"�;�3���%_�������iI���	���� ʝ�%߫V�JpuX�	#�㇮�����F�����P���\, �S�P�*������E�W H��A�Vg2Gj��z%��6�Q�;>@���^��,K�:��R.ΒA��G��l�{a�U�f��*?e��E����:	���O��pZI�M��V$O�nZ�׆��?�. �Ca���d�׽��������U���N>���ҮeS�򉤛��մh "��	��k�FM�ѠB� �"I���2k�`�y�߽��)˓��z+�?yg�'��1wk�4��v�;�Z�����J��'�����YK�ĉE }����9��P1��o�C��{�ٔE��rX��؊�7̍�-����t�JS���X*8�>8_
�#�wfݍ}��@w*�o�W1<��i���f��Q���e.X
��'��eN�W�D�o�3*p�M��I-\\ ���ԓ����nq���7�JH�H�b8�f�WD�2h��+@���d,�6����D�n��l�Q)J���R��ދl����Dx�W�1eX�C@������M�Gze��d��
]�-�!�f�6.ˎ~���~�	%,�+6��Z���<�wj>�Z�QRZ�r	��[;6i�M�hhT� ����i E�2î�c+�w��}���]����4(�S����-�����D47*�]R>���=� 9��ʋ��Ǒ��@=Ի����:�J�Ϣ��1�/��2��\H^2�/j�m����j����r��&Ή�?>����2VD���|��7�<B�tQ�H��ynq�of����o��b��ȤZ��# DW=�y�W��:流H�����';��7陕.֞�_����B;S����+0P ��v*1
�x^<<Ʉ���p��b��M~��G �\N��T��x�+4(A����O��"GT�ɕ�����$��mVMf����ګe�^�#��y��e���1�R:Hu{.���r� ������C���Ϧ���o}�o\E��������U�����JZ���}��^�ݨjZ�v����e�E����,����j�<z�P����ͫ��bt��1L/7\�����R�S����P�Ia��ߩ��6���ta�ӕ6�~j�'iA���o�D��XOg�kɟ9(es���^���v����c$82~?!�}M���{�n��h̀�V�yk��(m�/m�uE��Z��+aV������,/B��F��R�Y��sj�J�&E�v���rpO=���*\s���^
�1����c/����,z`܋e��ŢI�����B!A�C��4����A�1�@R 6_�ɔ\�'�[�>�(%M�n@on	�R�8Ѻ�{�g;^I���#6�C�b��#��K3	^9С�D�LPN�����ܨ�p���w��m����$�T�Z<�n��.f�C�G�q�"�̉Lɼ,�zkm)b�Hp���ڰ/��n�]A�V_�8GҀz��:m/�Υn�S2k
([Z̵������,��W��#:I=�z\m/ސl��u�������j����I�\:�4J^�O	󄋆ݽ�6�o��ǫ��%5Z�S�2��8�E�&���ў<�ȥb?[vփ�W1��lMz��O��K�¬�K�evG�<q�6�pbK���j�*E��J��N���r�	������RD��2�^�	���U�/��K��C�gH��U�����%���9�8��<�ô��D6��q6��t��EfN���}1%��\֩�r6��X�L#�iP���93>�?=oo��]1N522ڲ�ܪx��*;�U��B�^�;�0�G�'P�FTN)��R�fToГY�������o-X��z(;��i�Z��ԇ��N���J&�}r��S��"{-�[D�nn�u�r
e�u�qXq8e��x����a�]�ulŲmY7����=t|w���/$��QF��z�P ���@L8<� ���ɑ�;������b�hFt=�C_QhUn~�%����!�-�iDHES79���_?�"�`����q�N�x�z�*Fz��8��V����s=�r���H��5�kc[�-������8�H�N��`Xz�=���� ����v�h�^7������)v�+��
["�,x��H���P�����3� ��s�28Lp��ІI�G�긅�/������X&��-�%2���g�p���eO���l�8���\I8�țo�0�b1���~�2���4;\'K��/ow9O�{jڸ0ׅ�ǌ����G��9�+Je�|�T���Bbl�1'!/T*ԥ���)�gE1�be�wΐ��`R`w���-���<�`jXy��]�+W��G�6&�K��i~���F1�k�
�"<��Y�gqTα&p-^{����bp+�p�ਫ਼)�ʾ��H��	~�z��@�J�/��Ʉ�ӽu�82f	2#;SU#�L��5�/��$����RK�a;�z�#@k�e�Z �J����sZ20\��4$��2��?,��h�r/�\���州
�����HߞT�$�S�隌W�	3���tۄH������5�˛o"��`��vCw�
�XN`B��l�&n�L���=�T����Ꞟ�e�����4�n��ĳ��Ϲ [�8Y�G���Pr�Xhz���<����2 ��T�z�U��MR�9�io�d������_����N��ڄf��?>7W"�G(����	}� �Q!�4����Mљ�Wp�p�*��tN���[A��z�=R|�X�_�������T�`¼�P-1�V�"�E��W�:;pf�dZX��﫾Y�0�A?V�5z���#K��G�y������#S3�)L�Z�r�t� Gɍ��p������ ΁�u�M��r#�u��tK�.c�l�f;6�X�0�)-��$o�o��R�#��O�?t�SP��k�q�I��1 o�"@���Nu,�P��H�7���eUs��J#.5�P�^����f�=c�B��U�Ƚݶ&X�V&#�7����FD環��/T΁�Q	���<�)kKM;��9��H+�c��e2�f"�#ӕ�o����$&	)��m�w��V�=H�+=#;�߿T����@�_��H3�����h~8��{eP��؊�F��9����	���Dh��e
�3��ߥ���:��NN�J"�|�O�8P4$y�E壟f>Q��؆�R�&�;$v�G��̠�`y���}~�3��w������������x�[��F�d���'H����ܜ.|<W��z+]��_�nT��sҽ���xq���IxoGߦ�����+�12������83|Iu�sR��Ga/�����rNx}��ɃSoqҿ$S9W�v�C�"TU믥E�������P�Z�J�D-�Ng�?�	�Թ&�Op�#��=�+�XcyQ<N����ȵ<��[QH�
���WIc@Y�f�^��wƱ�K{�i�{�X_�4�}�pB����}�˦��EvS�
.� >�p���[��N�m��u���F*Q�I�l4�N#y�d䊵ҕ���4�.Um����N{(x�m�����φ�{ƴ1T+��i�^����� �%�W��!���C)^c��,_�{�,�ʛ�C�c�KS�F��^�7�n��5�`(����~<���|���IT�sT9Qn-��qཽ>]��s��2`8;'���Hu�j�%g�u�`V|�N9�{���mh#_�<�Q�~�"=�>�/N��,����\���'����IF�]���%)�dA���<4���l.x^a�0\�TTa�$������>=�^��;��l��Zأ��s��2���w��v�T['�%���^�l� b�)CJ�u-4���L^�VZ0���Y�Uc��f�eHu`�1%!�9>�����/�7qk�n.�j+��ѓ�E�ӆ:��3�����UV{���qQ���vey��>f��]�D�N�B�l���")�'�m����.��U�99��޿��s4#�3�a�چ�I�Ζ�	,�x����K�}8/��?) �g����\�<!��H�`��Dtk�8IT���с��6-?&�����]��d�]��|D�����=�-��F^1��*�g)��s���\�e驖��<.�E_��h5Q�u".�$v�ĝO�����o^����tW,<�&���}1�����h�%����b���$����P�9��Q��8��P�!�^�UC��[u[�͠�/>o��[o��I�,�I5�̔yB�U������o8d3�R��Y�"�bt�-��3r"��:��/%9}��e|���[�&��"CP��X���i���7ru�J���v��.	�2puI����'�\���Y��p�����x(���戩x;bv� d^�f���E�$vI��TaP��i�\.CD}r�#L������Q�ZR�~[�q2�/���p
A��Ջ�j��O�>)�³퇶�q�׎����Lu�"ZgD� +�q]��w�*���{�d�#�u[�<7����d��(+�ٯ��H��dXm=�G�_�������X֣��b� �'ݧ��>3���۟T�G��1�7��Z��R�_&B��ͻ��������;F�3]5JOP^�`]VM�q�?ӥ��2���7>7QL1�JN32�)d�l:�9�,
�[�i�g����@e%�x�y���=4�������7,>���B;4I9	�7��h�(�c���rT6+���L�M�#��`ף���^�މg��$���:�7����P�B��b��oP���)fD����_e�.�x��K3f�e�	�� @��<��]��@�W�m��&e�>�	��z#zu���p�]�"]KnQ�7��RƳ<ʜ�q^�,:�>�QleM}*�R���]�|���bX��S����8H53^O������\�߀`.�-#�ʡV=F���e?['^�7|�܂��1�D�;W�-m3C�6�K�<K*��S_����#���F�<Ya�J�������!�Ɩ��t_Z�I�D���D��
������4�P�B��*[��}��t�Ӊ_4�k��d�IZ�:Tڈ�BG��M	V�A;�ϐ�C��N����*�<����)I���7?��<w�¾�ܩ��0�)�o����(8�x�ɰ`!,́��<e�.��}M��e��6�iR�q��<A��i�,�`�{C3�25M�lp��B�ic�cC��<�]�o_��dh���P�/G'�`�����Y�/��q��U��U�H�;)��tA��P��Yɵ5?���Ň��L@�JK��!�ȉ|���A12�/i�m�H5��uQ��?I>�o��{)�j��k%�-ԏ��`�}G\4��|��['�eM$�E�,�O\���	r�@-G'A1Ę��=��j+��f��7��*e�w�����u� [B����zHy5N�9 _2K'oi���((uY݊C�	ÚC�¦J_��OV,�꛲SOh�]��*�J#�+7c�X��|�A/�vx2P�c��?)��������L�T�K��w�I �U3-�h�f��Dշ������J��ퟘU�������IB���|�R7��9�uC	c��?��=˦t��2�;����EI���]6]�>��/��_�J+��]M��Y�R�d��4��<��"*^\���JDoS���"'�gcA;�-�좜<�x(Dk�2�d��;RJ��o�i��a_B�Q�Y�ԲX�fo �$|)�(P/� ��/5'9�[hSz#{�G��:ca��
fw��-9}�mu���%��P.�k@��
 �����Nt�e۷�eDG��!�*n�K�g���ޤ9�Y�p�C-��`���ם*[�?��G
��v| ��G��a�����l��y����I����l?*��&w�P��/����q	)4�`��B��yH9�k��a�"�{&x�lU�h8�l{X�w%C�n���i�yW�{c�G���h\����#Ug�޾y��i��D���"��ܵ��A�$ց�g�"�99a�S�����<�T@C�xhj+�pa�Ҳ�*���F�(��&,�\��@��ȫqp�! gN:�b�9��΍�["����w����ϔ~�`���=��s����H�-��-c&u�����&� ��n�����y\�7#���S�.P�p=�xY5F�p/G�rq!Y-9�\F��F���)F�{v/x��j!*B�ۉ�$�����UY�S���3O��+PrĨ2b�뽌J�g�����j,���Ų�ʖ�Ά������H��������Ga�������u�AR�Ar�"�r�7Ǔ50D�n{v�x� @lU��I/�v���A���C�=���A`�I���͓���~x$�xQ!�53?�j~��������l#��*�����'�T��������<m�(.Հ�l����]{s^׎.�?&пr���m�#����s���Չx�uOGͿ�f��80t�,�٧��2W�P�.A/�C]i"q�>�{��)�s�'�=WV}���s���)�����K��Xc��q+�V�.��<��b��U/���.o��8�tm�7ۏ�=�g��?�V��֟���������4<yM�B��'_c\"暻w�+Z��?��U�¬�m��MA�B��ޥ��|�'��@�./�B�)f�xI���L'-���^z��u-1ؗ�Ϋ�x{�}tc��ڌX'�.o2�hvga K��xa��A��:���{�#��Ҝ6|��w�� �}��8)�'�˳1>��
�%O�����}�_ڂ��)����[ic�<7�Db��<�J��� ����l& p�u=�LLxxK���>9j�^�B�W��I��2y�?���u9��f�)Z�I���=w8���3LI}�F��