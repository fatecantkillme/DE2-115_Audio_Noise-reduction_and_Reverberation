��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��&���i} Ĳ?���3rz��I�{��1MZob��N�X�����0�D�ɣO��ad�U��e9�3�f����Rxe����U��S]#	Rk�ݸOq��CsL<<��?
�[E��G,Q��TN��P;�Xlr�͘դR��[���%�H����RS�u��b^���	�������"L�\��q����è��F(�O���v���F=�H�<I�DZ��d(�(1U=�/���*�إ}�,�n7H"(��2����bt��ZW(�5+�.W���g��0P���N^XK�Ʋ�65��0۾�@u�]��"�	��v���!vg�	4ś��x�WM�yWG-zvP#�y���e$f�r({��4oVh�/]	��}�k�M�(#�6��z�U�/^��e�k���y0Nr��EA�1���!��46�����4�=�>ǡ@��J�p�tx,-�%��A�>̸��
x�
��?A�v�c5����>]�;�u�ۄ�mߖ�/j�;����]Nw|桢�v��=��b���NI�B���5ND�̜��&I����� ��������
��d�U$�
�Wp�nA�bJ�W�D�Ԣ�#O(����Y'+s]b>۳�#��Ьʚ��X�h�N99�,pjA��.�>�iu��nyt|�RʞZ�,O��R�t�ĴV���]Iw����#a�/YK8����8-	������b�a�|N) o�x!l��dmt�f�<���#򂒂��s	�z\?`9��D�Ή�,��X���?r��x�߭��u,���O!j�3U��+|�y��.�<�k��\��>Y<H��5R���e]�F��sS_��8|L3`��x��2q�+14�6xH橺S�&^����ڽe�+|�(k��(&�P6$c��Z��UI$���-����>�`Sk�0pC"8�X(�U�j>��>����i�"�����=����gG&#��6� k��Go�GN^�a��8�� .�P`���f���-|%ώ�;[>A��i�3�*N V)����9c2pPm���������ܤȩ���[�K��>d� ��~Ih'� g!k���5����>�Cꮖ�(n3��i6m��<|�#rc�5�kf��������B�1)���f�q��ňg���(�S�/�nY
�������R#~�Y��� �4�h���<#V>��|�i�¨>���R�6A1��2[��o}�X�]��
�>�$|>Q,�)®�Et;��C�C�Bx160�My⩡��;0X�o�iW�X�d����iW��z��iC��=��8 .k@?ŢӾ�F�U?�ֹ���2��n�ל��o/��7W�{>��A}��8�C��1I[�;�[a~' t��	:PwR�/�[2}��L4�( �N�����#�W�Ǉ��}[N(�k�$��m��j���8�y E�Ⱌ-��E%~3�m�q���5�X=��"
�3j8�!c�G�?�Q/�+).�Yf#���
c�p��Fe���D���ϊ���*UM���ej���<���ȱo"r`g(����]���\!�<׭l��r
[��ET����wv��r`��fƋ߻^�u���$J��3�N<Թn���;��>J��~���W�qy�fH��G�~"�X�yGs%,U��4�-8�I�P����Z���X�Y���tryq��K^��p:^��q^�d	�	H�"�{��p���	��e+ ^�$Q�<c���$�	n�:� w�51��7)��#uB-��_>��cY�׹��˩��-O���c�2'���z#�U�Z�G�Qs1��Q`=������]b�q�})�t��`���$�!�X �[�(���"�!��t�)��,���� ������#�J�L�6v�������С�{�6n��}J��`������:U��S|��y���7S'zFwVB� d����_�C���|���TI3m�i���]�΅��ɻ%�ˈ����I� �� ��}�N���;�$R���3�r{�͜%�W�����0���x9X�MR���C��7�_�	%�>M�:�����3o��Tb*U7�s�8d�� ��I��N=p �����b/���Z�7&p@nX{�,�d=Č����Yщ �`r$�E���Z�7/���Z!jC&���%PB�p�*�Դ��_��g����^H��)_,}�DT�n�.�r~�}`��?T�a��O�E{��u�� r��3��8v��+�L�°,"��I��FLS���d��k�s
@h�ɠMd��G-����d�(ڃ|۴zۃ�����<��+�P�ksO��.&-��T��V8��ƞ<���\$��}�>]�v�BǙ�/�b�T�<;A�����d_�"����1�Y�LL"����v�6�T�D��%#�%�Y80�5���aA���BP�B�� P|��C��@A�rt��h�&mȞ�6,h��y���
ܡ����wԣ��81%�;{^rx;��S)���iZ<=xzg�z��I���ޮjpL �n����+"-��+sl������W_y�����:Z-�6�ؐĩ�컩�KNz߃�m�ߠ?pFo��jL.��9Ju	��^��<š�������&ݽ�5�?�)V|h
{�g��^�r�eRQ�G��P�˱�S�� i�f�ڱe��5��t3䲁�.�`���vH��M�2�O�"��D@g����a ��O�w�ݤ�vh��� 'Dɧ�qVwf�-�[��ķ/Y$�8hex5=�{�� b� ��ݷ�a(}�4C���BNhd	m>C���E�$(d�zO��E� �M$�����9[_����-�����<=���Qq�p}_���x�0^KC���(p��/f�8i�� �K��h=���۽#�$�N/Ҫ�(��/�o�O^�xDwG����Dt�,��>���*����\��na���R��й"hk��9.Vm^�U�8���a�$��)���l5re����Ȩ���G}!,bUU@�]�7B���E�e�D���t��$Җ��j|�a@kw��,��C�Lcא
�)��@6B���9LZ��́@��׋�_+�}������[ԩ���+d H]]�E��#p�횥W��)]c�w+�zeŞ����SH������z>�:�����t�~��*���3aK�������)D3��T��%GU��Rtw�M��-�}^�m׉�d��P��CI<��i;�4ؤ��=��R��ql �|��}�a����''gW���S�YCP�b���=�FR�b�q�&oP��qZ��3�P�C(D�8��@?y��gg4e:���H�鱒�����4��ූ1�NI��!ԗ][�s���wb�h�X�U�ԮЅ&�4s� `�+nVϴ#��um�>�#�9��ʀ���wD�^����mc��ࢀJ��a�k*,�B��ͤ���Q��	�p_���ԣ�R#�+y���4t%��(AKAv?m.� ����>���A'���	 ��D��}t\(�\r��Đ�h�'���i�=����4�L
��A�ߤI5��t��ԷA�h�$W$����8˚b���N�T����i�6!���e��B%�����Þ5'�j�wr
e�c���N@��ZO�s�\=~.�aY���o�L2ev��ݛ=��bd��ups���r/ܸ�&q
u{?��ֻ>���"\��5쌠�Iij��ϗ5Y�>�&(�)���l+���T��4d�[��.O���6�/��g@�xk�j�d8l��w>��|�[�{8��"�3���,�fXɁ��u��i�����7f�+ݬ������� d+&�'`S$���f�x�ugk@fʺ���W n:��a��o�5C�D�9��#-ד��Kyd�ڱfb�:��>�`�X�B�q;T0x"�z�K�c�
�sHS�~�5�[P<�LK��~���O��x�J[S�����`W?�]��6���8��a�������B,)k�����n���c�MC�Gn��e�BUq�}53.�n>�%������.�}h�p�T����PP��$`��Jۆ���A��+<�{��~��|�qq��*���*�WFq���k�X��`�%��R��ҳ��-�I� �w)��Q�e���~����h^�"%��
J��Z��;nʂ\�l1.S�oF ��^���Sd��O��.�)c��8�:~�t���i��v�t�}�� �6B��j���2(H�@���ȥm�\�3H95x��Y�M���1WW=��2��Vf��R���\��C�;P���{Ϊ���̨���_
�?�i�J9��o�~��ۺ:3f�{ܯ�C�
$���Z�Pqj��^����ۣn��y�+��/�(�W3x\��~�7��FW@�a-l�]�XƇE��U��od}�~\Z�d��]Q��{�R����W�v��(�ˆ�{[fR��0m7*��� ��uͤ *t�+M���q�];�A��"�r75�=�}�q`&�������8�=�O�Z��*N�k���5(�q�C��t�|R�&w� ����1��¹�|K!z��@��od������\z٢�)�?0�:d� ���r����{!�\�c©1*8�	k�1�a���f>����5l���e�Y2D�aS���69�ԧ�)�#sǳYs=.^WR��֤����d�̤ѥ3�SYC趰�0[ ��%�^��ˤ�uy�0R�J���D��g6�"皧`z�.t�.�/ot0�#]��r1Z��r�a�-��#�牉M���VR�U��o~Rő��7�&��,K!e�+��Ν�">��	��Z��	�(�yW��[�N�k�xw�XK�+�`ڱ�P���2b���<K��]�^T�h��J�^�#.n)�$C����kL����p�ת�NH�m��q.DUW=��.�qі��{�*=p�ťWF_����&w�<�S��]��q<1�D������­�S6�%���K��g�־�+�P��O�ѝl�L����א+��z�[漼B+k �9�&XI�4�k܇lF��G*��t;�!����. *藳�'��4>�}�%�|�Urjg���_��,.�˞�ё-5����p<�SM�Z�wC�vۉʿ.wB\HCƒz��]�t�����i��� n���"����.q-X�ks�PT:XfՁ.�q��m��F�c����+��u६f���vz$���~�<w���E�~VX�{���̲�:�l��~�M��5z����ݣ��]��l�"(�!I1������n_Y�FI\�!-	EF��b�+d~��ܑ�"������9���f��*�V��7r��H�[�jv���}��D�7�TrUY16�A����C�>��$\�B
�5�nq3��O)��wՉ�v�8ɦN��b�(���R�f��*�պ#��F�;�P3�a��~�ĈY�N�*�O��#¹Y����_: w�LEV��e��b�Ҧ�f��8�jH~���<	I1�5��C.���=��1'^��HsB���t��T͗=����u:�b92�F�#6릭^�8 -x�;�͓�	%h��q�JV#`D�gw:w��3�!�cy���;6\�Z���9�r��>���8��R�Zҩh���Ֆ��}=>)�
f}�Y���S��L��"{I�ݭ|�Up�>���(RRC��R�R��r��ќp��Ye��qvæO,������y�|�{J)�n���j���@��D�g�yOs}����E�f{��E
>�Z4��?h�f��Vz�]Y3z%��X�k�z��~1��cF��N&h~O�i����hW%4���M[ث�J�f�\0�^;��N��!FM:�~$��tIөfu&���".����0Xs�Sq��k�x�Ұ��4<;�9XO��}�Z�'��1���p���P��=�.|����`�����$gJQU<���<����� 49j5�!p���N*Ֆ�:�B[#�x��d��_��!s�W ����N��H?����y���[ŏ��Y|Sk�c�B E/!8�4S�����1k-��`��b?l�Mu5�MA�Ý"*ֺ+��@6D��?��E')j�')���U�;I3o�U����Ƹl��V��g;g�y�T7��d󑧴ybڭX&�����"��)Y�ɒkv3Dz�	v��?��`VU��[_�m�M,���-Z%��)%�_� �Anpn|XB_Ђ�Y����r�I�&#��Ɍ����>z��q!�e�u�vJ��K���4�O<�0\c΢Pf�2�>���Y��Х���I���K閪�kXXΚ�2w[�GC��{M��Ftz�ј��@*�K��͉�O�y���0|��i��ۧ��  �ɽ�C�Ŭ��p y'�=k���娏^���^�=��N��&Y#�QPbn4�_��3��ԟ������t� E�,QbgSq���ߧ���x�Ux��֐G��@�K`��RBJ��4rN��{��Wr�p�`⏵��6��+Ow+!����n[�8��򦁰��IS��}<�j	�A�.W6��.�8�?9jSƇ�FoW���^�����r����?����S���G���䇍_��=��k3w|ޠf� �1�J�O���;�S����k����*���
������sV/z�s(�w#�&̘�E�ng���냖.'LdY��	�%�y��'�jD����DHA������[�[]����8��3���BcٱXP����>�Z�y�����P���hm��:�TGY���s�6���56��G�N[��B�zw:���\�gM�"�sVQ��?��EƏ]�&zI����l&�.��'�9֪���⠷��˅���|��@�<&�Ƨ"%g���`���H	u� G��X7�_�6�9�t�@��t�7*���W�����vp���� ��/|�I
C��bᦚ�dCȂ	�#:�3�m<�嶣�-�U�#"��\�?<�I�aN1!a��Ã�u\�'X����~dy:�D흪=�H�Cf���g��͵�Z2���n���)��(Ry�%���>0�4�jj��/b]g1�c��,���2�ǁ(��m�r����c�o�v���B�ƄU�ٕ�DWF�w�����>�K����a��U�?�8cp�c�Rr��"@�^������s@�P;��Nھ����Lc��u���"���9���}	�;���Z������f·C9��{܏E���y�2	\�Gˮ�g�M �H|�xĞh8/]���	��d�����f8�\q�!ү��r�|{v]��V̶�e"�3o�)PQ;������B*R�������Xm�'����r�&v�/q�&`���B���¸:�3�����h�~�8F	_B��=|^��S�=hQ���RS�ho�� ���yHx|�/�r�+�p:n<\��0ܵ�ATN����iW]���� d�gD�Fy�kl���U.'[p)���d�S�|l���蚴P9uImp�+���"mQ�>_��ij��}\�USm�' B�$��N��L��(�!)?�j��D�t���0�V���p[���w��%��8&�o[��g}9����x�������S1����ͣH��v�[ܧ&*I����WQ����w;u�o�<mS���|������`�S�xwS���Є�|�{T�'KI��,�2͂����6c�#�̕C����dN��G �laG Ÿ��b����6(�I�jF���'�ɛ����E*ć�U��"Z;�Yc���uϷ5B����ܺ��y�Z;L��<���oȑ~��U�t���Ӏ�e=�bNd��������6�RJ̏[�� F�[(ώ���z� �����.[}au�to?.�Jȁ�Sj�a���K闃F���C��lm[�Խ�= -̑X�C�3f��8��L�����}�P�ҵܸO�B�!\��7���	]%���I[&�qkl^�jv1��֏�����e1���(0��bj��zj�4�BD����ҿ��W�]�����!�]m�Qn���M�)'o�N���[�z�O��t�#6ol�n6�4�
��dKօ��G�1�?��g�_v�uk�Sn�:��h����'r+�/of\���l�ձ�ǡ)�-(�l�9>�H��5�l#���"���𑔍��k�ŵj�+u��ۤ��}��b�X�U贑��������-����ʘz��#)ӻM��j����z�!�Hs4��D�����#Lee� L*x=�U)���$L�u�V.5d5�I�;㱱^���F�̡�T7=~�*6���sw��A�S�R�G=�0�eN��b�̸���GsGߛ �Y�l��^ZO�_gs�O<*k��Oc�x�0�s�}ɕ��q��������~tk���P%��Ap�Mg�1�D�P���w���w�_��Zl]�Nm묉A��3{!Yzϯ���t�^0�C�,3�M~����U�+�h�@J�i�u����u��uU�P,T�ͻ+>�k�#_�~N�rn_�*%�̸U�CfTr��5��n �r��Kn~�aĒ �������"���;[��T�K&4{F�H������7O��g�u�<��!�yr���+��b�q��h��Q^p^��>���F~����
;8J���ŷ���qs[�pA<B�.w�����k��:��.l�%XA3~���Dh>T�Ƅɐ� D��	x��:ٻa�o"����c��bu%ë��!R]�$G�vvC���� fq�A����Y��*	z&(p�'��M a��K�u2��� ��.��'�j��X�n��ʈ4ʬ��j���� T�'�2Mv��n^]�a#��K�30�a��Sg%&^�1*����Y��͂ɞSy�4d]��]]��,��G������t�'I�RuL�r�R�M�3�eأne>�Ӿ��e���(�������~�\�����"4F�5;�s��G��[�`e�AM����e�<wߠ��+�:3q��
Kz���r�-�v;�o�����B��OϏ��lO�Q��m�|	ٺ��Ss	��k������*[v@�9X$�o�-��j�����OA�nmG)����u�����ŕR�����7�|[%٫�[������)�V�4�h؟ٍ$�~&T���ܐ�-c���L�_�r(�D��	�v0�!c�:	Փ��Z!t5r��8	�)'�	�یE�80/chMа�t��O��$JR4`��j��	|��">O$���5�)V~$�z���q�#Xa<�İ
����ِQu���B���j�FyPP�>�
	Sp&M��k�~����ˇ͂?��LE�q���#>��U8wvؾwt-߿�r2����r�}=�9=R���(��I|T� u�.���J\�'b�J�PS-z�ij��(!�F�5C��׋�[�l5|�J��_{�E���
��z9�@
�:����'�8�ٸr��JC^t��<���H 4�[�#H�aW�1n2�/�������!g�P'=�P�,
��!���g "�K��<�u�� �SWa��޲��h¶�U���骥�r�C�=�9���a����7_~�Ғ���r�ˤ��5�4ӠS�MvФyID
 ��� s����n<<S޸(.̛���~�mͦ�G�2M^�o�.�F!5�(2q��[�����{d��/' y�oy]��md�C]�W�(^[�;�7h�5/5=�Y�$x�E3�H�&�I�8I����}Ƴ}��m��-��Em���p%h�/Ѐb����k���������q59���7ߠ�B�_�}Λ�؍�h�[Bf6u}�ҿ���w���E ,��'ep�3��੫j�m����mJG;�ie<�w�`�B�1�����jLd��״0��	�Jr���\#s� 0�-.�NS��A"TD�K�H��{+C��_z�P	#�D�B.����y�� h�)���=���&2ģ{Ԑ1�%�b$u?�Dr4d�~�S� xl�3�ėx�W�]��v$�d��F��wT�܍�c�2%�>Px͕�8,&�,����!��$�H����Y(Ħ��:����o�Ry��3?��L�݇�Q�<�]�Y��
�W��%%ti/�Y��
)��o[x��t�[gy�t.}NJ<��߹iդYJ��<$g��h)]��Iԧ6
[�^v.)�c��f�^x't�7�C˸0�+^�)�jP9��ظ��d̉����Ru��V~C�P���ϙP��Ҡ�����$��;������Kz5�*�� �[��4>� j|M+�30���f�(s �[6߷�O&	�v�lQue������<��S��[�gs�b�
*���j����̷�[�&b��+�FLI����N��ayO�+��Z 6��M��.���m��'�P�,S{
2�v���b5F%ZP
���i�G�+	�ohZ}������٥ZP�3��v䋨�#�*P�f׃����%�bM@�!���3f�H���F}��w#oé6fnl��[e���P���sk��Q��+�i��.���QMױ[�ƭ�J�JE�(����o����q����ݾ����쾃>���.x�^'�a����\�1�tY�%�֬V��HN�`��B|N����v]�=�Gb�E�F��W0����*�����>���7�ڭ@�iyjG�RH˗��1�%,�>ԋ`ϧ�o5�vM�#<�j�R5,Q��5V��y֯�1F�ڱ��U�@���{"��� \�9����Kw~X*�-2�5��q7�JI?R���r�2	�ӕ�Ps�Y���lhiG��. �d�.\Jڲ��b�|�/����H��.�rP؛��~�QlQ%F5�<�LiP�}f$������ ����A��l����z��Bv��Hp��p4 SnA�z�q1�f��nwF�(U�8������܊�{�t ��T�?�=u�rdcK�bܫ�%\���v^�4��S���5�h�L�5�%���v�M�]���E��5}﫝���1FH��B�$J�62Ȓֽ4tx���M�R�u���_Ը �����U�J���@�Jk�v�l�G:qu�}Xg叟?K&��'f0:���LP��� �W��;��|���ߡ�Muړ-���Er�>���㜛� �ր�u.��G\�Vz�J�Ӄ(�"���IJzV��m�Gu��c���"֏�.���{kĉ���5�'�A/eym٭�mqr��ȏ�t��Eq"m��k�W6Z���@i~�0)-Qn����F��d�lg��'E�����FשA�FИ����Y}�.���2/�#U�z�o��윦���".$r{k$������|SW'�Jâ���#�Uӹ�A�E���؏���(��jY�#��-d��\�/�©���H>�?"�d0\�c[PϞ�A�>�c���[1z��a��/��fQ�+�=�7��頁���(��>�*����OO!:0��B*��oba��gQ�`-3���6�ղ�&�R�����KA���֨�V��]��p;~�݄b~(��蠜�����1���k�d�
�zYY��^*��������5g]
�h�M�Q팁?݀"?�0����@D^!�[�:T�<���t%����_�2J�'	�"��p[��a�c7�I�ڟ�,�Rk�<��Y��!���xZ����Tcڒ�F�������Gw�V�Dy� m�I��k��j�"cM���^^a���I�̣��	K�c�Ҝ�������ճ�u�x�/"҇h�%}3�|��ah51��4~��R���e�\;q����q�
`�IC@�U�|צ�$��y�K�|&��oySHc!�b&�����o�#���E�������*$�I��μ��-뻔��bz�3�<�y����ަ����c	�/8sވ�d衲�ԡ�6��g9�����<#�!	\qu$��y�/;hSB
^�	@��{���1E�r�Ӧ�+(����$�m�8)����L��В����[:�Z��}!���
�>��*�`A-��u�t�W]<>.��fJ�?�x3�����}avN�^�!��ϭ{Z�����}��gW���Xt��|&'B��젴�'YO#K�߳���'�d�O�� h4��!�	R��4+��A5�CF�Du{���!�b'��T���H�� o$t�!`=�=��Rc��%}�/�ZS>,ec� �Ǒ�D��6�fE�	����;|2�2���JC_!��9%���wr@��k*�m&kv�y�r�_�~���;�2>v�(an����	�;�*ۈ��L�\��� ��B�B���-��0�w��7���N�<ٴX���4��R�)�o�^J��n��g�܋H>���0t�τ^T�KƚS���	����{�[�[�1d�=�.dX�>�f�Თ���x�$ʣ��θ;��k.~iG-�K%7x�%鶝��H��e?���&��Yփ�y���/j9߬>��@��� p�t��U̮��,�&?��$_���ݻ���"q�Ҋ��iݩ�ݭCrN4L��jXU?Ei��ցn|���fG��L �p�����,c�	.��9p� �i����+��&�j�.�;���l����-ȏwYZ�U;�h|�剺��6�搂D���eJ��QSapT��I��D)'�]��!�����ָh<�(=�o!�H%>C7~��]��̂��xE*x�d�e�gAS����Cc��:�ҩ�q�G��� �^��tk�3����[��'rK��@���nX�Z�=�R��W�8������� ��V�=�	c�h���q{^��W��ɝ�����ߩO��B�(�̌��Y��B5���I�ygh�C� KTaUb�g��j駵��u}��u4��C�`Gr�����m���o�������Ǩ{��WN �X�G�K��4�e�pe�n�%�M���g�ci�~�ɶ�ե?�1���ޚ�>{�?��U�ԭ�n0�]�G�@�n���AB9ܳQ�?U�6q�+�C��ѯ.�L�<W��9�ӷ#E��>]\76$rV���5�*}�Y&zI�W4t&tb��RcC��)�d4,�}�#ԋ4]-��,)~0�_�}ѩ��)C��Q�.^�M�)8��L�7'���n>�D��.d=߂46���� ��n�\�?ۑ6\\j����W��U��1d�Ɛ���ի3�v�a�D�K��ø����2�/��ą=@W'�W��CD���W��֠t��8��[X)�B�a?a;)V58�(���%@1z$uR�jN�xS��5-��1���i�'�+R�:)�N��Q���k}h(iε_��e�E-��*HK��1jE�������B���M�Yv0��������mf#	 �3a {"h.�����g�E�k��b	������Y�nI��Y�Ѹ턁���?��uKk)�5x3��"Y������]k��G1�_/u�¶bcک(wBO�"�xV�pg��XHV �H�)~����U_��6����ݕ:��|F��%��lrQ��o|	|JD����ȋk��qux��˃������ ��P���/3�e�l\�����;_������l�r��쌒�VccQ�D9M\3�]�)�U�1{h#v_1�*N$8�<�����Y�)��*l��]��&d�H�_��9ب3x�SX��{�D	y�F��k3'm\?l_���w=P��;@�$�&<���^<��w��o��Ļ�BΊ�ý���
�.�'#S�rw;= D�o����P,Lf$��%���SP��|S��V?o����s�#�斸��t��������r�Д��9�|2��$WoU�C��j��SS���W�Ch����	O�b�$$l�R�[�� ���'�6�����L�i�	���۱��|��\Ы�q�i"�ٕ�v�/6��7Gl����\�W�.�U2��N��?��D�,~�Ƃ�(
0)���w�o�v'�ƀ��<��2/�j]1��A]�nq��!��l�2�]���@˝Թ%<m5m���4M�/*v[
-��9z��m\7�Z=�����һ��<mk�����Y�̱�cQ�t�57�Ҫ���z~���*���M&�C�H&��F��:r���.�Q;���փkԌ��)���˫�ί?���A��dm��W�×� �PĹ	�In���:�à��� �(IS���>��?p��6dU<@��F���i��:���?�<��$��5z!�������l���� �F��6. �r�X[�4�P�;6Ӛ{)��30>Z�m5S���&k���LGC�ѥʧ`�
���5�߁�s�o�5d���ܒͿb#\� ����Eq���t����`��B�;��|��!��|,�����O��O�nyA���}L�?N�����i��D�7O��d���eU*F�	R�XG�U���%Ch��v讁 ��ܵM�Z���"�;_�����$�5v_���NQ�]%�X,�;�g��Ӡv��ފfh��dq��S�G^��{��pXM�{��ҏɈJ3��@2$�� �*����ve|f�F����Z�\������G9��U����ܵ��[7Fp�B�>�>�un�D�� Yst���ft]/T��*�!��FnY(O}��t7������ɧ��Y��=NG�>c���]�q�Y-�����p�h�zQ�"�32�X ���k�6�9���L�o��o �� #j���9��Ɋ��3˃�&���
@H�RŊv��vp��׆&sx8{p���{Q(��^Ȁ��k3��Rx�و�\�y�̆갣�z�س��M�͊G�9U��V	���c��hr��{X�Y[zY��V82����k#�~���<�g^��H������N����\�P��I��ų��DE
��c�X|���*���`�
��*`:�z~��}־O�#ނ�$����ۡަ��\�8�$�z�^$�k*�*-�.#w�&�,��3Yʜ����N$����:[:�u�[�l�e��& *�� �a��;+&)��ؿ0�V�O�;�Ԩ�P��;
Q�#���@cvCN�`(�e<[8�s�ħu�t��p��2n���ێb*�}���4a�vC��^a�-X�K
@���&�ʴ��?d�8�!>��z�����.��X�N*��x1�T�c�j�8�W�Hd �%g؜�Z��<<DQ(���Mӌ3���p�'��u5#sX�iu�R.0ӊ��DI���v=N��)���e��kZ��7շH�|o\���Bhr`�����P��Y���[��:8�����Ns�/Y/��:�� +��_N���p?-@��������+
p@�n�(�j�c�(wK:f��s谔�H��ipF���EW2��NB?�ů������6�~jP:�r#_MZZw&��ƾֵx}�ܽ^B\�b�խ���'�{�CF0��Oj�l�����9� ��[ ܑ/l���_�i�K��o���,��В����هD�>�[r��.>8A/���̷�e�>��H�M�L��ѓo\�9j�&�6t�go�#�O-l����G@��f��DQ�~b���0��;�>;z3��$& ���Q���6E�X�i)�(��z�� �����♵��sZa��g�c8[P`p�s2��gI�e�G�w�H��2M)�>���ou��S>�R�:�"�/�Bm����Ȃ��O#�n�Ye->�i|#��R��~w���:��I��j��HcOP;ϒEv%N��b��Z��KJ��	ۊ1��#X�����Q�$������6GŹYG���j�g �$�O��$D���M�&�����r��:��b:3�g��ʿ�!��0����9#V�����1�`&5QK�B(*n�%+W]�9y�r���a����&��Y�+A������L���)��4݊����Eb)��a����6j vy#^A�C��]�����8�~At��p��+^�G�j^�@BH^�fh��cY%�S4�V�(��F��v�kA��Q��BĔӨ�J�c�B`����+�2�4�XUuuo���j��i�Դ�i�4�:-@��������
�l_3='i?lH��'|��'ٓ�x�;�����;<��TY����.�s�'�s^�G��Ϻz�J^�'zͲjg��6�,��E�/�}�i})�#qʘ��F��_�FPl,S�H�"8�܈���e��D�R���"�"O�m��*�=�!��lK��H?q�<��e�h!㱃��|�M3-����q��O�$�S��\���� � �1��S~�Ԟ���e1�V��QG�!ѝ�1#G��Q"N2ݏ��a6I'����`�L��^���j䅵-�`;������#���b�9
�^l�N�H0;e��<XU�n�޽�0��@��"L ;V�m�O�\wJ�����>3q�$>(Iw�?O�����!
e���n��:�5��&�(��B>NӅ��4w�G��"�ޮ0�)��k���ou�]����_JO&=Q*�*�����e.��(C��3b5w�P�߲&��j�ok��S׀[�b�{�/�Y�4�gGp�z�bQ�fP��q+Ǧ���O�6s-{@X��E����e� �89��z��E�vc�bp���U������3]1��T��4AÁ�2dD)veP�ޖ=*Cf�v�L�A����c��,Zy�Kl��޸���"߯͜F��@�����\)i����Ro��
M2�}����,~�@�&�l0)�I�*.	�V{R���Ɇ�E�i�!Z����"G �m�8-9�E}c�w���U�%�f)?�Z����{]�9�����/�k=y18�A��Og���f�"y�M�w?8�cY9Y��TgC�d��U�=���|!":@T0��q`�0��l��4L=Z���E&�r�w.�dWb�|�!��)Et{K{>�e��-�?<��oA��~0����v��iv*e
N<t�(u�;���3��Ӥ��@2j��a�ɼ6�l?��^���6��f*IJ9^�wy܁(��xE�`E��i�����{���;���BՄւ�e��/c��uo��/%:(������/����*ӔP�[�Z���'π/��-cZ�*m&������p�gh�?[?�7��px� |4��󂖶V��%F���h�5-B>�g��F��)|��o�e���5)o�9�zH��Q���h���Զ4��Յ�dPew�w����	O��u�ͽ���.�3f�����f�:������4�o4
 C�R�r�{�m��9T_����~ڛ$�#�0+9E�mUȖh�@O,��0Ep�2H.��3e�:I+����vh���9��H��!�$�3��G���!�B#Z���	�cZ�KL�Ķ\�Y8 ex{��3�?VC`"�Z¢Ǚ��K�o3�X??��>�Ӫ���<�b�}߿+��e�ȏ2�/*�$���Wr��=�^p���w��J�-�]��L[�_)���p��ӭ8�RR�[-�jJN�Y����dvI3�?r�9ޔ����5��]�rd��:�D��pyz�ie���B��'��=с��5]'�����&�Z�go�Cm���ʨy�~�����M������`�!�*��zbBd��[��Cf'O�￭n�r���/:��M��������C��⽣^U�w�Q.M8-��xz�7�͵~�=�^MkF5)ktR����]@��W+�U����^O��Vgf����1���>��U�C��D*��r�;H	z����!҄����KAu�VV�
zl�S�Z��7��W�ט�DA����iEK��`K���Yp/]=�BB���|^�spB?�sQ]�hn��I�������{=-q���{&�����$��zk�(�����_��� �ɼ�*�(I�o/��
��յ�?|{�0TȎg���unRebFU��=]_�m�����e
5�����q~F���$���D��`w���g��@��*���M�0:֘�捋DG�q��Ĥ�Dch��9��wb�����]'��9>p:��9��0�;`� ��(ޣ	�S0"�z�	����N�t'a%���i)���S(�~㰘6�9-��O��&�h�����`i��ȏ���Xi��Z^����q9@���[d|{H�@f�9Lc�A#b�y��[ �F��_�7^�����Båcc5�Jtҥe�r�]N�`g��
 I�q~5�~��"DQ]���.�&��y�k�҅zp�a�o����L�/�a��'C��Qtq��-ɤ�;-N N�<^ w����̛�������%�����W�fU�D9H�p�Q�)ݼP*�4�3-�'0�0X��4�ٻ8�� ��lJ�!�f:��ї��Z����5oL0�n`K�PGT��%���&2�=�7���������}���}�~�Rр4?�JT	�*zP&�\�{p���j΁_h�1o-$��,c�3�e���� �duv4��-��fgц��IA����~�^����	��c���MYc[F���=�צ�X}�5vI���"4�Eg`��W��Ģ��F����X����v�0br���:��b@��ь]Ԥ���@�O�H�>-/3��9�z��p��⬹���-���WC�w�� �"f�̢r����z���<��q��P���
Ly귺L�|dO�������伜���TmL�/�i�Y�.�u�\B�_�nɪ�(C�����Obל���$w�EC�M�w,F�!�����Lg����=���>X^�+������y�xZnO�B�>;n�(|+,�-�ȓm���
윌*55�x��2�rt$�ǉ��ZDA7�Z�0�ݔϥVۤ�׶��q������>%��f��X�����ȗ�W������B+�-^�~��4����
Hb�S��P�K����E��q8$�^�.P���@
�Κ�8��;�і$�>�J��L�ү&γ'��,�S&U��hU�33S��:��dW�h��9���E�O36zˇ��H����ȋ��n�H�T	4��Ͷ�}�EdIz:�7��Vo���>��<-p* ��us�`�� no���� ����}�_�j�>SH+,���3@:�`�-:P �t$u͔D�?>m���c*q�)8-��NYf�����+6d�C�\��*�,�ro�/���Q��$U8$5���,�S�秀��i	����>ъ�r7�Ԙ��AE9!_��bW{��8),|f����r��I	nӄJl�Ψ�R�.	�)���G�Ѯ�n
�:bK�0�C}�]V����b�a��?��8���&��[�����z����"���%���ŝ����g��֥D��MBX�َX��e� ��Y�r��G5lk>�e�pq�Qg�>�	���\��?M���he$XrZ,�����$�P4��:�S��|+��S�O�m�g�+���|�'Ɯw$b��B�)����ݹ�qo���ߖ��b�*�)s�F�聆����5�Vou#�y|��l{��/4g>���0��i�q���-;:�����<���#ġ��U:#tk��$\�@�<�&Ck�\}���>�v3+���@��,��]f=X	_���Q���^��ߣlug��)�BP|�^0[�	԰���7A�]���[ׅc��e�Lo��9��Êkhqq�ŵ��,�o� �S
���y��uI��?%YJ$���:P����>�5E\ۅ�oKp���O�Ȳ�
���sI���##P�?���q��y.9��'�9"�̌�Mu�h���񏡁�tF�hZ	3�F E		%��C�T��M2^q�|�nۗFq�
C�%�F��؈2(+K>l)������p�䃪=�4d9��:y��M��;� ��#��$�="H ��3���{��R�I�7���2U :�g�'�s�[+S�<��!]�?�����8ňg�A���+ޘE���ѵ~�^YÞ,yPN�ec8�M�S@��S٧�80�ո�w�V.�D~9���@��4I����E�En��+�kJ�L���7~�BQ1�5~P�p� ݽ�CkU�z�������G�������a׺"@l��J,���W"�0�P���I�x�$��2���*�'�R�wd�c�[F�ڢ�l������t����A�R���X@9:�\o)��O�%hd�֨g�����}��Q�(�V��{¹xM����M��J�ba��<��o��cbw�-�Fhs"����p_p��F ca􁶿'��4)��Q�p?�r��D!U���D����xB�0-����_o��)}1� ��T!W.i��:����֜��	��ys�T�s0N ��2h��i����i��D�o%K�1�j���ĝ�1Hߚ0Ř�Wq��N~~bh�������=�-���
�U;L!�Qª�\��e��l*���� ����]���9�1@�·p��� }I�ztPs;��U��O�{���[Ǚ�{��󿣂��p%M �����BIX��M<K�i��ߐ5�-LF�u/^�,9H��о�(���Q��4+q;:�*�U�a�^A3�����}��%����|��f����Q�����ȸ+�(n:��~�r^klN֪@x�Q3Ft���Ͱ�)K��  ���0�8��").�M�Kc��@�2\t�2%�&��:ʀ�<�q��Eͻ��Gɹ
���	���8=�X-���?�V���}<��a#�� Z r[/�#�dl#1��������a�V:r�|%x?2� �8�n����`�������X�[:�|o�tܵ�B��j2���QO��Q�&e�5��8��^}�,�h1ذ�C(2�I�ޫ �5o ���:_��H���`�k��p}���pP����X(#9���E��L|ȼy��h�K뤠��6T�ɜ�y3�������"��2`(a&����.�����R��96W�_KwݙO'�O���{|���wV>E��d���}��������Ri�@F��J�1�Y#!I5
���R�� ���Ч������(W4�����Z:��� ��sx��p��OC] _���Vyf����'�3���� s&[�Ġ�U�P�:s_�W]�ST Z�g�C��{I'f�N���s��5�2���e�1r2W�p��1����X� ���$V:��wA���n�l�.�����͈ |���r����T�i� �l�� ������k)�T}#lZP��F��V*��i�u�3�S�2z��c�v`T�Su�ht��M?�R��Wl ,v��!r6��V�m�v�	Q���5���������OoT�D�o��w��kVKkK0��fd3��z���'�ג�:e^���^�,i
��/�XQ^����k�ѥ��/�]$ߋ�h)/>�h����$ˢAh��d��6(�,��ְ�g�f�/`��8��Fb��3�t����ɭ0v�hy���������,�F���<�u<�K;A�wqA�W��D5�����VuwO~ڪ�;iѼv�ۀ%d�4նY�	�	9ƴ7�ʔ��w`�vj��/z8H �\a��W�������VNރ&�������Y{�?�CJ�V�]���&:����4�n؜���G��W�O�
�ۮ�����|�¥Y{"�\�s�^p�����N�N��X��0�󑆯Κ#z%�}G��DZ[��g�DҖ��%�㞑J�\�EQ˵;N*ktj��N�=�r��0%ԕ�����p�A��$�sF/p���!,f� ��?$����)-iJ""{;�P��WrA��U�F&�\��h8�R[�?9[8U����cjK���hX	ďu@|/��Rڸ���DT��z�M��W��J�������rz9�����]��FÓf��C%~�	7.���fB�~�x<�O�{���7��xj��1=�^:�;�����II-�eĿ���m��X^Zb}���,�$�-���
oq!|�h%� c�l�W�p��5F<��q�8��r��+�V��X����Λ��>��P)�po���l<�T�|�UKܬ��q���Ӑ|�T�C߁�.{��r��ќ=I,k9Ј7\MYŦ�9��,��������E��C�T��Fܮx���<r�)��CY"r��s�Y�����x����S �;���U���2�&�wN�t�*S��1|pr70���й��?
�mX����á�7p߲x�aԚ2m�y��tFב�	�T�*۵ ~J����ߦ��Fi�z`��Qq+�|xo�FwOtM8���q��8���M��~��f{ʛ��k㫰����Y)��	��$^:))hǀfI�mN�%�d;�LБ�랊��E�c�<@ 7M6K�:�
*��X�"�t��=k�vY\�د��N]�)�{X�F���)Q��p#���sȪPh+DF����:ȼt�
U��bq/u�~�OrM�ߣ�7�V겴N���C���a_.��df�%��Yz��s�f�����o,��^m��W�MVW���������*R]6gц��N�7՘�W����/�`B]����6OH*0��~N����u��w�v��l�l?��Q��� �ҨdL�?�*,�3�2��nR|u�z��!�+�Kd��pUP��7|�w;��"�	�	^dӼ�����MZ�	�.�KJ��B]�-�����̼����Q��j���Z�=�mgW��!:��	������'��+5�{�VѪA����d� [&��&L�Q��휖I]����*�8+�z����᧔��4je�[����1X�tf�'�]�yҳ�	�Ӫ�N���S�W��8S��0܁O� B^�?>��ߟ�~Lc�m�����ځ ��-�g_ſ�k�C'M�=�=�I�~%<��D���q����1�q���$���f�͢6s�%��b�- g����Bà� %�JS�tVU��LmD,�E�.���瑓���#�kc"�=��wT�>���r^ / ��&�:>�7~:�����s�����*P�`2��7O<C�
g�_����Օ�W��a�O	�GG���H)�����>:���H����Ϙ�%z��n"��"���1\��� �'�<���b[ ���b�LX��<{�����r�g�t��R|���:<?�Kʓ������"{	� L�(�;�"��I�{Z�b� ,�����i"\Q���"|*�~�]�ֻ ��}u!x���ɏ�:7Ww(����*�sM ��n1$�m�i�.��0W���(R슥�Vp*\:���_p���u^�5�Y��[|?�m�Qj.f��0pK�2ڬ���'�d���u����z���!�o��8��u��f���N$I�>��<�2�'�X�M������QTr!��ڸE��@�?�0�4*P➛�Ȧ�H���!��r�{�,{j%u*_�K��[r����S�cm���Tz�zOx�#���U'��Ú��KFd""�|����KԷ�ڵҐ3x�ޞY������AS]-D�eb�+�ѸT`��E0쀓�jd�%�/�m��Ӌ���֟)p�@����n��	�޶3�;�:�fu�4��
e�����_��v�vkx�p4�>��x{}1�5��~�%)