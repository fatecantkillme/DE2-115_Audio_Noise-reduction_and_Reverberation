��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
|)t�]з;�Y7�^7/\�ǘ������W��O[b�^��nJ������`Zu�i�[��Eu%F>�,��ry��� �]�U� D!� `{�RK�ф�9&��nZF���(s�w��x��ѯ#�V�D�D������]ӵg�d��j�\ �X���SBN�?�&��~�o=i���	��n�����«��>Y�7�]Y���ǾW�S�H�������'qs�+{m��-��7PE�=���D��3Y��po!呻�-�T�\"�����K6���OMŦ��G�$��_C�p��%) I6� +k���k$�ϫ�ס�κI�~'5*�/�'���Qǘ���6������|@��[R����.;e$N�VݩtV{-֎�E۸�7����T�2[�-�7qN~S/Ѵ{����=��=���ђ��;k����$ڦa��D�Z�,�����4D�+Wv�4-,>PhR��������P=���$�#O�� ����&��mTm5/���稰>di��[b�������.c@_p��x�`	���d�;�uP��e�J�1dgĐ0�_��+K������.b���w�o[��<�v5_�*�!�mA%�2�F�~	B���a�a.y�*�c���ܡ�m0Zs���8��k�h]6s^�Kk��;�� ���y�!{?�ﳡ���xk�8���k4<��owdo�w�����%�!��afc��f�H�oP�X���p@j�,y������T���*0�"��8�8��2E�ۆt^����oj����y<���/
�ym?V`E���eq�L��m�b���/��q=z��jO{���t�sG)�A�a�)3Aeu�u�pq~s�8�=�T,ך� ِ��Y��(4�?9�pouv����{�Kv�?�<��72禲����y�� ��ZI?[r5���"o���1d�h�<�R_��	s-���Я�����N�E\[z�hwW�*���3�qx��J@��*	��% ��7Ը�����KA�a��Ր�u���G�π6~Ng������_i��%���S�]dHw0�$|�XP�j�&$�"Qe����� +}5�!M
������?Ħ��t�q�Yx=�9վ}477Jި����"�����х����^���.mQ�?��R}��?#�����xv�Yťl��V�g��]_*��\�Wj7��m̔?�����{��k~��j0��޵ ���#N���ǒXLI�l��_��d�z����yٺ:��U��i���L;pvSo\R2!nE�=��,�SJS�JtR�>YɾE��*�����6+/8�+\))޸���:�������7T-��-�t�R(�p,G��
E����2�{�����ocJ9���=w��|��*�$)�As��4�f��+e�U�hG�\��thN�qb"8�ktrdժ���YnNx᪱�1\�r������%��c1±�h��X�R[�]�m��wy�!����������_�Mз��.����߂,.���;���e�)�>%:gϟ��Q���nz�GH~�(� .�˘�Q�ʙ�mg� aάH+\�cV�L˚_%��(�?e��=5����vgc���+��h-�cN���	8f��r��U��"����n���fZ�>�C����'��J���TxZF'I�4��YlkP���2�g��C�,6 g�6�|���O��X�ޗY4	�A�':��/���X'/�������VL!g������'���n�5ɛ>�w��g�b��'ף���TA��e6�P.O��%�U�ho����6�}kצ�Qo�w��;W��Lk�R�(�䛾k�u�l�����1\"	;��/m�e���Y�1���>D�����֒>p���X�	���vٓ� H�MdV�+���m��B�׸�;i�Dd<!��h
�l�aM�&�jD��F4�/�~�h����R�\(���[�H�#4�R�&t�5赧�ˮPf�H�.�G��ޘ(@�_ �����<~G	�H�Fe�V�`�}���PW�r���$�������&xC`��aGF���N0Lt�v�56Q�<qY��op�E�T���*I��*�Z
��ZEs�gIy�IM�����ۅ��]�I�38����1���I�V�.��4�'�kc#K|�ks�ߜmx��>��R�w�]3��@S�b5���گ�*�L�u	��}�~IW"M���3��2�=`Yx:�pcB���n�DV�B*�P��ELp�j�N�D�XT[_�&�6�D��FXfld}�bn`F`�.9�������_�ћ��Q�X��(���_lA�D=q�p�5e0�z�"��
X�mt#(bL&i#g�T����:��$XPl�����ԪT,����ڄ��O/��p�\>w��$�Q�U���|#H�䍋�A��̹�����G.nOL0�ݨ5G���
��Z����unYc�%;�7X��cDS3p����(c�me���b���4�o�y�鷦���)q|��tڟ��A�G�+��!�h�fs^g\?L��5
��W�iݍ���:����Ϳ�cPJ�+$mM�8����ֆ��~�X"��jlA�|�e��V�v�ɵI�[����ա+W�X�[�2����zy�'-�DT��}�(��`o�|i�/�:;���J���>R�A�?F%6�x�m��S��C�T7��}xtS<�4C�g�Z�>� =�W%`?��-�5��XQsޑ��1:�I�Ԕ ���QW��{ũ���R�,D,�����yR`!��fteNx �N�]]g~8s���|��_��z	`��Ι��m���:?wη����E�ID����m �Y�'��WX+����?��yƑ��r���I�]���z��ۦ�toδPB���^' 0��G
�,^��,�F*r6$ي�V��!t~AVt\�7��֦Z^�WL}�BOYë�����	�h����]�6v@�'m� ��:�4;�g3v`����:!� �pJ(뽐irYv�V�S ��?g�]����V�e1i�>���&��C<��d�9bn���G��S\ݼ�[�4�z9N�$~��8ō�6�2@MQ&���I>w�Q��h�K1x�w� y?�
{�a�V�U�KU�oս�6��uM℉�v�9��pI�����C@�L��:���������u��]v���KB	���L+�+㟕�t�;3GGѾF��ek$C�p����=�!���F%ʦ�rVs���F�<#��QP�D�0���w�܅��*k�b���X�����bqgH�󹣼�Z�R�J~��v�X�����������aUg����|�5��r:L�[+45�o5���,��Ov�hJ�"8��ޮ��&8+�i�L_�+���=�>ɇR��=�d�^zUQ�?W7t2��R;G�t�Z!�z�K�ߺ���'~�-^)%��}21j�����\��(��?)��V�m}ybgڻچ�u
~] � �O��aI��؂��]������˾M���6�)T�'�����,X�5po��Z-�����X(���7����o`$~�ݻ�3oG����BM� ���� �sa��H���q��I�$�0����V´Pϑ�{��i7��,�"~�]Sw�T���;l(B��\Ӏ�{ҚlP����ŀ����w+&�\��� R��يKS�9*q��V�D�}8)��0�?/v��dRru{���g0a.���y��ëL��l�dC���G��c�gЀ#ǘ_D����Oh���6�Vu�*�Ns�ї
ݏ��o<Z�t4sI����E�%�}���(%9ŉ��T��X�(�H��킮�n⠳��-j�нa)�0ke� &:����A[�rn8�zj{���	�u��Z��]��tF��1E���(y`���8`,Ye��G� �����K]�Ƃ����u-���,H�T���f$i8��.g�od�C�{���3f˼��E�!kD�.˛n?4أ>���ۋOV�w��3*h�?ov)�1���B?&�\X� ���_s<�U�S�����&�{b|�Z��g�
A�K�@�Y�LB/Hϯ����/:�|���[���S'�tW�Zق�*�B�gC^�Tm�/K�5_1�K{�)�q��ar\l-Z,�"	��?��hC�?z��������l�>����3�ЇB�퇑+�g:]MCP��ڟ�
I��\v*��?��	��[�<��w�VE��AU%М�S���[E�$B�x�^^jv������$���!�k"����a������ڙvG��G�*|�7B�xR��⍖����a�
-~�D��쇈��f���uz9pS����c��ˋ}4�̂y����թ\�#M��X�`c�ٶ��d��	Z��5۸����ꏠk\6�6�B��q�!�"@�Y����
���p�A��E�΂{�=3*f�8S,�>m��5N��:9�Mg��1��t1��y�K�p�s��W���E՝G	����������හM$��f��o��2=(a�MdHL�.
��ƯR;�MT��[iPuy�!�r�Q(��5�g��GM���
`$� �J�<�����ۛR�{��~l�˘��
���.N\%�Ia^��@�S�W[�؃�L���>���<c2$�3���Y"��<�)nܰ�;XS�e��ȼ�[��@G�D���[��_mc��!>nyS	���F� ƞ�2^��V����#<��Wt,M�w�G&\�@!�h:�3~�"ާ�o�,�*��!W�S����%6Ic<qw���根�d�΂ߧ;_�c�"��H����o�p����PT�EBR�+�Ɨ�'��H��A���p	�|  `�q�i�{�T�^�F85�����u\S��i��mf���!S��Dg)v����P-sth����K��2���)�B�gQ"��2�&OWl]a����ٍ�`|,�x�0���3)  ���,X�>x��V �Ij��Ӷ�t`)):�C��u�F�s�B�F�<�Sv�(��$*r4���˅������?l�(y!9�#uШe��ms��LYZW`��qm\r�KYWG��]��*u�;_Z����$�2��-x��`ds�3� �Z:�um��+栱���]qH��F���~A������LA�W���+�U�C�,����m�t:$�S.G�l4�5:�"���՛6STC�1CWU2w�������ʛ?�9�{��5�b[*�*)�w�N'D�;vq�QR!d���-�Ӣ�zcM�%�LJ������ƨi~@(|z�-�ς�c���.��(T���H�,�<W���׬l�u����s�cH���A���05��E�(�9f*���ؖE�����P�M����`��X?s̞Qw��#NBC�`�t
�C�cTU�& jY�Wm��r1;
#^���N�[�긞�QdK�� �a�'�Ǟ���ܭ}*��	Mo�M�HkMzV���ԙ�^��2P.�/�,U7��Ʈ�Q������ �,Cn�
���R��~�:B!�T>�B)f�5n�(v� �_n��J���S���%�L�0�;�&L��9�U�b���M��xP��L\�����Y��:��b�����u����<���(���͐��ҏUf��g���t��� ^�ʈ����65�ߚOi��J8l-l|�e#���Ҟ����]C��dpK��*��Dy%�����*[z�4q^�I�������4��&O�m��iO��C{{��v�n�|b\͡�wB�!����J�'q�"�oZ�����۽����x��j�#ll$U��F��c>f:�b3WK��IJsv�nY��qğ�
U�x�_����8��AeZ�m�n)�J�0}`�m�����}�Z��ɢL��?����x�.�؞<=b�gl��-�V'�~�p1B�D�65�I�2іj�H��=ʜƾ!I�!�-�Eya���\�/�1m�&��{��B�)BX7��(Q#�px�Q$#g�K]��Dĸ��_� �hlg��6`�I慦�?Hi+��)�������_������gd~Y��|�nA� �3<E�Z�x$>�o�'5#��P!u�|vO�c�����GC}��_C�t1���6�x)S��e%,��g^Ѯ����M\�b��s�]��iڢ�^kR���b\ �17��@/�`:
:;�~S����t�e�vͰ�w׸�w>jPo�s���RaK�@���C�h�U�W��c%�I&�6�s�_im�>�,J��ީv�����B���FųP������b0P�Q݄����w7 ۧ�7��
�� Փ�7��ê��H�OE�j�P��-�d-�v�nHk���S��!��i0�(U�y�g 6�D�t=���N�;Ǹ��w5�l�;?�z�����qnzx�X���ϰ��>2�S���R�]�]�j�rB���5��Xo�^h���5�d�X��U��XU��0�ӻ��og�<͓�w��ݻ��)�jgg�q*�/�fl��z�����;�u⁘g?��4!�w4��g	����0<coN�4���j��F��.`S9�'�������~{Eܺ�Oh�z�!g��Np{ǶثzԠ@�pR��e1İAy�%ٸ+^��{CO*i��h�2A���So�]D��/t��&;��.`&�W�֑S'
?+��Bס
3�p^���i`�fS΄�h���T��sE��ʅW��[*%L��_��V���_�(���6X��$���	u��_�D�U>��Z�Z!����+�ۀ5
�}/C��;pA_ۤ6���5N����+S�1?$�W�����O�yC��]3x��@G8v���щ��{>�P�����N�L�}�g�\�����ꮸoOevZ2���a��U _e�����a0�t�/8^�Y�U����>|��#�Hq�N�ϼ�����4�r]dW+�'�-G�-�L?�xa��r3c8.����#Fɰ	)
:x
N�N3�Z���_�$�L��;M� �6�����7��U-�M��&�4��i~ş4tB���٪D.�����7DG���1M��F,a7���.�3Ք�p.����R�;���(�D��H��Xvπ�"p�>T;_�D��N��?��J1_���U�_�j_x�rDA�p���2�"���Į/(G��N��XXH��y��RCka�E)�x���Me?�ц*�x�(Ei|^��7#sq�����������{�	�J�2r..?�y۵u����}�Qmo����[�v;��Y� aT Y�$�r�̎���G'�'����``��H�]t���,2�!�w�7M��\F�ɱJ&�,k�Y���+�z.������A��n��d�	��J?��.(�.|�KZ�������,�E耧�+���Pn��jh�
�PY�?ri�3�,�����-�u�fД�wR����s
9u��Ꜩ� �h�j�G�P�@�ln��a^�^�c�@�+q���'	7����U�h��C4�<�1�>?�����Z��7��蒍��b����RP}�����8l��</����Ķ�G�و�#\wVt��Շ�e3aX����r�Y���R"o%`%�G���������LƁq�Vr*2Y��Ȓ�\�!)�!�ת�b�~�HY�[D^��t�I��<e]��F�6������N��͡��2Z���-0�����z�e=B�_�E�@������&vN������h��[�L�Ԁ�����~"����w�ɵ3N�(�=y���]�(��%q�����D�Iؗf�̦%�/h#�9 ���vR�D����G:=���3:��8�~�rZzP�ϐ���_=���t���AvN�Z�1�:Z��	B�������c��нI�SՒ:jߦ���6�ח�T��d����sA��b�\1#I:=���H戈Q��@�	_��"�a����]��f#�t��8JU�ւ���-��w����n�4�-�����L��@�H�յN�Ւ��$���i�:�u+"-L��	�� �K��.2���a�cê�*�kﴛ�a�L�;Ǝ0%@�����zOz+�ۺ|�Pdp�X].u3G�x��9|�&�9�u�n��V(I���1^W�C糂�1��\��t�6e ��҆�ӝ�at�HV|��F�_	 Sux.��qfw\/F�(���[|��R/���Ě�[��o��Z��ܵZ��Ў���X���a�'�m;j����2I*�놫v����I�bD����<1�6����B��[c�D��[���ďw#Β\������ �	�a�XWB��fw1��M����<����s�O"]��D���eL� 	I�p�o�FH�5$��.p���I䚻�m�Dj�(ɅH.�v��y�Fa��>�$$-�֫�L����>������Q<������s����W��9m�M�D�g|&�! S����z�K�*3�z�i��rn�}��$���#2F^��?�{}���S	������ouf��<�.��#ByV3�+�]y�c|�Z�fa���5y\����#����HT��l/ sq�#o�@�e��#ϭG����l��b3���怨�ZY�ݗ�/�e�ϴ2$�[�u�a��Ti4�����s
�J�F��%[���Sp�A�����/��Te(@�u�� �ǜCM���C�?����2l�6ŭ4QY0ҭdI�薹��uv�P9n��uyͱ5Z嵸|!�=>�*�n�?�NG4�.t����Ϋ�Z��Q֕
��%➿���z�I����.9y}�Bt��9 �Ȟ��n���-�D�\�%�c����Hr���r٫�D1�8J	�@�b�"�*�%�$��@���,��n2�b�Q[J/�\���B"r3��7�b�0�	�b�7M�W ��ق��\^�8�(�B��L��V�H����mЀ�{:���z��5X�S��$��C,!���)7ĕ���[7���.�Z�hb���K��I(�q	p&J��QH��N���ʳ��m�ie���=�ß�H�Ҿ(_����v'��	1pi�1��$��\�e_� XS����_̬����ϑ?���Y�&�^�ǐJ��q,�'@D7�Y���X`D?b�]�P����m	9*���i�C�ɍ��$�u_`'b���>�J�-��Bx�=�6�<��ޓ��S�/�Q�!k�]d��&�:oZ��hH#��������.qÌ�㢥�6'L����c�7cK��"#�=a��3M�� H+���(,4��Ο�v:��f�%��Dp�A��in7���܌ۡ_�Y��f�^h�Ȏm��\�Z�;�칛��B��8!}ǽ9E*�A���YY2�f��IJ@+��>Jp��((�)�H?P�l�a�c��w܊(�7�NIR�r&��0��ZbáZ��[.&�b	bb�O�3�*���������S�I;�}��*�Op��%�̾����������ű����4��u#��4�k�:��/��� =���kR�z8��+�
�#����*�^�[��0b��7W�����ih�k�\�Z��s�Ю{}�!�/���J(=��TA��U���j��Z^��Z��d�	��������v��Y�C0�t��]��gRq�aN�^�I�Jny?�t*F��z-=�+��ؤ���{�{�ևW�ә@���A�ݞ�~���oo̯0�����v���o�}.�n���~3�~�qb,�,�����!Z�iU�Rh`��>���MO�C�q���Y������������o�(�:,�M�e�#E
O�:��X/ ׬#�����l������cp��?q2�w�����e�`f����P���	�R�z��j @V��k"%c�����g�+k`�8]��X�Sme����h"���l_�h0Q�SV0!~�۸�QL������e2���Ki2�q��a���1���j��HFdKvK`_��("׋���r>"y\��,�a�3rд�̄��L��9��j"/n���>�b��Q6��v����Ss�ET�j�}��n5�0�ʆ�oV��e�� ��)l�H�
l������ݥ8��Jn���]W���'��T�0"L�r2cM,w��"�Gs��r��]NC����浍}��'M�A�o��.�ܣFA�!	�m�9}����<������fӐ��`-{J��Ge)�8��G�Gqzw��rZ�������J�ux�}b�c�=gH@�u�_33L'N�����Ҩ�����ģ�|I����śͯ�U�ͮ��2w��>��;�ս,X�ac�w�왨fF/D�hm��]U��>�l]ձn9$��,#��AN
!��f�[t�X��Y0$1?_sCھR�A�9�hU--rn�.=Q$#/
�Q)G5Z�a�a�33j�P�L5L�NS��%��]	d0I#��"n����� o"a��B��M��Ύ3��g��F���՚���.� �����O��̪H�0�*8�FX>A���>����ougFD�UFL�5�#���-�.C�o4F���~�U� 0�A�@H|�Xt�Z-o�K�����=���fH�Q��w�B �x�d�:��K��,�B�e��9��(6Q����g鼿��!�y&:/.ih��$gJ���@���Ġ
-��IϚF��аb��*xm?L1tU�~�݂��$�]��)¡�i�$��(SKKDZT]㴳��^�S�������D�'�d�{�sL�̓q�ix��	o./3%Ald����-�<��y3dȢ0pC������J����V��f8ix���Z��z�I7�\�yUQ��O�ȃ$h(��DX�hd�E��x��^�{G�˓ d�ő�L�4	�V\�#�;����ٹ���R�ӷX&.�
�ؤ_鍪Ζ�M�L��g�>J��G}"�[��cIas���,'�1���k�7>���Ц/��I��P��-��-���׊`z���q�`�Euj3������o�|w%�����FU�gBZ��-d�{�hc�J���4�/xZ�b9��ۻ:�?՗��������Ѥ�G��ᗐ�w��B��rj�^�m����Nz�{Cp\B���ՠc���g^4OD�W�t)1.*���ƀ��N��h=wQ%*an����kP�&JA���U�J��k ����[L�i >O�g�DK���A�d��6@��5���(�1A��R�j -s�$_��W��ȳ���3�����qi#�_��t��cf���#��p�G<���qEVe��pT}�2���ְ�^s��)M`����3_.m�$�9`���ԝ|pT���{\[ty2lsd4��<U����1\6_�C�PP��.1r���*�&��
�KZ��d���փ`7�����Cp���J6���hD�jgI���l�Sb�)�ޛϩ+9ڠoP�Fa�?l���؃n���"��.��8�����9��VvL��f2|���܁(6�޸\�Cw	w ,qy]�Z�WQD���J���®�sO<�
ݳ�ǯ��������ƕ�k�_Z�L��,J<qH�A�ec$˿�G&xe��%ۜ�=����"����l�c��b�����2��4���:?[]j�}�݈C�v���V�Cq_j�F�0��^�Ȇy�Ǆ� I!�Я�L�Ӧ�PjÙ(����D_`��M"�����+0*�7"fEÉ߁5�Y�N�.��|�b�����S7��/�_����C��T�U#T
����!���d��ng+�����ov0ڎf���iW��hu����I�6z�wk��oru�(j5�Ջ���܁�`X�����Ü(�P?�/��Au_���Cay{);sjc02��/��U��WԿ�ߢ���2Шerમ��=�d�zh�O��&��֎#�.47:~!�擈�,��K<x4�	�� ���XvM��E"��ZV��έ�*z�j�؃��h�"}CL���D������Il;W�J�|F���|9�i?���߸S�t�d)+��r,6:=<\+CGʨ4���~/B�Y���s��(V�2�$�Q��qY�����R7�ӫ΀fen����[�gs��2�@i=��X���U>��S�`"����,��|��u:�"ܭ�c����?A��T�+quo�Y4�)�j���sQ����R��J0�j)��0��f����4~�o�
�vyl7{H�1�4���E�%u��RN|���@@xDr,� &3�r�,�'��
Os��^M��,�Xܨ*B�%�G.X����;T�ϊّ�
 eS��l
B	�8�5��&�1�s�9�����D�ED���n#pkѯ��^'q�2e�5��s~5ʟ+L�,���0t���F�.��˕������)��ZD��Y>(���!#�.?B��濦�K���FJ$j
d�UN�������(W��r�ts��&3?���Z.v�.���M�B�YR��N�<�0C�~�f�w�\.cC�zM��9}`�y{X��n"��&�f� P� V	IW��x_��,���l����лP�f�m�Np5�}X2.�SS�k_<GC;��ߗ��(ӎ���&��{-��+�Q_�}�}�@Bu��Clh�L5�1W��وɁ�S��Q���\Ĝ2�~y?1
�� zr��#k������jV��e	3
��d�Սrs��N��"f�d�ü�#?{Gfʪߴ��(&��zn���y��$�L'������J�����jh�0�
�S��̕�ìȴ�+W�~1��b��2Q^5������9n"E��)b��2����jb�|^��=DP�emF��3�݇�z}� 	� �������q��q�0Q��8+�r����53{�gMa��~-"?z(Lbj�����-��K��wdQuO0ǽ�$�5���>�p�%j�6��3�ћ�fj������h���J<�#����T�y�6b��Z��e���ͷ��l�o��/�/��!�ȼ�ɧ)Y���W0����u`��y����[`��PH��� ��%��I��,+ tܨ��R�*��O��Cp߈j��_z��^K�,�L��\R�	ƛ� �tN�[hZ{��%r2J}�Ւ���lug�6�/m��T��~�٫�/%_��j���˹Տ��S���%�ic!۫D�Iz+a
^�(w��#�!�q�څS��)�*F2�PT��)	^�s7���k�}MU]$�q�.�l���x"�↬6���!��K�D�d;(B8�D�zX)��o��#x~D�q#M���f��^���r5N�b�4]w�$�-�ߗ�虯�x6��G��=\,��"�vPh#`�k�[-K�ә���L�[H�(,ad�~��8\]�&�ˎ2ٲ
��ì1���y!�j��ܭ��]�52�Z����I���ELN�$F$�^��p̖u߃�/vx}�>��ݏ5L"hs �&�9��ɓi�ꈾӚ�k@:�lu��z�cy��Y����O=��#ii�˝�o�6��q�G8�bH�r$���g�$Ƅ��m�0A�!/����_�P�ZYR�m2��@s ~b搙���t�ăK��>�1���7\����ie��#n��l��>}e[tw��bQB�E���zր� 	�V3c��fz�Y����K��y(�+Ş����<<�V	�:�o�_B>��D����Z"��&��s6}�+l����6V����z�pgHA���u~AѨ�=���g ��{�p�w`���7y9{�j�Y4SG�O#Ğ�b^�]�VW�u���,si�(�j�)|�	��1�S�����E�9�f
6�}��g?i�6��ۏR����P�1�,�j�7*I|v��������,�WY,v�~�����e�~An���ݔ��*�;�bS@�1���5�-��#��6O���,�I[T���@��(@�������p='���V�};n����m�����A��d_����iBFk�/U8�-'^}�W �b)Z���)�[���7s�x�vQ ԿN��C���iRg}
������������@�ݾhM��q���1i�sl�v���6����EtZ�N��߉̰#�(d�{]���7@X�u�LT	a:�g��cس�P�<vٓ�����"Ȧ���m����:�G��|n�
�S	�V��V�ϖ�3��3#�
�i�٩�)0X�~N��Bo��]���#�3��c��j���ͫ�Hƪ&��}m� 9�>�o,#aF?BW=�!�`��^ERG����5{Қ>���<9�e��X!�G�RE��ї������:79�Q�r���^�eM�Ǟ�0� ��n���<���K� lm��;$�%�z�2���<u>j�A�C3�QT�/+v�]��bh��z�`���&�M�=��}wK����d�J�$���e�
�{�_L6�ƻ�7��$���r\��� єz��=�D���]Z�d�_�dǛ�\�9 �
�=�<�>'ܴ�H ��x���1b��$�j'��߮�����ߑ�%E�:�Hi�	�>"�
֣�I�x&	�(�򤿪d�/E8����#�l���ӺЛ�7��2ŌY��l ��������(w�~���%��p�ҹc�$��c��z%�c9N�R��v<umb���*�M�eܖli���ݖ�4�b��4�0E�#����F?���$���@x�(�5$/�ɶ,b�gފ��%�[��O�
���c�:L�A�	�.�K��0N`̴���,�ٝ�p�ew����V���)V��P�����N>��6� UK&��`�퍋=,����
��7���th�~w����I�m���б��k~J������x�q62"�06�r��omm��d��׆|���`g����񡻮�8���^�vO]��ڷ<��Zd�VR�4��#b��aXb$A�F���W^@�a3C���¶v-�a�l�u�h�_k���7�s\���gm�]�dA��`��3iS��б#�r�:x�Ak�o4�˷�������m��a�-mS�I>���JZ��.ߑ_���E�x%ڷ:6����עy�kH �+�eX��_���zU��p�D�ۇ?L��	�{m�5+ؚ|�-�q]7�����7��J	jLza��Yo�pj��VY��"�vJ.F/isH2{�Cߥ��]/��7%��-��`�Rs2j�/C���e�g�G`�չ�F)�+�0릒<í���ݓj;�U2�⃠�]7����|U�$s������(�2�M��t}���0q�x���Uث�;C}�E��oE��}}E��+�9��:]����Q>J]k�uֿKd�Z�7��ZZ��v��A�����������T�1D@B,q�ZK��~/�F��!�M�cU^;3﬍Q:��&���R�9-a�(v����|��
h�����p��k�ϓ�%Q�]��u��([�+���� ݂0��)`�K�8�^{��#ϵԞ��
3n���e�� K�&�xU,��[�:�}���J}( �6�}�'��֊�?h5<��R����N�"��rP3}�%�# �Pae9���8��͚vq.V^��a��8��Td�MU�s�Y	H5y�o/�OՔ��$�*\�d��W��5\�V\�Ύ7���bL�2�?�_~����;���UN!�w�9����qg�I�3G��G<�����(߻�\mlV�����"�X\��Y�ᔱ����y�y���lʹ����rM��� ;71��['���!�xH�k�a��k����!48(�e�-�6 �bHj��qP��&d.�f\=a���4WU�ę�%)3t�垩J'���� (l���Fg���m`,F���E�R��B+*b�L�(�����܂CE�8�T	qsw:G^���f��Yt���O,�4s�}eQxje�8��#�q5��ң�t	���1�*���y��>�\���	c҃ ���d.�Bߓ�R��I3}�q�g/q�n��U�,k	�bev��-�{�<�����*̈́���~�?�ɏ������B2������ �},���q<���h1��E�m�X�~#�d��	4|k`m6l�-w+�]G��Si�E�c�RM�کF��=-�\OYI��^�8�۶4 xG����-�%&J�g�6׋B����������"}�x��`Z�Kx�B�D�y\�� 2��u8��V�8�I~�m�5Ubћ���A��^����)�*{K�;J\�b������y4������'��j�
`��v�x�ٔ~�փ�Z��Z	����{z]@Y��]��W��]�g0�ST)b�ϴ}t_)Na�0^+ų7"�ey %>W��Â9^"�K ��x�`J4��{u���R�����d��F$<̤�7���;5�⨣8��XJT5�!R}�>8|�'*g�kF�̘M�i;g�"8�T;�6�ME�KL������%>a���up�⦯�T}�C+l���{
�ƝmW$�����iP3 ��d����ׄ�-[��+ѬLډ.9�c�����IA4mX�r)J�Э��˔8��d�q���uX	_Y)�տ9����� ����(1��I'z�|0:�� �?�=Ť��r���j��1PX��0�Es��
�n�x(x^��ک�l�aS �,�ga�8�餷�̡����iAz'ʊ�Z���?�|u�eF�.�=�W��*��l�_7`�<��Ä����(�o��#�e��K]�\U*��C1��L��}���f&��J��
�i���M�o��t\��J�t�^�r�-��rVؾ�
(i�L)ǎG���+��V@���O'�dc��?v��Unr�O]�[��%7��u.���:6�2(X�׼�CZM��8���"��^	 �m5���s�����u�L�f��
���n����i�v��҈:�q�L����!9�w�6�kpA�W�v�a7Z�8�F�x7~���dm���LvP��{��0��H��8}��O�6����%y�9ȂJ�Yr�����Fi�h>�=��ѥ"����-:h��^kr'��k�t~/7(44��,]2YY7;�G��Zt�� �eb��R����c�f:^Qee�������;Ju��a�;2�^z����]� �j�h��Q%��v�#���y�P��8]��r�(�����<��m�I1�盁'����Z�����J)U_��_Fl)�w9�خfRp��F9�B�1܀d/�A�����A:��$x�_x���S����@u�Q �(kͤKt�IW�����%�&
pc��!��o��6�џc���Pn5BIےD�?�(U��K�qX;���Gx�%o�)3u2��K;fQa�.��]��Ξ�������J�L? �c���z��x֢al�l�'45�:4��� ����g�����ܮ%���f��Й�J�����p2{�@�I3��nC|έZ?�5�}���Ao����������<�JwXI����pw��k%��$e�B�{�	��w�'��e�s�m�ՍV��x$�"WR��6M !P�Q����5��^�Uwm��^/��ױ� �DӇ�ܣ�J���`��pwH�Ѥ�^�'���Q�������6B/L�<��++�Ϻ6��%o	���:�i
�&lQ�`�؅��e�Ը�k�2�n�Z{P�x����7Gh^�������1���X��{� ``LaM梱�t�]�� ����AГ
9�v�Ե�R'��h_X(v�C��%{'��ߗ�`�z��_Ek��=.�y{��&%�@m��\���2����F2�wD��G�f~��G�s�}<�)�cG��<�8�j�V$3	��7�O��t}=����Cb���G=��ǹ9�R,����v Ơ����i��H�Tn��7�s�>�Z���DF��z�mf����m��C���.�H߀`b*�TH/��|�B�e�|�sm��O=I�L1�O!��(��>�~�J�q᪮/��]z@� ��Cx����ʗ#��C��s�kF������hU;��h�l�7�RwR��C��g�,����GFl�����'cx�`�R���J��!�m
�q������񚲆k5��&�U���r�B�F�]QU�[�#Am�M��Rmǎs(<�� W���4�ezј�R��%i�6=���y5�x:���*�_��<�0իY���<�6�s����n_\;Wڹ	'�c�Nٗҳ���ӡ�w3�r���{(�M�t-���e�I��D�jw[,���{�=%��;{"���v�G7��J��z7������xb���HưTH)�>�ݵ�M1C�}�U��Αe�݆�1�J˃]�j�Dj��؝����FGO�&�:Ǉ7�L��Q�ٮ�j�@/=ˤXS�����g3�F�������s�2�v��y� �_�O-5N$}�Sϫ�ntE/!Ux��^e�atדY�H�؛��2⌥�[0�a�E���x�.��ɦ��ԁ4�*Mnw%}p擊ل��&;���D�r�pR���/�����TI��MCYDG9���#����,�LL���',�\��v��d�9�������P��)�X#�����E|��!7�ë�$��3���e~z����b:�U9|�0�s�D������0�_4+�0��.l��E^^�Pp*�}uCȚ'�r�S���c򄲾k+�W��X��D�3$�|.�/�J��,·�B��Ǜ��h,ᴧ,��Y�f邩 2�`�t�`kC�?�y]bp��(�O�\�I�ԏ꣭��������&�b�'�R��)�XNN"��v�'�gs���*��-���1e���%�(\̐�K.�	�8ټ�`�NS��Ԅ٫R���Ǆ[�X}~��G.�Ǵ/�,�m`~�"-��ǉ�S��z�.r�9k��Y�
Ԟ�gS�I\RV.���K: �re�I��������'�+��+��H=Ra^e\[P�*�U��}@��������F�ca�����j�ۧ��脣��MӘ��91�0�3��zOT��c�i�:-��P�;s'��dX��2�.{_�=��5�6�1�=�3�Yfο��t�oL4����T����L���L���;ak��B���|�xg��/KW��b��c����:b�5�ή6�1�,�[hhz���f���x�+�g��A��
��}��	J0TG�/� �0���	o��c�H�H���Bm�W-a�����,��q��h�g�g:^��<��u˺w�Ց_�J���4�@��[�*�q4��F�%�opQ~�����OrR\i��ޜ�DFh"��!8R�Ք៉�N��"�>#��&O��%���D���|\�c��W$�=s	�Mr�Ma��X��9�v�FA]]�]�5�ruj���u|$������
Mg�7";�_���}�xS��S�n���5��N����t���d�p�tn3c�R�4�4�fxC�L�*}f���8�o�}��- ���مbBf��2?�U99Y��O1�0!Б��\r}j�ǯi�I��ȏ*ݫ^�@m�!�����H.4�������m�1�+2��c"���X�V*,�$�>O sq�R��C�6y
Wkp7�9c�D��d�V�D�<t>z� �5@l�r�z������%��\g�)��%�y7�w��׀�5k��.���8�
/��WO�aD_-�JC�-��3�#O��pIapr�v��`F'�꣉��9�\X�ΝoC�6)М�ݘii�(u�s�lf[�d�M�)x��;:�N�R�ޑ�~��:g|Eyx"����&�`X��t��'�f���R<���	��<b�@ǆ3C��=��hї���<�N����j�P�;��T���)!LV�L�[�уk�H�u�~uQ������S|���"�\'U5��{�ϥ�v��ܩ�#�w��Ĝ�8ЊR�*��X�:.�19P�s�u���#i�i��Z�����&�Ae)�C5�AiI���6\+['&�5�=EE�-�,�DI<G�Qא��H_x�ۢ��5p�I��c�jG軔/鍑*>�3G�)V�G��6gJ�XG$�w���jƝZ�������4�0G*+ WW}3����a�m쪕5(^�����/�u{-�y�?�B$s�}
�㌣ʬ$_ѩ�<���/`�?��G�KV����`g�nj��@����06#j��� �`NC����0��)��tȆO�����}�� �c�<�m��mX.{���P��E�!P~Y�UE�Df�t�#;÷a�y��8�'�)�\�WU�F������eg��"R��wV����*7����.�y��_�!�fdt��ŕ�a}��M��A$�W�7� u�l��Of�Þc�~��ޭVTR�Xf�L�P��\��0���;Έ�U�t�c����@�QgѶ������z?F/ʫp�W�cB���U%��F�$r�� �v���Gl~�c��:�]�hi��Й	�[]�Iݟ��Cn�Ma�R������׈��a>��0zn@����i����~���hə�-�l��ޒ����lT�A�����̈́�gb6E�3�-_�LP.��z�F��d*�|��0�C�;oO!��X:�����G�xs��Tgi\槐c�p��wG�M���$r��̽��$r�u�_�׼k�A�)Փk G��6���!h7ܥ j�t�>9I��D��F]�?�P�R�op�<��%>��Caw�]�N`_zx�KZ�=B>$H�#&�� ��j9,�@7������6bX$�1���	�z�u���uHfT�b��C�%|�da]���%}س �:�;S�!�E{��P	~t(9�)4����´9�~�V4d\i��G�bT�K.q'�~n+�/����@�x3���}��_�Jo��� �>R���f%f����ݚ#`N���<+W����Y���F"���	�D�#���M��sF~4��dmH���G��2UG�
�d5([�\Tvջ�޳>�s�y�r7Ct�Z�$���i�����BO^#!h��]��2NZ�we�RdC