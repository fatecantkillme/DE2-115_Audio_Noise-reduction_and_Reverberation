��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<S��!O �&a�Y����4璻~௹���Y$�J��kyOYꕘ����	�����zS�Jb�څ>æ>_[>|��ϗ	��4�x�"!�/
`acY:���F��!�V�_�!��r&JJyu3����ZE!2?�=`�"�d�>�e�Q#6.�Gv�E�g��72�l�*�+��g�q�$��=�U-B�=Z��۸��Pl&�&Mc�me7�J��V�Ք��������
1?I��m4�)Gn��7JfEq�'�q?}��.wI�{��XM�[�ܸx(G���|�h&ň�71C����a����:��7LK���?G�h{�� >���^�YY�_�7�ٕ�>P@O|�"-��^�C5�GEKw�ڒ�Fȣ�=�4k��f�l�m+E�_XI36j>����=[]� ��8C��9�O1���w�������O�bI��TZ�Y������Ot_�r�����I( A{1com�d��?�r��n�j/�`���op��g1vE%.��U]���H
a�*Mݮf���ؿxlB.�����P�V��-3�x!�����4Mx����E<vas���qJXyZ�.+��F����ms��s����X�٣=��q#J�b4A��+��I�ą��r���4�癶j���Ų@W��wc^!�%�%˵x��qd� r1�Ug0~��4tK��-7*^�__1���2޳�l�"�o.��ՓS�C���
����΂�?�s7�3�vs�0���*�fY��տ���:�2�PVfl�R@�F��t��L�w�ͧ/��}�/a�ҹg���t�Mw��	26�q>K���;��u��
�}�<=Q�'�sw|J��Hd�i�V�9)3nŔY=�H�8T���L�"/�ҫ{|�^�'�v�r\�k�Y����;�[��T��Zw��;W�	��K��p�4(o���q���*ipe���׏���+h	�./����'�&�uH��I����>a�6��������[jlTw�����F��'t<��H�~�=���+�q�v��vP�Q^��sv����Y�Z��-������uYh�v��ͩ�כ߻h2o(V�A>�d��J�A�I3��X7��3�LG�Z1R��NJ��V:~w�\�}���i��f��[*~/[)R�PǽW�2�0�
��� N������T���4m�N"J#ߺ'�����8���\����ٲ��76���鸂�>@}ᢐϊ�#������K��ߔ�rB�9��k��h%P,Y��G�.Q�`�~��W��t$h��ԧyS�PB�I؈É�HSKa��Ȣ���e���'fKPN���h�������ɪ����׀Y���Ǒz�"M_J���k�h���f��SW$�GMq�Y:�#Gv�6���ʏ?.�s�&��*N
��v���+8@����-��1�7<rվ���9���2`������/^���ֵL5�R�jHf�q]�;%��"@�&}�z;�.DI����G���AÁ���u�IgZ�e͇@F�7�!a��Z��W�9�n/�А�W&�i�/�f�viP����ns�+5������!���A�-M`���t�Xեp	�I@AEA�F�{ е������aG��E$+�k���H53��V���p��֬��Q�cqCS����*����@�k�vxL�
yh�G�s��%��)=�g�����#�ji�D&�����Q�࡛���q�&?��  c��H�Z~QnT� ��
:�?c��[������9�:uw.3��+EG>!��	[�t2J�����1�䩹���-���1Wb��3}�N�I���A�-S`���q�V�ڄ��j��/�"0n%�:��^F���m�����|Ra:���S���gu��m�+���m�UJ}#hD�\_�f����{�̮b��B*�Nŧٛ p˔ʌXV��m$jd�!�.�jaK��z��95xz�[ j=B�@��o
���A�!�v�e���E�4�M(�M����;Yk�TN�鈚�H�-�,�mX��.cg��E���p#1�A�J�A��r��q����>��N�{w(`�$B��4�� ��JP���uqv��"�G���,�|0�yH���}[ɩ�F�'p��$� ��1x`+:bΟs��s�*�ґ��^��#23r��G8?h��eA�i�u��{��D;�ڇ�*�S���?lf��ņA�U/��k�o��d�A�Y���eɦu�{`6Z~��04D�;ʇ_7�v��D��"c�l����xb��~g�ݫʯ܋	�=D�˞�ހZ�RD�H�%�6��L~��'Ilr��5�O�,{ۤ�ә#�Av�(���f��|56��; �����ݝ��r<E�J����t�fCwH�Ԣ�d �啄��e��(�$��k% ԣ�yNˉ[�5���:�Vc�ۍ&v�������2Wǟ!J�T��+�[k]o��d����:��4�+��͛��)o�|����ǂ>�7(�Y)�����rV�ac{x�c`��+�S~�Ԧ��4?^�j$
gI��O�(�ód�]7A���JdG��`�8p`�߽�IS��.5�9uX+����!�� ���z���F\�&��(�  ũ��������LKޡ��N��KO�~�1�t��4����ڱ܌V��j������Z8�ڭ)�|��xv�hLşP����o`{�5�y%�
ɾdK�3�Vrp�B[��������G+-�s��tx�~OI90nD�=Ll!+�&Sgڈ�U���$MU�ئN����ᴲ�K����%����)F,T�M|V���@�y\c%q�7�D��X�F,�OjJ�n.m<�'�O1�Լ+�g4��W3n��N5K>�V�(kpe�o�s��vܝ2��Q���}� O���S4�z�+������g����\�p�,qafD��������P��	��î��������� �eW胣E?ĺH�R���IxЬw�ԁ�%-�SL�iE~�D�����g���p�h=kr�҇�u��d�{U+��@��/*� Y �z��a>�2�� W_�b,S�Y¿Y�S�G�!st5���lN���u �RCπB��m/�^�a:{a�%��Oų���/���p�:~
k�T�rF���� ��Z.q�d'
A���_��У�;��j�8�j��jO��?A�,}���W͉�B�u/�����A�R3>�F:i�ࠔygc����1�זky&Wħ~$7�z#�STZ��x�>�hB��}�Uy����aw����ٱR7�,
�j�X���NoT0�?,ʹK�+�0�� �T�09O$c �7�8���sA��>��O��n@tDa��=���_��+��.�g�1):+K��M�߼����ߙu�|�oY;2)�L�5f��w][a댡�*T���	�V��B��u��4���<��
KY�߃�Lt+W���Axwi�����8k��lBt�␳�%䪉f{�H+�a��
Y��ZjFG^%�|�m8�{�����gf2m�ԫ�N"�Ļ8e�b�*}Ճ�Eמ��V��?)��@r/�d��͈�
Xs(���H`J��;�<�⦊`��҇w�r([�['R�u�Kc�m�< ��$x�����:���C�����ہ㐙F=*Kb�p�P��@�c\_��P��_���Ep*l�s�	�
��@U+�Y�H�oR��c�PxM�@'d[�;-��׷��g<�����	N3�����
 �?�f�$�ة�_bF��\Z�}����xP�!�}���>���;�I-���}�8χ��jh빙Z"I�-Se���[i�+^ �Z�/� C�#�'"�!�U*>���`�>=<J�>q�J̥�VQy���'����3�_@VkW�b��v���g ��7�o:v�S��'c���yT�:]	���H�����	q�<��L$?6�m���t�v�bq�r|�/����3yLW��!$�*Jw}%Ea�����t�?$��MKeQ�,�e{�&�ъ�~�w�<� �8fq��v�o��J"�_�-��� {1�k7�z{ �K+� n`1��U1u����ړ:��BE���,<�h.�a"��"���c��X�.���ݺ3����%0��0�[�lEɽ���w�����m뤬�[��X���,}":�N�4��e-E��"NB�J�N��֎�
�!��n��I��7��&z{�?��3���.+�ȼ,���Ɂ�	m��ju���sԘ��|���z�C��s��ރŬo��Z�O�j�zSH\���s2��"� o���j)2�r�P����y"���v�.k}.|>���pP��i!�=ɒb?_T�ݻ{��h��}E�����r�	H^�G�x%�{ qmw�W�ՙ�� ����Դ�s5���d��ռ;�(�(��Uy�%v��~tf�\/G�&O�c�`�l ��s�1:�F��_5���\3e0��b�� �(~>�Ϩ�OE�Zp��o��+ﭷ��c�M����0�ɱi�jQ�����V�`p��ա19n�W��_��[*�s/~���_�V5&ߣ�;��n�Je.ݓ���@�)�3.�B��ɓ�D�h>���V�K�#ۊ��М�[��&p��$E�8�RĶ�t���$�I�;)�|9�8S|D�7��--�A��x~D�k&~�C?qf=�Ʊ��!�GЊ8�;���袬̏_�D�j��EJ�U�G6 +x^J8O�jU$�2)�Za��a�mQ��lϰ����M*�2�udC�hlQ"����'(DF"�������=��E�F��5N���m����[�k�7�!(��`����z˃m��i����U�u����9�{�d7G����ÄѠ
Q���ke�5�Q	Z���x�5�샚�4�e*^�z$�n��ߖ�F��{��1v)���w���6K�@���X�1����s�<��06����u9z�giaU+�®�Ɓ�m�z֚V�M�������扶t��:�w�t�]���/���S� ��;�)l���R�ެ?�4��@��"�PK�}���W����=IF�uG���32�Dlm^�˖�,^w@�Aq�|�lM�[���0�ҁu�c ��D���%fN�ʠ�ɮ���-,��Ӛ闬O���ҙA^���<�q��6�����RP�Y��s8|#7׻��?�"qV������E���G6�L�,.�*��'�����J�J	W�L��~��MQ��h��s���: .�o���7��!�77\	���RM�]�� ϗ��)�����
C� `����s����I������ ��ܼ�T����+]��yQj��1䩺�=:Q��<�r�m�t������j��S"�36�UTW�,!�6 ��g�{M]�K�O7
�jS��N�e/=,	1�G��a!^���En6��,��2���=R���a�<S�К��4��G/�]�R�Y��?��T��J�W�VhA%m���u�p��/	���(o���f<enaG���X6�������T�ɒ~g�ڝ�\�1S�� ������oZ[����(��C��&s.�P�4��Z�nI[�4�<� ���ډ%��cEADzO�$�=�Ƣ�y>n]�v�<�X{�xӼ3�,��9�@���d���B�wz�������DA�,������w���?da ��YF�Ơ�^m����/���7R촾�<�Q�~������;�[v$�4H�94� o����~(ׇ����R
f+��4=�<��]�,~������(���ǋ}en�ı[A�
������`,��!#.I �(�ܠ����S�����z�S�zLF"��q.mY���љ���$4����w2���=��1R��������$��	�Q�m� ��2L���������BǼ���0��H�f�<wz?\L
d���^�్����%�:�I`h���FY��;E��T�墶�b� ���e�#A��ԫK��k���r
sqUd��IҦ�ږ�ӄ#X0e���v��z��
���%n �����N�O����sl
���XS��ݛ|�ﯓ1�g�9"3��(U�?z�ʟ�51;�.@�'�!�b�"	i�f��`^Y�	��?�!��Cڍ���[�����t?o}�m��}f�z�]���Y��}!L�ʐw�� �P�6���S��:s�㙲�O'����$����K�S�@�;G$��;�L�l�m��}�� _/�?~e�P]0�}Gu�u��HAN�a�f$��y_��X��*\JE�?��WZA��*�߃��Ɗ�t����#���A̝YJ|7�W��pO�		uY @(l*o҄���F��q@*���lZ��\[,a��Rb�O��]/% Y�Ttm ͞k�a�^;�����C�o����(�؎���������;]�@��&�pIM�QU+�m��Fx���Ѳ�I*��K�;�6+��2ۈP���x�����h-���Al0�6�sydMZ�ܨf~��{�gɍV���_��f�Xv��QP�|P�^�)�c(�YQ�juVM���!�2hV�W5P�yV���k�Ux��@R�� 3��P[dSqd�뙠`��"����z���ԉ��f�,�w�JRc�bq~"Ye3:�t�ML�3J�s���	�4�ċ|����oT_SuN�N�?�Gd��/Y�Ȅ�iS; �Jͩ�N&5@V ����XtU�\b�=H �{�t*���A���i�I���Aҭ�&fCk�	QX��ŪN������$Fuhm�sd�U��C��@����{���	���o5��'�D��xb��&��#l9T�7�#!���p;wi��Rm�
}uF���3F;1�Ew���F��8��sAu��H�r����t��A�'��Pvļ��w��_�T�(���Y0(>_�f4�&�����q�gP%�.H(^P�`��Fݛ��Vx��I�_��M�ǤŸC���[Z��<��O��]*KY�M��	"5�񂧙��)��D�+�*،A�y��sx��G��]��}೜j{yP������L(s�D{j59���o���ƂuRm������2��q8(�)���v������}|�8�5]BF+���
���<Ұ#׾�ͬ��pуr	1��V%L�kbC/6��.���fV�T|��[�`����Y�W����p��e�6J�-ě� ��m��|��e���'wB�X��7� t���VKً	2�7�KŴ|�o�?K>����q�O*��?�U�Yq_$�o�gY4n��otyWO�h�ݰ졽��Ȋ�6�J�.��	#os� ��C��ԕw>O�����akO�}�b�MX��w5�0S)�1��xpZƊC/�<�9���؆��D�����fG;�$d��,2r��G�2U#��|"�|��߷b��xR���6c��&���5����Wy5=$�e�><f�,����b�-PEqacy$���Z���sr�
����f+Z�o�r��6��Ẉ��m����z�$ܹ�_�5(
1�$���#�F5ـl��o�*�q��Su3W��$Fox�'<m:W�%���i�7�9�� K����F�7!aG�=r�A��w'�;;��p�"ֿ�.V5�5�:��0��f��z��3��a|a����rq�u����5˂]9��i�C��5ݪm��{�b>n������#	�Bɝy��~�:���!Ԓ�n#�<�n�VY��5�W�w����4f���W��.��V�p�(� i@M��fŨ/~ݍ'���i�WNTs�b�X�x�顿��Âꋄ�o�`��a������Bjeu���{^G�V' j�Q�ك���0=t�"�_|�w>ãf��R������A�Cc��P��xe!��JU��|��1�W�o��*x:��e�����\�� ��q�O�g@b�4��,��l"���g�j�[ZHRĤ��qY�F�����&@�?Pr-8Z`��4H�� ��J6	{=����D=c��u��M0��ܵ��V��Q����B�uL'[�'^���V0���L��X�%t������8�M3�/�g�"֤r�&_d�S�}���i��e�/�&�jsc,�T�/�_Q���|tK����+��s���9҂gi��b�qP�.1zbz�?��w�ˆ�x!�f���WC��}��ؾ0%t��T@�u-����c#[�wr����}VH�[L&*��,?�ހ�_˟��S��n��bmP�m�9�ê�EH
��¯ǀe���Erz��d��7"J'�7�Ұpڼ�C]�N�&��Mϔw2D�[�\�f ��ɽ������s�P���l�Q�p�4�>-/���nZd���h��:[p��ꃄ�&�5���ёM��kݒodo�Y,�e��ت�^p���:�U#������T}'r�2��M��q{%�>��,�G�3��n8.�d�<#�J&"��1q�M>�T��,�Fj�`�s���z����M���o�~ T�U�Ƿ&o�r.�W���_�b��2�l������sSI�U��\F���)!,�pP��Iӥ��OKԚ�M�x��AYi@rq����<8���^�r�}�1тj�h��Hk�c�ʹ�z��o^MI4.�[�!�� �!)�J�z�q�-�������u��	�A�y ��O�î��l;S�#Ƒ�h��UL��D:�=T,��8hB!-���/,.�+�a�[�Ϣ��H;'\vȈ�t��9��ӯ�����O�Gi�Z/8�v=��5��(�b��V3�*�����kڣ&[��	�ξ��������d��4���~Lx׷K1Dgaǝh��Ӹ�.�Ò�7s�L�]��ś�����)��@�	*O�=��/c�>����:��Ꝡ�K�;r@��{��㶱3 u�I�{W���s��Q��E�H2ho�E"�Q�-=���	q�۬�ڕr��Ɔ�O� W.���^ȸ��8������'��^�"h?w_�Dv��޹w�K�Z�D���?��