��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjfm~���*9&ʋ}�T������%[��Уt�'�}��������l�J:��	�gO�p�?�LkR{lmj$��H�����ey���t�@��cg�/�\�����>��`��0/ⱳ$���R�� �K�� *���g�Q�J2'�	�=d�E���ϠN)G99׷���h����cm�x�xI�^ٟ� �E������狳bֿ�h�j�T����(Ο7�5'��Ҳ��ǅC�tbN�jx��7Պ�}g������`�[pm�\{?s�J��������]�vIE�}�:����͚���g�$D�6����:zZY����9_�U��Srs=jc4X�J;�qs�RC��*�$��B	[��{�C3qHR?l�^g�+7�Gِ���z�.��Tt�S�U�g��q�J��9��7�RkդcT��ǳ����ĺ��� ڹ����*�a
�E[�ey�5vw��_���R�v��^H�9(�&�!`> ���:wp,s�w��`:J�Z�v���	��	z5[)9�Q���<��	�/�O=>�f1V�/��O�f4qN����Íj ��[V�0�o��:�M��c1B�����C�����vs�ǌ���Z�;>���93�@G��\���21��z�C	P����hWpѕ��)JQo 0nQ��5F~��eu�`��%8d�b��j�Ypi�6K�"_�8��F��U��u�K�������<J��\2�j��EFD*��V0�q6`5�{x0� �c�X��ډ�<K69�O���!-Q� +Yw� l�òx kqR5˕���w�a�b�#�,���W	�����<yA���&�AGtc4|B�>�ԟ/��[#���̉���!�(7-��X{&|Wxֿ�4�z�6(��z��<3�"�s����<Ne�YU	q6�Dh��.�p�o��n���t��YH��ϖif�����a�����-��:�HGq��:�H�*�(Y�-X%�������Q`�#���X�W���6,��_�j.��_�5��Xp&��p��D��	xw�C��Ej]��Z��(Jj.ꚑ�7o�>��=��1�r� ?�2o�	��6�: r�5�����gӤMhX/U%6XG���Ր�w���S׉�.� ��A��8%���ر�M#�o2��U�ݢtb���'S���y��"eq����ev��G~�	�"�X�������R��ʕ���*�5�Xō�e|V�*G�P�(iw�-�yL��Ѽ?��⎉��t�fM�7 �*�L�r�Д��������N�J��8Z]��SV��FYfw���ƽ���o��zF5?�1�$y@[s|����gA��9�����τ����?mc4n��
�WR�	R��M��ߩՓ6��b�
,J~��|*���ϴ-7g"�1�=����u������cXF%�ɺbվ��%�`�}��3o�M@�91t惉���>��iY�\�f�:;֌��2{c](7w�ϣ�Q�	z6�+"�ߒm	F��3�����If���L���M�{�1�W3�J�Do�2��!N�2�2F��������e��H�,e���������1- ��L���gUlZ�r�Fo,c��vQ������i��T�u��Z�y�x��m�C[a�d�͌��SY���pMp��]h)1��2��Ŀx���#�x*��{����Q1e��Ј�
b�5l��]!����RR`�vO�'*��֎CH��K�N��Ά�!3T��~Υ�g��=������r��!�Ac.5@�Ү�ݕ��c|Q$�? �'b�$G�`�����Z��l�7��7�L?&�:w�R�t\5���y$���B�x�A���I���,N�|ETL�0�
������gM+�� N�wP>�7t=��q2�tؖ��v��r�[�1+�Ό뚦Cg(�㛣5rE�
g!��#�YZ�L]�\�C�;+�4c�F��VQDh�1i*��\	��� �����u�'/j�(T�B�uTA2&�9�L�R9-SH�e.�=ɛ������>r)`'b
_��pfd��< u�t��ߕ- ezvX�s�u����p����~d	�=
,��޳���)p	;�/!׷�X�?�kVc��w�ź) 6;�3-���rP�hk)�M�0\Y'��^���t��q*����=�p!\����6�-k�A������F|[�Y�{L���i�LEͩ.�r�r�zT��u����2dF�C�H�q[}��ȇ��}��9��L��΍���!�Ba���s���U�������ill��%��`�x�ތ����3˂������`�mؑ�҉��.�)0�R�'��K� \���f��U��9��5a�B�q��e�F�*5�����r��װ0Z��+�r�9�.�@y��{���P(1(�0�O<�D�g1M��0��^�`n�!�k3�
A+p�]����·v����A���P�����*��'Q.���\�p�.����~���9��3Xдk�
�Ƀ졭�LY1��۲N��cn�fY�4��:L�pK����𹝠�h�=�bo&\�P?F3EzJ����M)ɡC��m��F�$�lL�#�T�kԩe�oc��E:�"g�ѭIs$�:�S�<���_*�j���3����%�����5?ǉpc+IC�[�|+��e��o̱��w��b��ρNR`-��@��D�XMj52��74��Ο�R3
�R�� a� he����O�rgm:��Q���C��c��j��iڟ~�ig���7t����� 7�gެ<��6�b�')g�L���ܐ5[+�ޗ���Nz�N�����V��;0AI��N*�X�U�j��L=�Z����=���	�oK��Y#?@b�M�{�)0����� J�@�٣� 5�k��r��]uB�^�m�D���<t�����.��YD|p�4�@�/Kp����A�ܭm'o(8�`�����@<���.a�٥�U!�|�����Ic��934QV�N��V*��.lՑ��$�/((NZn*|��Bɩ�fm}��Qϛ�"��/��o�G���W��9|��_K��H<���M�j��/�C⺗�+=)����d�0�^�s�@׫&PrǊG�	�VO�{8Y�J��	bL� ��3MPE����SR�b�~#�z���0�DD]M0�V��ŃTѰ�h���R�^l�k Ҏ$�����(*U��M�9 �Q�6uƘ�����K�Vo<͗�����ڂ���Ț��f��\8�Fc��:kC�)��U�95��OH΍�O�͘�/�����}��d��+��\���r�βh_
�\���q� ���f�����-J���Fa7�Ch �����!��x�{��0i"<۷1G���tVy#�a��P���@6/�r� I=O�!��6[`��J����JHD��ZҬ*�c�$#����%��
��B�ؒu����`�wSD�i5�u�=���me��: �]��I�us쿿}03�g�J2N!WT���D>���� �,��7BYA���eg��,�E�ih`2�ٲ���H-��|�r����Z�XR  �Rz�S��A�l	j{��E�0��$��0+�^�sh�^D+������t�g�Ln��
$֝�l��-{�~F=��	��ą��N��7'�fW�yf
VkH���[΍ d�J#����.���7�]ü��Ā]��\_����b ��i^N*�` ��b��U�i��<%j�|o�+��!�ɫj����#\0����ʑ�P5�0�4>.�#��L%�1M�rP�ܝ9mJ�C��"���&yQ��<0��q�**�k���l�T� �x-[$Q8���Ђ�?��4XLP�M��B�ن�!n��P����$��;��������֣K[E-��僩㥫�kk�U�-*�����g�o��G�"l��:��I� s���>�a���|DR�sU&�������j�f}�*a�I�\�.&�Z6�]�Zh��u�ڭ�ub0�o�lMt+�:�~7�zXCz�L�k9����{�Y�Z�l�#�Yhc��A�E^ǹ���68ԯ��>]?gRu����A`zZ�%�wY��X4S=�J�4#!dv��B�̧jv�\Zşƿ�wҭ,��?f>�����seH�#��I�ݓ�_ �
ב�O�/c�A���8I���r�k�Q���s��<�<8Ɓ@D]�P��V�3͍��^>�������k���Gf2v�F:��5anɞ��cXv�B��Q:njc����s]���u�2
��p�s�����'mjՒ���[�m��X���!m[�����f��W��昚"�/H"�%
Ы��o�L�f��k���X�}�2�/�9��#*��ʡnn��,��o,��<��ϼ0֋���O��re#�6ջ������$�45�L���,ϡ��(M�En[n�H��1B<�c��q�LL�\��V��ۨ��n�X��֭H���l�o��;�v[Zz�1��[����e� ����K���n�����L[��ŝ+�gP)4�� ��I��w6�v�@��z"������~��"ܼ>Fo����X�ѩ3�60��`�3���7#t/��X�����?"��u�Mf{�4�����e�cn��d�@��NM��L?I2�Gi�{�i%V�����0�̼M�f���e�Ƴ限��T#�;�os�P�K���Jl���5ʺ!3m�d�)���lL<��>Cq
��lD#�F{�w���߷k&j%�3Y7d[��2K����iȊ�^5Pǈ� &�W0aՀE`��3�R��P��#Ri������Q�&n����݌B,�y�z��pp�����C'e�J]H �]�$����6��<K_a�p=�u�	��S�Cܾ��3\̆�௖#tN���܇\�tېo�Tm뺳���|T����b��uh@u �*#)+P��_e'���t��@ˏ��3G������4�.�ۥ���]�
�ո���0�����A�?�7J�$���g&�%G�|�.c�G��P>qH
'>�qs�����p�Ǧ�r|0��ܦ��`�����{Pg�0�s���u�A(�����J�_)=Ũ��ZB�ދ��g���
3�� bg�2��q'�A6��4�e&�_�{F������~�E��
���b��9S�_�=pw�|��O�K��%�:�#�\l޼)#�?�K�ʤYwg�z'q�s]\���C��1>�����À�w��[���Z*�s���e��h���`��L�0)�Ս���L�ώ������%܌f��f{罪e�:	�2���;��j�K�Y���Rığ_K��ZЭ|�MLL�����g�n���޳M���Ǧ3e`��.+%��Vp^��Wzi&)�����9H,�C�y�e?��-Q+iП��}�iJ���C[w���6�|j`2P
��~��m�Vc�}�N>������\�)�ң"���۹��n��|W�ne���:x��z3zP��Hk_�� E*�S�G�0���m�=���3G�3eQ��j��K<񎖮b��u�FR`��1n\Vcg�&k{qE�>`�CA�s�Q��ۣx�7m�q�n?��X��ҿ�m�R
g*7U�q���"���=��ŘR%cõ��坿�,��_`�����U~v�~��_�.�|�D⬭U����<^	��MY6���{��"P ���n��S�n��Pő�8��[�;@M6aX[q��z}a������Z}���qt�\��z(ܮ�o~��U0��cd�6���a�[�V~�A�)�Iq�W�/2�t����+n��R���{o��<H-�~2��\�tg)<62���!��r�f&�Ƴtǚ/��%0!�v ����V?�A���C�������&V����ڨak������c:��&�h�L>��Ÿ<Wy����=�x�1�״m��ܟ�q�7h�i��~^:��
!�8'V�Xi�b�v�r�G������u�ބ���Y���>Ѩ�M�d0�S��Ffa�2<V��h-��e�5��z�`Ĳ^�e�=4cɅ���*zȪ�e�#Dm\�@h��$�D)��q}�pрH���"��R)E���d\���6s���SD�+}4`����I�B=K"��C6,1��4(ٮX@�R�������h':p�J�؜V22� S�D��c�Q�ē��"P�>o�pG��D�Ԥ���$������UhF��34=�9AB���v���o?F��}�Y��=� H�Q֡kJ,����R�'}ݢ�u�h��4}G%�S��V%cW	��s��gxzpE�s�5���z�S���,���ލ���Z;�0�ҧd1e�c��*�r�#�����3>.�p�Դ�q���'	��:��	Z(h�6=��Ej5��Kس��[=DJ�?v�y&T|����R��5W��A�z�fߦ�Q~Kˈ��9(��1.s%�A�|hнoG��cr�KLi#��ʅ#��y��Xp���s��?	Q؛2�n�����=�@��*�S�s��Pg0����xƻ���QVN�;��y�&��S*�/�z[S����'1| �OCd��q0H�C�CSL�r�a���Δ�|n��1�脺��,���2�.	��6ת��B'�@0.Z{	C�,���cn����BC���I'�#�,`��:Th��ݐ���X����5�� ��{:/��"��E��}Bs
.��m�Ű���u����Q|��H��Z�l>��V��e����R j�P
C�ì�M:�x�"�="3��$�ك���I��^ճ[0��X�{�7,unk�|��Vt�W�4�<�5�*���m�͇�f���p���$�b�oW5��!fp���-'F�6f_��P6�~����5�M���2aigy� �w��t״�ƥ��Cp,u�l��M<�G�\ J	_Vˇ����_`օ�ga�R��?�v��#y	�d#p��X�ުѪ0��KV���_�	0���������]��3}��5�-KB���F�Oa��X���?E�c�9����4�	���W��t�.���]���O�K�6C�fhŢY���`�}�`xC4����ɺ{�>��&y;}�u�/��9���'�]ώ�s�|i�ێ ҫWMP��^l9A� ��Y��uó���R��b���|ʥFă�,��ݕ��RQ�Ə�3�Y��jԡ��S2� g�+n??f:�Q�H9�������	��*~�VK��n��Ҍ_���L�{m�|�K�J{�2�C�:YtQ����ic�z��Hw�sj���ܑnT/%�c�����&&�~k�\����+,8�3�o�����G�fc�� ��21Fچ��Ң�۬t��-��7��ʹc�eͩZu��}Q"����#`2��]-[��{I޲�ē�V{�9Tt��XPܳ!t��NL�:k�EU~��6q�pч����Fc��x(j����AL+����sH�>-��1`�7����ۙ���_Ѷ�A����Xͬ�ٸ�f��"��.�Z8�?oË�\���v]�o�6�+.۔n�.+�3 `���i�F��6��W0��P�CP�c�Y���L\�y�O�C����#ͅ}'v@�j���㏬`R"IΘ���i
n���ÿ�R�����ٔ�?zj�5��f{1�9����O�ʱ�#�D���-#�+���(��Je�B�.���E��0r:��
]���x�V��s���x����s�_~$h2�^ܛ��xx=ϯt�	�}��9@�Je�$N�[�Q
��mL?��H�(h�L������
�#qn�pw?��� O�i'�!C���8Ng�}e�a�Y��k�e������̌�'i���J@�_��!R�)�����8B�R\�^@ ��r1�NM��C�ã8���Ӥ@(�۵G��a⢢��%��+������Q��;UNf��p�����~�4���sZ������@b~�@3��;����[��i���2��K�71�Q��8e�҂W�J�j�*��Mf�Ȫ^=�Nbm{�nJo|)�<��S�^R&M�s�c�ܕ��.8:�λ�O�٧L��)�#��/%�k�Q���ǎni:���������7�����e�X/c�̚8R���Vq X�n;��WU�q_����!׌��߾��ʍQ@q5Ѕ0��y���پ%)T�2b{#��OeH��r~�H��>��]s�oxް�{�0�P�o֮�����?���<���`r-��F�q�i�()��E?�T��1�r�p}�N&B������~�,h?��mn'�k�Yy�:���P�c^�Ǒ�̆c�����gw4��4Ac�������Vl��0�&��|�~�)��`/Υ�"��ǒ$��E ��t]?��ӳ�ܚ�66��N�3�|�M��|��Љ{���b�m*�9H�c�Zc�\{��L��E(�e[���
� ,��ۇޱI���	��y�}��`��᤻���KR�m�9�.�_���L�����r���q�/���v'�\q̹���BE�5p�>��w�Cr��g�q���#h�W%DХ��N��T�(�Ҹ=o����[���V�+b�0��2{ق�h�?�@H$�*���s��:?��~��_	��ZL�z�c�i�C�)X{'��+3tA�\&�qH@+�s�U(Q�H���ql��Y���y�I�H'!�.1�K �w�K�� �\�am"� ��������Gs�8$��1�V��00��C3��5-S�W?��6�p�����љ�4
۟����1��F�J�0�$�s�]����#,�X1�R��6^�n�$z�{2�7�R�>(@-qԳ~�hb�e�R����<��R�N[����յ0�Uדǐ��p'J�z+%�J��A��WV����w�YsUp�i���ͭ�aΣHK6t'��z��G{��O�]��H�ջSHј��8�[�D����|B�y��*.눈�6&%�	����GȆqk��v�nc~���9zү�v!ptf�:j���v�h�b�~��+���*m���n��G>�?�|�n��s�ܧ��1^L:��#sJQ��F]{�W!cv�m������8�'�n�đ�2�"2c��o�� N�x��I�3޼�V��t�6(A֜���&�S��6���p���!��<�z팝� �*�� p��}_nl���OM(2'�M�L��x����ue�v�s�G���z��o���c�B���,7����	�To~02��
�����=:�K��J�����r��������JKP���E&��f�	LdZb�?cJ*2��@ʊ�����T�UKQ��#����:)��~%b
�mіWv�6����Ƿ8ۓ�`ԍ��UPb,+�s+{���d`�ȁ�M./4�vTI��ɋ�1D�T�hN�9X��/k���������B�6?��/e*)h��J":���o0%�3��4���2����m�����{&�ɥ$~饣M5K�*���Yg���&B�M�]1aW�(���U��<��6,�܃�C�$�� �J���G4�sP�[T�K�����7�d$���ʤ���O��7�U!�7��4齝]�b

��'�[�]��_�k	C90bYU;n'E�E�4���b6˳��e�v���&�o���HL,S�:��*���l.��xH��!n�fv��Bbٕ�-1M�n�?Gw��ML��������Q�P+�R7;�t�Ù�Z��tY�n���6�&��3��װt'�U���Ơo`b��ЄÃ/Ad�_w|x�=UUĪl,�&8�=���.��Sf�y�Ud�7晝�b.C�h�$�V=1Li�9t�[��bSJ15/����~�ߟ�-.��.��2o�Rى�P��)l4^�!Yb/m����\�+�|(�l��k���n�s!(!�������e2F��`o������P�5>��:Q�>}e�Pe��k�Na���%���<N����R?B���{*��BՖ@����9i�݊���;�^�����=�mq��GH�����uKۧ�ZN�/�Vˊ3�<�<69.ݵ��ǌ�����\��8��1L��0��xI���c���u �kD�G9�#N� �ڙ�J^<-͔(6�
3`���q�-~r���ʹ�K6Xf��e�ICCGT&JS�[h�i�B��n�?��8>���6{�F�'��3�&[��Z?@�I���X��h�ƹ�Lu
k����ݫ�<9�enL�D�h%{�H?�ێB�;�	��_��.�[W��R��������J^�����u�@���Reg�BkmU��0h��CҶE���� j��䰖u_0$q� ꑶp�� ��]<8��%{%���U�]��aՆ���F8%�Ѣ!��bXZ��! a�6 |J5C�JR�b��4>����?/n�3���F�x�0�BL�g%��N`�ew郠�;FR�_��h�tP�8 i���A`�Y�9��!�[�)Zd�#�R��b$z'?�&,�Ip.���K̰�7;G�U��v%c��~��R�!Z6dH���ť�M�w�_^(��zv%�wX+'d�1l�ޭ=��ۮ\�H1,b �Y:Rɾg�-�}�=�����"ֻ!�yo��I5�1�aA�Q��O��%�l#���6�;��z�����.��{���0
�Y/�i�O��}
��ߒxM�9�'��ጜ�fc;	hGF@j�����<ٗ�d���&�Z����3�
)5�&��-��e�4%n���/�&	��A'O�(��4���������cU,�%'WΉ���h"���/��9�(n�d�'� ��Xh�ƽb۞��]��B���u��|���U�7A�~]n��L?`�����y�I�rhHe�]�3{��� �z���^,&V��X��r��`��`���x�I�ɳ����E�ƎB8K��gbzT�*���+���� *�f�	ş��J`R���|��#J�!�Y�3QC��G���n�,�l�X��~c�c�p�9㑀m�Q���8���z_#|^aE3�xʟ�m�ߡh���d~��P/�^v�9��Sx����TR=a�>	�Ϭ��@9���bx
�0�ң]Hf�@n��7V�lP3�[�ȇ̬)�O��"��'Eg�k�z�:)US�~}]e�5sV�O*N�S~,L���A	@�	��z/��8PѲ��<h���<�3��9��#�Z���W����$�G^)[��4C̾
� �m�4��Q���}d~q:�TS��iy��aH}=0���T�^�13��T���dg�/�L��~�)O�p�.�h��W�
]?����*�Cj�VW�/�"2�!1�\5��o �U��L��q��:w�m�E���7���XV�H�D.��o+�e�:{Y՜Sē�����k��)���Y����m��	|�L6���؈ΪI6��B�´��xy�K�a������TGg��Xέ��jK'1$�fa��o��/�\|l�fW	&��Q�Ɏ#�9�
��������}BO�ώU�ů�j{U� �E'�/���m�1gwVA���>����7!t[�o���_J+)`��zZ!xW8��ljZo��c�B��}�b�S�oh�������z��tF�K3� �)��kD����9N��*�gH&�'������n?N����nm�W:���#���n�`M�p]�o�X�,�l����˓���n穾���.�����ف" Hy�P�/���6�=<p��[��N$]�h���N�lkHӇ�zȐ�U����P�׵o��s��{���'����v>��.^�����'�F#M_�@3�[lOX�^�D�~���Zc��f���<�m`V!qO�f�9�FiLK@�T��@�9��g7��X�H�6pT�����⩝�_��fX��]�Ԑ�;�ҧ����NTC�U�p#I�"Y��~��*P���A$k[���#��>{Eu^�8�Pg m2�_!�K�.�^�j��������X��Z#\��e6��?k�CA�4�\��W�BU�:G9�����>�؃8{���&&lMk2,�f*� S���2�]��Շ�ł���5D?Zf�v��*��g&�e�Z�VKt�C��*=
���Y��糕�D����,Yd�����O����./�W��8�M����_���(K�ՙ����墠xz�q�����qONԔ�g���, �[�k���΄��9�S�ܪ3S]��,�}㓡��x��k�a\�4."��So7m��; �U�OO�l&���YSluO?q�aY/�%Ǐ8�r�=b���<�Җ�/څ2��T�8|�js%1Yp]*�V"=��$�����/DEc5AxT��EV?8�1z<�����.��ޢB�6^��ѡ�+V����; ��h^�y�y&�
�e����Z.j��ޯ��F��p�#���QH�Z�X�����u�j�m�v�3!���"��]e0MuEwΧ,�|�e�qJ��Y���-��6ѹ�����4B���CLT�|B=j�<O�]o`K�^�1*^�dJ�k���n�\H~?��ݺw�Ӵ�f`Y���h锄*"�V(�Y�-��>��|Z[)j<j�99�iN^�\r�KÌ��bVjC���[d�nKc���-���Q8�Qy�	�aMӴ-'ܬ���(rL`0�S��۔f�mh�çt��S�}��y˅��ne@�+C�8�Z����i�)*fȫ����n�dX�k��Y�e�¼��{�p�Z� ��Ќ�ĕ�IY�������F)@����̽�n��;�i]�6�G:���N>t�:\L5𧃞	�ų4�����?Ya=<8�V5v+Y��������R���y�w�sw�&S߻�9��X< ��hu(q��)^��"��2�']�R�B��N�ŰD�)mɒ���M�|��B-���C7�}����G~2�%M����GFڴT�'��qN5����[pk��o��]�ˍ\y7�Z�J2G���ڔ'��8,0���B����o��.1���F|�|ch���.��&s �3�z�7��V1@�_��[Z8]�h�D�����M\�ݕ��t	��AF���N�~آ{H^�W�����D�蹶��_3qM�+�9�����V�
�s�%=2d,�LV�)p�3׾]��Ƭ
z���Da�h"r	""vܚi������y����Pt�w0�	�%� \Lh"�!B2�{8��s"�����(��nY�3[�9'ڃ�[�
����*�M�`.���)��F�[�Y�V�6dt)�7'���l��J�=[ d�f�@��挏u�{�p�ؿ���H�yF�E�?���(��(��J�/�B��]͆^�-18]v�n(�J� ��h���u-�8b�l,
K����fq����_To&�-�V��t� ����I�l�^�y���whyv�s�*�og8aH��Sx�%��(���Bv�F����)��;��5�K:����Q���6���)w�{�Bƥyુ��;��UEMR�W�9=�Z&�,J�ϟ.|��.Y����c0/�H���#@O ?��M�����-�'��^Ɋp�2*����uB����?�{=�Ӡ�w*�=�K�l��������Br�KW$e̱��bc�W��sz�#�pw��̥ ����uW�O�+�I1={�]��`������S�>�b�	���[�Uh�ʗ�]@0�ư�&�Ys�� �����N�:�r����$1	�p��PXxն���ke�i�G_�r�f�S�=6���&��f���-�	:��f�ȗ�'�m���R�������*�{�8�IV�D��e%@�2د���ô��
�#�q���e��ŝȒ�SŵЎ�@�j�QZA��-��
����-�R�	e6ە�Vf�;���5E�� �p�� �vBL�_�2��W�n����+�լ�ظO�ɰ$J�l��Z���lf%(�R���λ��F_єzOEZbX�i(_��Y'�q9C�F��V��l�S
�_�e�[��ɫ����-��������0q���b3e�Q�K�3�p��<�D21T����@Lgң��K���~����O�G��
�����=��V��� ��q�sT�����P�QÈ3�R�"���]>�9�� W�G�ya��s�+��UgA�E�ҋ���8�4j� �?��g����g;�o���-?�ȓ��w�%��c�]o�M2}�B}���iu˔�W���$3~�����+�ʫؚ�F���^ d"����	"��璆��I��������tM`D�2�O�]�zC)7���@�^��w��μ����%�f����Y6hv�{4������M�[{�E`��m�C�lZ,
VFT"/�y�s4i�z�4L	�Qrmh���ȣ�f��,
��/!d�d����qM��1P0�MzҌ��(���¡E_~Ի�<�I�O)+ ��I�kc�:��{��`�X[��W���ąb}`�j���PSL9���j���F��`w%��Nx�>����+�����$�7�[&q�y��ݣ�?�h��o80����:���4�ku� %SB׊��w'�8��bT�O�V�u�eA���"3V?��:jJ�����Ar%Y�	zAB�eEF�[H�����8#IUA���xb՟ZP<c/�0R��s�	��s�-�t�&;�H�r^`�r�������:)Jq�"Q
zb<�^�Smp�O�瑚�"���G��B�%����H�zМamր�/\�}R�ȁ`r�!��vN�.V����
�~�F_�M
aa�=r�`�M�Q�}�7h�f���Uۏ�#�:�a�4��̎>I�f�W��<0��
�j�R\b���7��B�=�8�g��DM�0�ݩ$x9��]�����QPuv��:�"J[=rr�,�-����钛�a�z۞iw�ߓ���I�-k ����0���W@W��.���t����������1�dH�F:��� n.C^�n�U^^z�(?J���3"_����?_������Q�I"�U1zy�����bv\y��;�@�Kٜ�����|��왖 =eb5c���u�V���u£�[���z������@�'�wY�qYl�����~�M��������ydcB�V��i3V��x�3<H+iF�&�����y���4T����I�V��z�L�[�#� [��O�-�`ߑ0��h��Gó�$un�)�� P�Eh�v"6�Z#	xs�I���bF�:ا��^�,����KɍJ�ʎD<eQ�.�6^�����.�<{�J|�)?(��uT�Z��zB@��S�\��*��'1�Vڊ�ֹȒ�#Lh�\�c���=42 mtS�g��5[��-��=$�'�q
�w��G���x@�]�����z̔�YjE������J����/ow����X�s\pf���u11r"Z�(���呙�YĐ�|p(6�i�Ѱ� �Az�����T`�Q��q\9�����~���T�αH�((ZH�ڢ����e��/�?��F䜛{��
�ഄ!I;��R�V��nHxKx��K�Fr�o�e�|��Hp���aQ�ϲښ"׫4�/��D�J�k6�<�/�#�O'w-���Ed�3�{�tG��.<Z@P���b���k�h���k��q�P9V�ދ�'��q�ŗ�==�iZנ��y'h`|��E:B';���m�v\ee���@��+\㜥=��y�<�iS�} )5?�-Q���˟�3�9ى��~����<q��6f�^���0.�~!���>�ug�C0�(�j�e��$��� =冖A�}������2ğ��w]Z�`0�sE�fg�c���e���wrS��s�, `09-O��4=}�Qyx^v��n�ռ�Ȉ�r�P���l�����'i:�*�y�D~����}�P;7���T��������0��cq��#���I{j��m7���@
d�G�O���  &C�7%��:A�M�F�z�+s2��$������o��F��âb��K���쩸��3��m�@\oVMk�>�jO��4� �<�$-Ш��8�}���u~��	@���߶�	p��td	3Ӕ�I�?�ӑ��o]����J>E\v��8��_�
L��ļ��v�{�/<,��8�������<��?�*�yeYֽ"�����ׇna�-	�I��R#2�:��ê��M�߆�x��8-�#R�G��/�Jpw�K�c�V�r���ǎvPKg#m',�)_l�]���Sg�a{���m8B�Θ����ę?�QȞ�J��-f�g�4��=,�(d(��i2�\"���l��Ӈ(<�+�!ji�� �|!=29q!��:>��Ӿi�����CK�C�ij@m/A\�*�E�f:�é���M��oo�^��̅�aN�X���O�i�uA�;m�m��p<� Y��_a������!��3$�xks�_Xr?�l��9'cXĊ,)߇��<����cz�]wB��!NK� ���.QQY��Y���$�.P;��s�<�kue�S}b�����юw3�=\oV���u���_�t�����4�i���M�B����	FA����u�>�Ʈ�N7�4Oa!`�w�JL�	���^���Ӊ�7[J�����>M�)�N@�Wz�ӪB�����1JVv�`"*��`5�Y�$��A��~A[��.!�Σ���I�kB�����-̾�=�o������>���I��ٻT� ����ғl���#J*�� ��\+ϸ <0�'rݰ��o���s�����p@����G\8gw�XިH��_��A�L�����9J\hȸ��~�i�J3a�ȥ�7|��ϣ�&�bC?yo羚ҷ�*sJ�����%��!���I��`�k���J h�aƧE4�cH��K��W묊ͦF�72�$F����}� ��W�b�[s���r��y��-'q9AYyJÛЮ�����uȲ���3ߨ ����j ��ݼ3��G[!�!��E��ߘ`��(��Z�H��G�����9�5���Ӡ�_	!C�cp�z�wg�,Eq1@�釓�9� ���
6�����oD���K��75ۗ�;�{��]㢎=o���_��q%̘!�p��vy �@��>�>b�I�@�9�G��4�:��w�?2�a�mbW�×>�W	[�c��Ĳ��N.��r�yJ�aDA��w�&�nE��οBF��Ԟ(b�6��W!��q�<�zw?���� %s��.�4�{ �5T�DtV\$8�=n�"�߈��N�`.�wP�U�t<py�y���D���z���#ջ2�mfz�N [��W���ƅ&O3�	!QSM�?���\�U����*�Q�}ϒe�WN����½�@'�B�8
^^��1?�:�gcq�?ݫG�J&�K�C
��2[`�k����G����jT�N�[��ɳ���W ^6����cu�W]�B'�D��8�|U�~� �bygMg]/`w!m�G�(�p�@���u��s��(���~���rg�c��3k�W�d��+s �[�8Gl��lɔ�R��(������ា��h q� ٢	1y�/�Z��?�x�.&n��WT�-�zW�-\�6.����5|��_���L{�k�Ԥ�O�rN�qۧO�q(��'B������ �%' RP��GdTi^���"�G����N
Ҽ�d\������"���D�L,��T�fT��s(Ip=�dX�����m�ǟM�1dD�&���I	�LQ�ؾ�W+��^;-3]�q�/8L�|���b�d����@�� ���qx���; �FT2�*�����6����� ���eQ�M���
�����[s��cE$�#�Ŗ4�/9+����zM~Ȋ�F���BU��ђt��W���k��$�F*�8$Kɓ��v��������^�Y� �	���|�!���P�Vh��6����M����o�՗H��V�5-�n�d(B�ٍ���ʕW��Գ�HtG�Ҥf�#�"2B��K8���u�f��AU���S��Po$�[-�T3qBȳM+e}��x�[�c#�6(�^�.��ڗ��~�LF2��!M�L��Sd*J��	�xڏPt5뉨⳾�j{���4[*�0'}`�e�*���$�Y��/2ū�~������ �t�i]�q������,��>��� �����n��UOii��ԍ��9ae��j�׶BI���h�¨x_+� |�x�xa�i(�3�H�!��?���&��:�r�}�t����զD���
�!�:���z�����Z�#3\5�~�B��[kp����\/\H�oԥ;eP�*�%Y�]�
!���0�<4%�A̰��oq��17(t^���$F��z����2��~t�[F��:Γ7��Ϥ��P�,���$��l��	�ѧX�o��_O�5x�N�>Sz�	��N��G��[J��N/5�i���> q�J
�q�a���P��P_�o���T3g�h��#͕��L�n�i�po�Cn��\��9�!��Cց~��Ɓ��v����.S,��;�6�8��>��軇��,�oY6�~����K�[��22z)���iw�li@q�$ÃftO�vD��p�@M��.��1����4����a������+\Z4�m�\‴�@T��2Q�W?E=Bo��<SW+�c��/G^,\\%]�K1���$.ToQv�$D��G�H߄��$�ۢv�6�H��+��ź�kp(Ǩ�&n���Õ��YWc��X�&�68��j��4��HH���E�m���#��i���=&��۞o'�Ác/�aZm�g�F-l�6�3�_���#���H�Hm&'��~-�*0"|X�����QBv~S%]#�~� y��;��"�;����6@&��K���ōV�H͆6%�i�U2I�JQ�Z��}܌�xgI�u�r��G8З��~�v'U����#x���DF����Hx����_�J�g��G�𛴺7Q�o(ᡕ�U�	Ϟ�z��������.���	t������g����y4@��������wΑa�D翆�)�B��Z-j{��X�0�0S�	T<�E�H#��D�Q<�����P��5��̠��i���ΐ{p�����IV:s"ft��#�1�m%���3W�����?���3�Q���Q:�@krtʷ�z�������{*�#�򻸦�N��E���	�IJv�^��qF��u�M���[���F?�&]��]`u2��QP.��"��O��Bqk�M����/�c��S��K� ��N)r�Uz� syϜ5��w�O�Z����n$)	����M�+-s~���O^L�	3R~gS���*���+岜��>���bϡ�rvI$��'B����XD�=�q^�{����Z/��c���ژ(�Usd!
���~i��G��zyuo�z'-a��^���&Y6X��[_e�!� p���B:�F��5=�(��\D�n�a	x�;��)���ӽ��N��`�1�5u�W�x�7��T0tB���Q5)ia��IqtHpH�=��޸<Kk��~[̏!�4Ql��JXFvǍ������H���R!y_�cL�s�U�n�^��0��~��Z�Q~��+.�za�?�!�l9��'$o�3��X�.���H[	���V����,�\^�w&?!a7�#,'H�-�d�&���Y:�Az�7��2��U�����u�
����:���OO?`����B��
T�x'����]7D���3Yʗ�iڶ�ɍl!�=���7��9���_D8	��C��A���^�6�d,)y���c!rm��I��F_M9��օ�����������A���<�W�����TQ�^c��QR��>"�CD�6�`~��В�"�lF��ګIJCsi~���v�z
 C���L�'%뙣?넢܄ D�߉�J��MZ"2��ɦ��$���Ǫ��GL�ǹO������{`�gEK�,�FT���vQ��5,P��1F��:۪%~��6�r�p�����d� �P	N7g����x)fO��.����K���G��#!��L�N:���W����Ŋ�*�G�V�R�Y�lci����}��B~�g�ѝ��l��Ő�M�E�Α�ȝ�����E.Ǥ�:Z��@�s_�̘�uv�"r���u9�o�@�Ds��hؗT�e���k鴯�{���b]���=�Ta���鱐���VcOBX���svbj�(�q�0��m-�ċ����\P&-O_����Ӂ����|�4Hq���:ҡ��݌!�7�3���'�� J�pŢ�5�J��5-'�=��s�j�ΕmiZ����Jx����^*����B���<ķ�*x�˰��X;g��dI�U��8>�9���>,Z�~���#�YIԀW�f��-�E�ȏ�w�ĩ|$D����=y�d�b͢���!���8��1P'�sW�!��OEa��a����|�a@܎��`T?�Ѝn�Ê}�O����l{�,U#��D(y�r�m7�t;�4���Lk�	��w�ƗsL΢�����3�:�eZ��4 �>���Q��"n��0TE{����y���Wn���Z�M� ��e�R��!ώ�o�H��^���F �\M��fj�R�u���	�P:J)�3��>�������֦:�b��5��(����6\�J�	�p9f�����	�5v�\�,+\G@3o��A�w�غ6^;*���"�+��i�M��BM�%i�A�CI�_��u������	��UB�.�ā �3�G$���*�$�����{`�庩X�γ/kH���t��?},H{�T{&r�N=��"����#p��5�86��PEa�J��us���0{�A��-����\>E_ܰ�I�tH�?�>A�g	��'��{-��{ʡb���/�Q�iƵ[���S<{����,��q���_�׻���ҙ7��厠�ɨ�k~%�1?����|X�b�>(�C��;s�N��L	�]�I�N�[�=S裓��}�h2���I���i$�<�hs\�BN=�"ڔK)�l_p�MD���h�H�ÿ�탔�I�0j����PW�,E�����Jd֭�"���C�	���ds�X���n��OOV��I�����1r�Z�Y���n�i,�l��ؾ?���O��֎B��o�	�\�fw��9�i�s��l��=%�� '#<2�#r���?T�J,�u
nz;��l��s�ޜ/�A����lf�7r4@Ժ$�*���)^�W��6�H�P��$�G�������5�k
���b~j����� ��g� Ac=���h������f}C�#���{�&���4y�H$2c�&���� �-����=��ǚ*ym�ǭڮ��1@Ȍ1�tF��*���4���l��R�,5�/>��jw��4�j\l�U=��@;}�nc^��J���N��U[sW��	�Iu��ő�����#�*�I�#2��݁�}3�GSh�W�|�e"���?�.�ȵW
g��h�g��5wWq������s�~�O1@�q�'���K�-4�N��g�v��7���)>�@��K]
����G�\B��K<W,(鉀Ɠ�AAM�*�y�R�,�V��4��#�U|Y}�R���f�J���|ͳL���[�hJ�����L7�	?Mzph�ýG�?�m�=�N>%s/�P�2A:�,�IIke�.ӝ?���4y�+kj�4ƚ�_j�����b:x�RSX�*~u.�զ&����I�J�8� 5`���R5���]�Gmn@�P}��_�œ��O�"^���Z7�Կ�\'k����Ί�1�9=(��:*��'�/����m�~��R���a��sM[1�z((�-���<��>G��0�wI���y�jp0�� ��a=��'�08��ZZA�����M:i���A��$�����@�c��p(P�ɝn	��B��g��2�g�~2�?L/Y�B����\�C���#�햨�������MS3�4��7��$iՏ,�����<t���j��P���,<��zߕIW����_���`uP��k�E[)rx�6��������[�׊�a���`(~��uؼ<�6�IP�R_� �,~��썛�oD�a��V���8S�wU��Ό�b�e8ul���9!���Cܑ�ay OY�s��ݹ��U�].$�)( ]!n�ҵoB�<������KsV޻6}�]�S��#a8Ɉ��z�\�P��(�*aK&T���w&�NbFL���h�NM)���J���V�9|H���lQ!� <#�����ƞ�䣓�3tXɞ�A��`����gI���^���CWG�&�M�疸u��ۃ�K
p|R���uX��װc\<�RM��� �!�K#��K6I_����5�&����H���}8I��[4����&ۚ�X�V�^�'9*H�!�S�E;\���Al�K�E��fz3��Џ�z���L�gv&�3��"�����pM�|��r��~�IN�G�#d�
{"h��W �W�U�׈�(.,� �ìJ�J:9E���M���
Y|0��$]S�η���)�;��.��Ô+M��5V�����DφI��ّE�y-n7i-L�(���q��"�o��P��C�x�a�VX`�Z!�u�A�ҁ����r�Jv��f��iDL�����t球�:���Ŋ��4��2m�k�,���ω��6�~����iw{`J�ۀ�|sf�v�k�%���rH��I����(�c�w��h8!P#�|r��:5�SY�p�� ]��C���؅�H�ϝ.�E2�d��#��3�
B���F[cs��+��K�YP�x�w�OK�㖐���ւ͔��U�,K�m��j^nY��a~�]"�d����W�bӿ�����\�&iS���N_��EJ.�t=\K=����L6"��S��r?��oA��ON�h�gY��R�¹ϝ�����U��DҤʜ�;W�������y���e�H�����i=l����s��Y1PkOzW�3,� [���������yu�Tp��*\�T`��YeP�)e�d)�pd��^�;z���V��)�GL�-���J>6��.r嘦:����F��w��|��k�$WMƿ��F��-�U�'�@����i�b���X���"��Tr�з`�[�k�L�Ʃ>��%�k�|��3KEc�PGpJ��ϩ��d7�� �b�4�jH#"�m�k�6�zw t��
R�1&�Mۭj��;�Ziz!�b}��kW�������HY�2�z9-��1	_U<vq�X�[T��tֶ�,��֋�+���ikY����3�¨�)X`A�[+��1Q-��zy�N��]�-�4�:~�C��;J�nM֍l;M��A},�����ͼR-�\��6̇�!�vE�����*l�a1�ϰ�j���~
{I&����$�r �Kd�����bք����t����o'y����=/����$CV!�~C4e,߱�a���5(�7��8Ю0�_d�+��Po{`���Y"��l��Emkj�^}�)�=�n&l�S|(D�>�����z`��Q0��:F2�Ȝ~��U߂�vݱ[�$���FO� ��,���j���8���V�p؋�7�I~H�ϯ�Y��Wn��
�{=�����S�P�.~F_Ԑ�hX>QDbYC��5�R�T�Rہ�����`�����l2=�r�Oo���iPB��ͭ���@��Fz5z�h�gB�"�+��~3tk�N�+���2A�����ط��4/�?Ff����H��+p4,�e�ѵ�����d?�|����Z'{~7|�`}k�4.�8 L�|/㾓/w�%�x}�A�b.f	��̻)��T!�����K����fז䗷��	Lep��a��Q���X��Tl�Y�:Vj��QFd�/�zQ���fDJ�n��P��O��c�?J�6�<E*��x|J�敘J���v���j�s�h��!�
�]�-c�2Vs,[�0J�m���"�1��s��h���&y�����_�+�����o��2�i���!x*��	Hl8:Zɘ��Ϫ�u^[{��J}N��ל��5[�q�ev)����2t�yn�R�޶����4�� Z�	�m�<�������[�Pi�����uOM�.��	I8z�p=�X9�M,���tz��N�K��}�e�ڍ�L#�]|�D���]O��|�.m~h��>�$Q�6w|e�Nt�:�~yS���x��5YQ��Tc؁i��P-k*(�e�ܑ��&��
 n�t�	%�WQf�BX��^��q�[�_^�{%$[�e'��u�W�P�_a��Mث�q/�ή�Ū���cQ	��O�ˠ9�
p�h��9g�Fv[/�����m�n�.�A[�@"�&(�����d�|6�+�?��f|�Z�9�I��֗ܖA�l����
��強K�[�˥=n8�˪	�E�!�4�yu���YVѪJ���25D�'���u�g	d�z�IVm�1�`2��l��!�܈μ��k�K�}��r8.��K�φ�u�:�b��� �>���U�ە�SG����z_�>�}h�2��|@R�������� ~C\��}�x����ԛ�����o�מ��_Ի�Ͳ�a���J𰦣c�_����s����9耋�é��;mG�.;��
��j��	l95�R�6�4}�����ӄK���-��
��Ɵ^Nd��Ǹ0(�WB����O1�}Cl�]p�n"��+�`���-���5���ƴe$ �h2�N�/��}=Y��1��T�ryS#S�2
� ��j`�)rk���OX��􇂎� ��;w��*�e�$�*t�P�s�} ��,�����@���̲��g���T�ز+�b�.�R��G��QW�	�����9�57��g�M,!g`T �l��|�����X��P�t-X�_0ԅ h�T?��n"�"�!����_j�a�-4�����ת�#n���ϲ~�A��q�C4������V4eB�#���7��t]���sȖ'�&8�-�<��$9Ƿ�BH[|@+O+Ag�syB~a/�J,-fc�į����;=�O�^��x4�0��AV*��l[����	��A5~�Y�u���Ҵ�)c"M����l)�I�e���G��$�	J'<���]�8)ee1���3,!Έ�օ?�}���^Ŧ�`W�2�A����w�g����-He�qDa�ÏLt��}��v�~0X�-�PW� �JZ���{'�E�� ��;���W�@�
#�O� 8��H~[B��U�l׶Ч^�%ș�OFz U��;�ա�Mꍜ�Ǫ�%���O�&�6�W8V�u�|��ą�ߧ�7�z�J�XwX}�l�?�r�T���p�ad*80o=�a�8��}!�
:a�5LB�ߑqN-�7L��CUz����F��;�L)O��273aeC/�����WO�/�GC����|0��;O?��D�P_�*k���n5V��aM.�;����vͽ��������u\��} /	�i3+jñlQ]�_��eՓ��*q`��D��*��:/��z!��BF׷���y�7"���b����x͠��T���q��ɕ�I[�}o�6*�{�*f��F'(�տ��2�j�=Z���e��g������WSkN�x�����폣�|�2�f��,����0rE~�*��С��ǯq{� �[�F;��_�:d4����$遠�u{�=$��.�~�,`�I�$�b�Zp����D��b%� ly�,�+Q#�ݴJ�0>F��#��+L�e��=1�vzr��:G�ײ����~�!`3�W�H��%$nL���#b��F��	E��<m�ۏ�e�]���ܐڐ�IP`|��MSP|�e�jwg�� ����j�u�"Д����T4�j� $e�Ӱ�̡i^w�Z�L�È~d��=A=���m(�l���|�cI�%�`%"��~����(�=ɷ��6���tA�S�3���/�1��ߣ����n�a�&�*�f��ש�_���Θ�XG�[ko�k3 �j=��OCi�e.��������B�ޖ��qv����C��ok3��ٱ�>و�̼,�'�y�0�
��t�S\��^���m-��y�l�K���#(�	:g1���/ե���;�ޅ����=�T��vɓ��#��%�����M�v	E�<[5�� �{���j<����6�� �ʺ]���9�J��en�C��6vۋ4ӳ�Q�]i		��B5P�Mt�[�	��想:� /�f�������+[�!?��g���C�E_��z��w~�VE��rWIB��y��j�Rvv��	�|B�a�k-j�	1/#T���Y��ӆr��.���~��hpA_�zEghԴNE�*��e�5z��O�jӐ%�d�>���D������l�ژH�9nR��WU��i�7��m�H��0-/Ui�3��{���*��92�QUF����$�F':m�*����@eķF�{U2V�T�lR��Ҽ=��\��;�ڜ�}��?xi�ΊrX'@oR'6�>A�(L��w�a��O�d�c�n���B�qe�������L�n���'���$|�)��±�W��ґ:+ߞͤ��9�Σ��1:Bb�#��3OR4&${�
<�A=q'�֥TI@|�S؂X�េhT��`+�ma�n �5҉���u���8h��yȿ�N�~����%�YhF�-����	)�V�gF!v����]��E�m�.�_)J�VL���pF��+Q=�/O_�W1�~�8Ί1n��"��;=�29��Iú�iŘ܆��N����I�����;W�͍3W)ގS>�MQW�1$��~֚��'9�'ѕG�c��e>J�jT�O�X�a )����`SaAYuK)�`kFeu��SJX8�/y�Li�_��,�������lM@����1K&�+�=�s+l��9�뇛4,ﻕ�|gZ�&w�ua�}m��7C�C�ӣ5��"��g��b4z�.�t�ņ�L�����|��
%���h��˷�W��Ԅ���u1:	���}W���ye���ح9�m��0|��\&��M�Zq	 &��3���hT�����NC�;�L �H����x��f�z�#o嗧����si�� YEHw�/=���v־{b�ьS+d�e����X�;�È�t�4Ύڡ	܉��K���ct��:X�9H#Z*�wE���˘�e�8��m_t:´Xr��Q�O��EV d;��|2��X���+��<�$r��5/akN䧔��&~i*
Y�]�U�����Q.C�HW*�	5�gҐ�
�KW��ӹW�N�y_�2�d�N�R��tZ�Z��j�B�}�a	.��[�E�IN��E')��t5�ּݐ����D2�5$�����b