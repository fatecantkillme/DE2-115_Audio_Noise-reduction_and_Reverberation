��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<JÕ���<g���S��Y���fߖN�r��1�S��9c�$�aJ�A=˧rOZZ�Qtk7ŏ	zXډG�*��_Y7��l$D:$�	H�-�Ut�X/)��u͛������J:�S�b*Afi��,e{T�)��Uc�]�� =ϹO	M��#�Ҭ�Q9�H�B�-d��/��P�g���76Ӡ��}��c�����b���[dx=]��Ru�o��g��������B�x���b�yh.m��,R����V����MoV��#V��ݬ�-�0���o�����[-ƔvZh{�\��Ei5��kH�Q�y�Q�%��4$�zVGQJղ5��y��xw ��E+�-��j����_t��h�;��Ξ��k�tA&���,\z���V٢�?���/�����̱�"񀻘��C�Z3��.���&�[9jB�e�)G
�O١
k�q��M���Ќ�23Y�B�$�}�W�%�� +d�52���Ź���}���Ԫ��yn��>� |�=O`B�I�pר��I�� )�C��k��%���H�0f�)~��m(�%]��V{���������܁���;�&��[�N��[�u2ga5q���Cd��-���üA�ꁡ6Z͉�{�C��)���K�*Ej���Ld!��s=��l��n�肭������Cp?ʉ
!������<J9�A��l���'�^��D;��>=��G+�r��5e��>����>o$���!̐����+Y58̹)�,�����ƽ5X��xq��x�c[�A�K��G8,��l^	��yj6�]8{e�(�������98���F�����N'���9�^���tW���t�E�O�ֳP�� �W��p)3V`dW�x��J���K��]ߚ)���� ۜ��52�fǌF�t8ƣ4�ۚZ����\u���u����$�o�h�D���f	��C6�v8��􋖷;�(+�@�lg$U�=4��-����^N���3z��g���}zw������n���vwcJ�����5(<4TI��_�8v�Ӏ*e_�.�6o�Y~a=���SӦ���Jk���x+||����^ϣ�e�o�*��@s��W$��֖�������c�Ga��}!Ձ&s�{���j�oZ1n�s��zZ�mŽV�g^Ь���j� 뚌W��ru�l�'��3f.�85�����)9���ϟ��b���_�e��έ
X��1��,I@Pɳp�{���ҙ`-3!���|�:Ar��bELv��t�5jn�Cw[�H�|��Ɇۣ��Ѕ�?�¤@4�����a͕��+��E�y�_�4Ʋ�;b'�}�lT��@.��d!��;���xQ|3��Ȯ�PR���쀽�S;�a}`����J�S?�f1�������3�'�߄1o�����7�*��R�}��3���T_�L ^Q4pa��K�-ɜU	w�+���y�/=�J!��U��B��BѾ�Q�R�-�GggG�d�R�&+kU!U�>M#B��yq��O���ϼ�C�F�C��I��ce4|N}_B�{A�)O�����%h�ٴ���8�!��zp텪xj�%�����#;���i��g�/���C@���i�@z��I�J�A��,jG�n��Rq'��K�F)�"���@7����>C	�`M3��ɑy#�
� z�!B|h�	݋��"Uw�CLF�����0���%2	��6P9��e ��rDB�42�
��z1���-q�����4�Z:I�Z2.ۈ&��T�+N��Çj���`���z^`0=���3a3=>n���=S*�i���t��wǆ4����C�LB��H����w������F���s�D�.Q�w�C���9���mVd���B��9l���
ߺ{�e\-�Z���u�v���5Ay&����ys�i����^�g�50h��D"�lKt��?<��>��@��LF��S�Z�8��!l���}���0�п��gBr]��D���\�6S����|g�~2�,3{`*AnoUN�+[ت��;˫�YRU_M��n�`2a���Bܧ�`)H��!7Ø(�/��P*[h����������VҁP����w�Ў&�s�]Ĕ�����v��SR�d��|��?�ay��_�w�����s���wD��	�>r�3*��r�ϭ��|�%���}��q�H�'�T ��e�ք��,�d��N�zk� !Xû�p�e��@��jA(�g��5 �i���-k�Hӄ6��c�DX�b��3Z���_jo��X/��"��Inn����]>4���)W�*�x�q�`�7���Z�=t�l.@�
K^ �܌��7�IoO�Av$��x��	>���9��Ղ�%�h�ꙵ'�pxصK)�-8�G�#��qTؾ�B_�$���nz���qy�l�C���4��h�C}���$�Q�?��ؓm���M�E��,ȏ�g�
M`�,`k��.�m��{�L�OH6ڨ�n"����� 7i�M�fQi���4��b�nU�y��K��� �P�IQ6.74GAqy�%�R����436�d�� ���c�R�~vos����v���ú<�)^���p�`���W��A�,=_���N=��[��F&;:��]����#���/�Gh�1�M��y0*�vbMfc�XO�_!�l��jw�^�8�K���mݥ��Lh)�%Z�2��{vѾ�ܭ���| ���1��6�ݫ,9�n���!�ɂ��c�-t���g��QKfֶ���0�ai������քo��W
|g�Q�գ�q�$��Pxa��C��6X]��@_�-��3y+y7j�٩و���Wn�W��;��@���Li�߽�X�Ф!B�b�����zw�%��,,XM��8߉xKB�S��?�/��/t�:!$t�q,'�$^��7�ZK���B�j�B���7+��+t}�f��f6k��λЌ�-�DG��x��K����R���5P�%8X��T�Ⱦ2����¯��"\�Z���b�œ��W�6��ܯF'���� 
D'ϰ�8����6�����>���h8J�ʯa!<���u��^u������\�!�ý�����n5�zx��p*� I�H�N2`l)N %��".ɇ���R��fWR@���IQ"{���n��4e����J>AuQ��;t	sHYy��Y%�m�/5MW�<l	��r;vRx0#|k����_W�� B-�fZ���7��$��fTP��yI����^6fdn��^�R=+K�HR�R�P�������m��g���(�QAb�BAe{W
Fhm2��Z��,g����	��S�	KFn���  ^46
����~޿�e��s0�g�'�H`�
d�"���(;O,����#�H�k�`�+�;��LϝQ�.�%�ɤ��aڸ/#��+�Z�Ǳ��3fk:�єwBD�9���qg�D�v�e�Ir�-��n�(�Ґ0�7y1%�m���M�����E��YI6�5���w\
%�2}�µ{��+�x��6��Jne�lG�Bk�㇠�r� ��yQ�4���*)/�5ݙ_�^�Vk��(��w&-��PJ�=�_���Y�E�F.�9�|M
)dX,�(I�g�wCG���!����K<�a��5-n��o3�����b0�vi�"olCq�t���v�K�!�z&N��.���R���T�]c������}��<%<'�͛^���4�v�]��׾�'�^|Ng�KgP�S�O>-��҅��8�k�K���T+k䐡G]���to�C殛��2#�g|��Zg����Y�3��[�_K����W���i�E	S暤P���1�Z\�C,��z��qh�A�tѦ�>���������v��_Y2oШ�Y<�-���i�~����>���,M8�7��Y�(�΍;�������/������"��'P�9���C�0��Ic/L�����f��J��b{E�w��;	q%5�Ci�G��d������㧅��6=�`k���~��~T�;2s�d� U�$D|��2����i
O���nM�v^�}���"&f$B둱��'�Q���N����d����?����B�%[A�ڋ�a��;�k�#�]���~���C�{]�AR��X�=������o�>} ��{T�VD+���:u��M��Κ��wT�n��(�q\ô��#BƖ��g/
����������m��r�걆څ0&{HZGBSH��2�p�L� �U�[z��ykU�-hڂÁh��R%aPn�W�?a�uXȭ��lYc�1Fu8,"���ˠ�Ʊw6U��TL捴��ʐ�[���G�s���/a� ��q����6>�&�g�Da�� �K��Sל26;������0 �0���?�Kp����z�?O���!�AԞQc��( ���1J������/��������&ٚ��iD9�,R���a�����c=�bVy��sA�.�,��JkL�C�3W�,Ȃow��	�>w�Cܦ�ľ�S);�A�V���'vm77�.ѸlQI��i�YC��`�jg�x�Ld��´�YAA��l�������*���S�߂z��G�R�!��6b���g��z Z��`�
�8�mɑ�%�r��e�+�BS'���]A��.� !��E��x�-��Z��0�^�d���"v�b�h?�'f(�A5�:�a[|�4ZX��U�}��.�L����V`�!��������B�_]e�Sl1%������Qs�E��h���k�~&���&f'kY��׭��\����Mڋ�OaI�C�����s���'tĩ^��^��'b�
:ɡ�Ě|���uܡ��x�^�"����Xe�]d.iK`&0����o6Y���|�$�ˊ��^��<�DS�ϔtñ}f��(��8�%���v�Ŵ̍�+K넻9�;#���R�� ��l�S8 �&WCCʅr��D2\���T��竖�����1�O��s6������d{i+�o�i��� w! CH�C�$\D���4>4~��҄^Pa�.ՠN����d�v���/v���鿻OC�,��xb�w_G[�H΄�4�����FO��Elc"r�;y�wq6���1��K�ܒɯF����h��x���VK�:9���NIsK|Ʈ�svv�nR�;�� y���3�.�Z�:�[D�a�o��-HA��g�Ű�쾔)�4�/�@H�M�<��:��,j_�@�?߇rnc޸�F�?7cf���$S�07A����V�d2�����|�O��U8��2����w
���:��5"��l^YJ7L}x���7����b��چ& �91�W�s��1sS��u=U�$�o x���6�3 \�0[��� D����MX=�|����/.|�@��^�q�X�50qo���#�o)���H}^Cd
�;r~�}�8��=x�&fn���ܟ�]�ѹ��M1�_�W�폿W6~��7c�L�䁼!Jރ�����2�����ϟ�U������-��6�)�Q���3Ds�n�Q]₏�rmO�7U�j�QK�\�9c�U�+���(ِ��Wj�̰�<����>��6T4?�I"qt\�g,���`?�
�龟�!��;X�
a,,J�7L{1�;��zҦ/KP��˞���1O����M6i΍g<��1��'�����2#Q@�m��� ��y�y} �������O���W��:&|KQ76�>r超JQB�z6 ���4I������D1�d�e9���@��&�SX��״i`-�36GteN��.�Y8�[���"�v����,w�U�1<c
������ϲ�^>IL���;��-!�)2���B$��%,�0�U�L�p^�8�tS�s��Nfɹ���
��Ba��T�3���T2+�lI�F�n�p�01��*i�=�|�B�{۸�s6տqT�AY��2M�1����Z����&�|���;�5�(�T&�:�I���d>�7��� �/]�ߑT5�f2u���;��	�^c�徏��v�@��'1��_J麈)�v��?NO�������8���O!�L�e�N�m+?~I^��+f�^���zi�;�t��A+�+Xx+�.xD���+Z�w[����
�ކ���U��Z���1�����ףG����/En$�nx�<j`������)׾7�{���J� ]8j�_ �g�:a�6Iʩhd��ߒ>Ҫj��=_�K��p���G/ᚁ'���%���A�3��!	�~���5pŌ<��gbs�����B����X� a��L�����SV�9�/�X��.���+��O�L���l���I�?)���%����CPwX3��!��}�����8I�ݍҁH+�]8p>�=FH��J�y��$�{Bn%�Iw��7���
O�I�#4�*&��|(D�L��7W��υ�͠�y�A[9^#�����+�u�MX ��R�o'��#(���R��:��K�2�5�M�\\}��̰mI�pW��P���n��J��eZ]ƪ��YS�!0z�������zXA���&2���V�M3ҝ�&��"Rh�g��*��o�u�� �a;^���"\KpH�-~��.Ǳ-��� dGA�P6!���;kU@�^yغeR�r�A��l%l�r��������R5� ���ј�)-�>y�Ol���;_��H�Q3�r���0fP���[���Ӻ��::2�~�N��ul���k3 �-cB�@��8�^�[�p@9� 9��}Lkږվo=: 5��PH��q1\��9���7؊ψIw���[�M���R*��&���U���K��1.���r��,s��o'h��yJx8 W�fp�2���);'����So�$�k�A�?����Uʤ���/]�����}ۿ�FbN�i}$z���0I�	7𗛽�W3��y��^�yc]�s�g�&��ƞ�x�?��cg�e�b)
D��|q�v���ʽ,��M�D m��Y���||*{�I��K���$ܸLҵN3 ȃ�U�6���Bq����b�e8e��}���I�~"#����0��D�'� ^��L���鱇;z�Ks4�ެ�v����k@�i}��{�bF0�U��=�� �\}��C�b�������\��(hf��֬��A9��$)����S���+g�.�*�0P�8�R�Ļ�r�K�s^���\S�:X��a�sw�}+���S(�v��((��O�A��b�/��j9���X�R9]¼T�φ�e3mvٍ�:�����9�l
DZ�X�uhI������?�G%�LxN������Yi�O�.��9:3m��v���P!�~��Q�qxb���i��;m݆���NFJ�$����8'�`��:bo�δ\^98��6BflZ�Z7Y )JHw���|z��u=y)����h����wB,��d'÷��S�o��96Z	HQ}^&8�90AP�%/p*���D7��vfб8�h�}`d@s�v��S3-�v�vW�k*��z�z���K��Z����Q�TF�m���R\�����P9��[�Eu� �����5�L�K����n��C�%=�m��5G�����4�D�|���h�d����{^@t�� �-���	��e"��k��S�%8t�k��2m���O�8�X�>�:��s�%���N?>�ą���x�SF��Euz=��2�#XA9�VN�v L�m�;V�����"� �kr̓�xA̞y�/.�O�I�}	s&����оח V1�J^t��r��PD�4F0��N�%̴�,���.�G��ئ���IP#q�Ϭw3��p��K�
��l��9���=?�������C�C���V��&��s���M��t��A}���3�����Y��o�&�+�� G��~��Q��+���2`_�Y�:�*P�@�H��]R�Ux|zC#����%�����%9M�\U�L�˴.��̸�΀w������Yy�;���R�����
!�TM��ɿ\�r|t��|wVҮ�8���ƨ��XE������ `�d��*�>�he���r�!f�T��+��\,T�GK��q���?�L}�@g]/*�����6���s�-X| y�֧4�X_���YW����t;rd��'˖i�|���
b5Yu�Ў��1���i=���7�{�o��/�����F����Z�v����I��D��:b��N��l����,��RĽݫ4�tV^l��]��Ay��R�'��`τ����$��B����D��GCZFe�l�5�O���Q��;��������E�f�U�ϻ镥�<m�J2i���̪a���+`����wO}>t��G�F�h���%�Wp=�J�+�-�@�-)k�;�6�տ�� ��)���d��k��6�2�������Sǯҕ6KE�}����� �����W�v�=���P��O^�(��	Tk$���7���E�Z�$&���sL5�eԝ*M��6�t����o+�Ò��k��Ŗߘđ�is� UÅL���<�WaW8�H��n'�T�:�;T�o!�Dxk\/ǖ��?>�Se��2H����1L}�3 ,�9+�= f�!ۃ��0�5��|���B�~����6�,\A\魿�ڭ�ln���`�=i�V�d���������x�����U$7]#�)��H�dE�,��Oq�SŜ�?%�D��c�=��A�D)
%a�!��1��<�2D���h�zd���w?���\J߰4��՗�f{h��E��u�E�}ib������Ѿ�C���жH
D��]�	�ո"�1R�9j�ǣR�]��BY����73m����p�Q�9[��gw��GȸI�VʡD��;��3��C7S}{�%�J��8�4�rҔ���ֳ�g��Ì�A��t&�s��QoS���=���7YR��tK��q���놳*1�����	[�Ɠ�u�����w��&ۻay��e^ԖYy��m�:,�ڔƩL\6��
�8a���C~����%�=Ix�!)B"���~�|V��]2���+h?D�C�SP-c,��b���%|}���=���-�,��L����/����Z3�8-f�F�O�9��f�pQ��_��%<�B�, �"��`��q��e"-)'�%K��~+�PN^�尷�:嬴)=T	Ⱦ&�H���񮂞���
���3����I�^Xmn�)<��7���X>�QkSX���<R�L�j�Jf�C�pv��i�����1ۨ{�[�K���=s�~�8�Ğ��?��b��#��=vY ������ P(n|��?F\sLG��ͥw�<��~Q/�_ ��X.�r{U[�e.E�g=��V_�f圶Щ7" <���uf��l��.do�K$��%ʜ�+�1@�U<7�K��Y�� �ֲ_Ei�$� �&����KIE�c]ٟ��sS4�>�r�ˉ������I[#|�W���\ ����uq�Zy,+��~A�hm�4c�����I��Q�j��DC�3HN�JH�ϲ�̪��oY[��"�T ��(}d1�DP��Kc�����u����h���$l�ŕz��HPЏ����L\�Y�7g��&�g���w%1�W��~�2�f�? ��Ўx�-"v������Sѽ����\�i�@}g�v�Q����֝�^i2&�i�J�Pҧ���ҩ4u��	�%��V�F�V�������48ρ��S@� ء�/tsT��R�^�Y�6���z����(\��������.�[�^[W:v;eP�+e��v�kH��7ǯe�>M���&4YU�D��-\�E�86���J$�:K���L�jM"ɚ���p}�L�a�^����L��-�(�A:��l��  wuzq�årjӵwhN��@�۱�Fr�ƫ!��5Y)�k��2�}�����F���eH��U�~�9<�f7"6��xw%B�+�ѝY��߂=���x�* �� ^�Nj��v��]ف�<������S8buy����&W��D^W���]��>7-��dl*�}�'�l�#~4k_h��M3�;}Li���Xj�R�wTB��leJ�@�ۭ�bjC(7xcRs���a���,x"�@����*{r��fG
Ў ���a��� ���xr�t��}��v�O1P���aȌ��C��e�����,���O��vz"B�Ӗ�`�=�E����\��%�)&Q�&��cBy�(�N��'��,6�KF^���rçF����g;tZ��l�����t>�/ b�_��1�1o0=37p.��o��F�������s��ܕ�ɡ��&Q��S��:�ne��h$u���UMe7M�0,�[�Sm����]�?�������f�W�n1�W�(J�â*�=˶�VQc�� ?���1�v���k�ܑKUS�FR͓����1[��,��X�̤�`<����P���@Nsv�j
r�1j_K	��m����p���t����I�%@q�G���J�2���^n>+�3 aq�{%fR{����R�;�;*ͪ	�{癜�����/R����ҽ���E���CAU�ְV�f7�U�*g���T��6a��	k�ٲ�XZ(>8r���-A?b�����v)� �j˒�%�U��ի�E��Ǹ�>g A�^7%W��ڏ���L��S!C9�o�� �T�Y���B<��4 r��'��XT/	��w�e5ϣL#�	_�g4aK<�R���4���z8��\��yv���ׄ�i9yl��#�t�Z�#��ҍmOvRO ��1��i��t{���"�_E��m�-�ȈY�J��#�����Ͻ�t����p��W}z�(U����G��.%���sI�����m��D��r[m� *}m���$����� �����S��N4JU��x�7�{t�q�:�j��j�{�h#�si���^�^|(�O
۪�܅����=���} BOqf;�j�� �5������{1O�����#�����Ts4<�\�w��$kΞ�j�u�t���**1���V'H��OC=�z�r(%�����>cdv�UŜ#-�'|slh�u T�^�i<+���"]9I�p�1����j�t�^��^l�*`A;j�)��e ��M��.�2]��	o"���rv��W�5=?���%G���D����K~���7��B������K��v��3Dwn��-�E�� ��|-�(4�X��X���	���u#\�"�w�L���n��h���P̻F�@���1���N(���K+<�����뛁w�q ���]���]��رa8���a��<$���p��n�5˹~����7W�((A��4A+�Y�dUf˿\�ߡ�"��o�_�
�I�ҍ�3z��Cѣo���ACU:�Z<��&@Hq��~�V���"��ZE����Z�=�t%?�'��ٴrw�
��{eF�6�v@qR����2���-�8m�����Ĝnm���9(f���Q1� j�rҢh3&���ٝO����DS_��� ��7�˅ǚ9��\�W���E%��W��g�[p�clەd2�S� �-��s��?�M�.�|E�6���j�$Ⱦ��V1������������5�ê��.<2{h��	;{���̐
F2a���9!�ll�;)c&�,C%F��B�_�:��Q�u��^	:^@��6��J�aᙽew��L��vN�T���O9B������M&?�Y�&E' ~�����p�� ��&e�"u��eJPF���`�ú$ˋ����l�!�*)���#�`�^��>8�}(U����N)�a��5m����k�Ɉ� �Ą�����PhN��������dV]��a~�]���*/h~؞-Y�#zk�����\(�H���;��M*c~��vw~aW��5�J4י��м�}��D����Dt��B:��9��f�3o���<��+�3 �I�W4��ܣ�����H�֑NO�#/�R'��|�����S���.e��U����F�E�<������C��$��v��]��e�$9Sb�c�敾\����a��ÄP�:l _`A��ג�|����k���*��)��.��T~��TJO��`�O���c15��/�K�-��O�-��������+��v�P	2a�M��Y��� n�����鼰�-�ץ�A;bG ���/2����R WI,�K���I@�*���uOi�����a�d\i�:��\������	u;��>��'-�9�V!�P�B��ꁤ�r��+:��]��D�x�ٷA/q���u	��i����g����P�!�f�TӁ�%əN�*�Ѻ�[�������B�g�7���g{�}�ugy�+T�z�(]c����T4�`�|:6�mw��Ut$�V��Ĝ�F�g��}
,�߻���u�Q^[��"�%^b��w�l�m����_i�����7M��F���'1jv��Wj�q�R��bT��M1oQ1bo#��V�ǜ�հ� �lG>q[$Vݘo8@�U��wg����1�N�{X�6�F"Y����}���q��a����X��Ĵ �{4ghG�F<C���z�n�� �N�gR�!n<6;�py`Xg\�P�X���A�`��v-v����n�&�:��ͼI���?~Y�(v�f�e�
^^_'�(��~�Vð�S��(4w����'z�߆mCww����\��ȏ�it��7�Av��6�����5G�5K���(�ʜ4�sx�,Q��k;���a{����O�n������o$�����H��zl��"o��6-]�d��rO�v���Kx�B� �9+=���E���|)Bٺ��7X�V�^ͻ��JkSZ������u�5�):�yf��7rO����\�����A@t�0!Ab�M�Pv4Ʃ־�n��|������@�(G�3��P�<���c����!��u�9�3����y��t]�r�=
�<[����r���L`�@5�8��j<�5��	��߸{_RXV`�Y�-AR��0�����Y�~0�j}��#�UƱa�˶�y;�^wEBG�{���ܯb�B��I�X���c�j1% w�S3��Ŏ��U}�J*TX��F��*m��d�i��4~
�����iU{��2�zԄW�7�)��ON^|���\Hb�U�����E\��1��UP�׃�X�O˷Δ(�R3��@&U��4x5)���_zqђ���X�˛�1��}�(�,�eD�N�kK���c��}�����{�[}�Wu'�l�@��Z_6o.��>E��8�w�_e�4�1�5Mr-&T��e��uh:^C�p��2���4H�h�r���lW�)�Q�d|�Ia���^t��+!wyRh��S�J�+!�e%�&�Qa�	=;9?ƾb/��x�@ӫ�e�0�������]��{W��k�.�c�>�B�;�3�p6�
�]B}� �ĩ�<���r�$�� �?in�H
 y���_jx,f�7�%C\����҅���o��[aNRd(�_�ϛ��H7�M#�k^�+�&�����
�T����3)�X<���>�`��E�ë���0$�W�Q�6K������/�������h������ *��V�&��n��1`������/��R�/�?bB ���I�}�c� �H&Q]�wTk��US%ν�	�D�g%����uf�xc�b!���r;L<ir�BjEBJ&�ߌY-[�-	��:ӕx0I���E�ܿ�N&�,)L�*?�gD��`J��	M��+�֊i�6����5΂�cҒB&X9B��(@�<�j���D��r�BUq��f@��������k�-���\�C{���rd��Ǿ����Wv'�S7��H�N.k'�yq@
���|[*yL�ݑg�+ze���M�r�;��z+��v�w�/���w*�2\@��FG|�������w��W�/�M�C����,��(Ӆ��,��,�bJ��Y����K�!Q%*���K$j�)�`D���}ێ�VNlBlX��_��%aN�N����*�]����s�D6c�gQ�����|դ��V��h�-IUIPUz�e\��Y��P��:ԇ!~�l�:X�T�����s3K�����Z���6�f�Ic��8��Ԙ1��O@"Ɨq�]ד��ܘ?�ڃs T�a��䍸��X\�:-TA�^�e�V���׀"���U�P�qPV1k�Y�2��ό�,�5�u�z�����a�|�'s��˟��Ix'.��|���D�V6��6�n�Dz[��gk�*u�>�����O%8[���B'����C�g�ɘ��Ɠ2�[?1�ZF�	T�(�h�߹il���'"�K�L"�qb�� �lfQ.�Į'AJt!)�R�@/[7�3�>��L�O�t���>��'��FҺB�
��H�ԙ���֭��-�l܄TX����6N ��l�&
�w���\?
#0�`nD�V�Έy��oe����'eb���V���E+�K��
�C�N�2+Vg�M�A��߮��\�O!%�+�n�,���U�Z����|Hj&b�5�G�X{��q��HS ��'"[d��x`��c:LZ�Nc/��s6�Zi�;$�w����_Y��o��tas3�,�$�&���G���#0�Y�y�m&+�8��]���z��m�<W:6~)��A�r��e�Vu�@[!2�����3ENzR��ɘ���a)�_�oڦ��H\>�a�
RF���;G{���~m"{�b��.�=�E{���
�ə+��K�v�e�uJ&Ke-H��~�Ĝ��j�DB#�?�K��u.�3��M9XնH�;JŁ�Sg~a��q��z��n)�8s�$ ٪f=
��dͲ1^P!�*>���,#���U,(������xsr� q¾�,��!͖< ��7>3��h�Il�L��pD�m^ڌ�m��X� �|��T9N�-�֑�j�&]�>�8A�O�����`� ��_��^�@V�I/ ��[D�j>T��M��W:;'I��l�;ʛ�(R���O"T�����Éw͌KK�h���M���s�,`��?:�@�o�q#���dn'p�ҡ�[a����������tLj�N3�>?�[��t����Y�SaZ\��������S1�0�'~��6HA�{`�#���
|�^��g'WyCO�W.��E-�0���Ȝ7��,<e��X]����?�7�tY� ��vf�(����&�PK�o�+yV?�@p�xq���b7���UG�]K�d�eٛ{��.�����[�Ԗ��!\g�Y���1B�9:1�ah9�Pv����]0ʁ���Ɩ�Ip��L��ӌ^O4����� ���A�'F�xN)�_'ɶ�0_��<SS�)�f��%��Z��S�4t����o�
�����|'\��r㠼㲤3��Z�_�rr�X���Q�%�U��'t%"����L�.��u�ۨ`	���dY]N�c��#R����G[J�=���bq���jju����:�I�G���M����_h��Z�e�!��&+
Lm�?�J�Tޱ��bAOu\B�4�qo�I.r���9��W%��k�� ����YR:!�_C+�����>��F0�-� ��R]����G+�Ҡ\p�w��G��K��L��kW�Ң}�3�_-�pj��%�B9�fݧ2��9�>b��X�F��b��e�9�g���(���W%"�`����b�W/zE]wmZ ������E�[J��y��,�wŁUG��K%�~�Ʌ�>��Y��wq�%ư��<J���Ġ^�~o�ro��۫H̓����.d�9=[�yR]�Wǧ�R��	^�Wˁ���TڧԱ���
�g�g��'g��Ǐ�K[𹿶��L����2/~� ���x�M΂��̀o����@��?�z��a� B�x{~���h2�web�V	��q�"v�Ǯy�.F2��p8��:��@Z��DyȌ�6x*F��
4�;��N�}�\�������ޫ�:����[�ǂ�%�=�������M����@�-̶�\`3�pJ�b΋�2�{q � 8����`�,~w�	�]��c&�ub���~M3��j�����HcH��&)9A<�D~�9d�b ��)�3�"�9����X9u�n�b
�c/�0?�Jxs�u�ꫫ{y%!�2<�x��ϳ5'��ŭgzfm��T�s�X���؉Z�H��AI���W��P%+fZS
�-��wŖV�)M�7�~�x����\�Q9�F��t܅W���Z�!�d�ŬV�tc�T���'����K�Y�oP��nH�w �lE�a��D ���;PB�g�d�rd�>�K_��26�=�r�}Y\���^RX�!N���L��Y������}E<�]��;]B�ջ�6�jK�$Ώ��0� �����,�@s:b/?�#t���O��E��L�x{�	�*}�IԖ�p�<�k|����%�v�u�(�U=+0�h��!=�B�>f��D{��o,�i�[���`?��/n��TCl��Cb잉7CN�y,4�~BC#���hl�+h6�����?Q��������2�� ���Y������=���-l>_O-���]�ᦩr��O͗/��}�*x�,�i�U�h�C��,�Mt2�7�]+��]�T�A��Y��8�{r�����#�]���Qq���^��,���$���V�%������$0�}桄�<D5�⊐>X�wf�:0ɝO˴d���W �凈T��7bZ��/|�����o�w.��3�eN]$�rxAV�b0�����;�t��@Q����%@y�pm�IFaǭ|�����;z20�엗���d���uRW�O���nA/u,�K"@��&fD�L�8�������{��EHD2+���A�f��b��g>Pz}�JE|U��%6J|KS���s^�vj@f�Z)�}���>��ֆ���X�
q�)�������c����	��'8���	V�4׶�Q6n�ߧ?�d�Z�����Z��v�G$Nm�r�ԦH��UB?@O�v>;� ��i�b\��9��nl��@�vUI�z�V.Ώ�\,Τ�e�����*&�o����ib�l�CCu��l�#�U���;e��У�p�&�ȕ��e)zP�?b�6�rݙl�3���B�V�)��D�E�˃f$�כ'��P�l�U��P[�[��a�d�lW�*@�-58��	���d�8Z��̃Tߺ�"��Uc��g��-�k���5ҝ��^�\���N�F`����3/Qd��0�,��	̨	�sMr	���t�;^��V�/w�X܍�RM��)-�=�Ci,��j��і3�#a98����]��G���A�n����?�8� �1�P���Q%�7-���DH�;(�� Z����Ru�^�L4yuZ�6������� �䂱s�!ɿjR��o,���D>
�_�Dg�籫��ZI��Pb�ܷ
Jk>�Ҷ:7*��xiS��(+�cG2�u@��2m���EA���ap����;ߘ��c]xVb��5)E���� v�a��?c@3/n5 ������=�CK�{�{�	e���P��Ӱ���*,gl��c��op�y:.n����;eA�F'ە�V�uN��s;��mj�j���q=d^�(�.k�a��WS�����?@��1J�� ��t����z/������

�i!��G��c���맙z ,�k��M����ʹo�K�z��p�/�|��p'�xYq���|kY�M���<}��d��w^��Z`m	�D�+i��^�@=~��t3ycH�SG��o'u� �-�6U>�3��E����U]�A�K�r�%�-��d?P�e����<������;k���4���������ZR�JU��Y�1A�4�8�Pq��.~k��~��V}4���|v5e��oPe)	<ɉ^(�*!7w���+6a��^ŔtW��m�?��L^�t����湝��,�\������L����l����M��jFY��>�(i�	;�X����uoL�[����5;�A_�zM����_���%�x�t�R���A�oC����nЊb~�C&��gu�w40����X���H�*su�vZ8�8���&+%��B�W�F!�7 �fC��*�NFP��D�6Ї�H�ő�.ۻme�A�<�>����Р�BF�32
̚�`lo�;|H��8�F�H� Bڇ����HeZ���/��׋y@�I*UZ]��%��)�M�����`��� ��_Z8"��Wn�f�<-T�y�u~I��b���)��5�J��"��yK���k�ӷ(2���%<o��*~{Ό�`��A�`S�j�M��3��ЕU��hy��O��|�ؘ�kN�6�7Hח�ھ�t�J�+����F�}�aMKS��B&�r���?i���r:�������-V>��/�����P~�n�u{�0.�X��k�����H�U7=]��Ն�Ď*g+	�Gԥ�՟W�}�ݨW�ֶ�rcK�&��6�,�&��M��D�l��*��NR�\�{����P�N�S�P���p1�-H3M$�K_�d�y��-{�RV�nC��Q^�%Ԡ1�9n۲���='����� ���XVl�T�A/�uA<1�H|���*)ڵA���'�0�WҎ�ɭP�M� 5�O��J�� �O�^�xb����K��؝;-\�^Ss�4�{�*��S�R�wL}�Mx N���W,g 2�5���vk�����#x0�&	7,�v�kJ���m�x�RI�I���=Ժ�����夝�ғE��e-�}Pw�%3��8�H*fۧ��\A-��Ǉ��~d�����ҩu��.��T}�z�I�>6��*�V!��*k�Ζ�J5�=� 9}5��e-�������;�֞B��H��g0|~�W�.��.�E��h���c����G3���?�	I<A������#�^䊖N��L�)���7ь��I��[�Co�'�5�b����0�-o�	��=I�$!^���-��D� ը\�-��	*�Y�+��K��x��*n�����	�
�.ӻZ4;�k�������{]ՈA����W�r���7�?5�1I���^1�'�*�H���g�t�\ ~���X�^g@���1C��:ڏ�8WR�� d�{d��zP��x�g��hY�����)��)��i������l͠���گ+��g��o�a#�g��@�PN��M�̧)�J�v�B0n���Z錏۰�n&���KU���n�~�Ļc��oe~�Y�͗���U�WBn�8�*�;������.�t�>���]�k�bN�!�c��4�a�-���jW�ٺ����BD�1�e-����G�֝,t<��$�v���\0��3���]{�UQ@���
/�N�s��,�K���H��wAGH�Y�������Q�3�G��s���IU�/�U�P�OG��I��fu1^�$�:�w�gȖl,�H���2Ճ�߄9���c�:'+İ�����>�>�d�&���=q��b$����c��Gv5������z3<@C�Z��NLL7D���'����d@v���d�|/օĊ�4}��q�n�����,�oF%��hИZ[�L$٥߉$����D��ċn�v�U�~�U�D)����j��
�6�;���3e>���Z�0���F�����e�D��w�7�`�	��4��b-���S�	w�LyM��T��׿�{P��)ןg�/��P���٫d �=Q�\��'[@��ħ�����W��v��[ �nt�X��p1����L���D��9��Ҟ�e�Y,��,x�*|��
m'C��AB D���\,�A�'��*?. �D_smB) ����h��%�E��V�����q�2�����F�oq��J�ڵP���5�\���D�stg���0��]y?H��(툊y3(x�qUxߖ��h�i�DI�D�3��Ｋ��0y�cȴ��a9�<��E-XE����-F�|�f~FXTT�����0�y��J'�6��ƨhTߣ�S�����C;c�VN�'&x�-�l��5vϗ97z��Mb�V֘}���	3������ެ�^��4� 7�J7oD[f4�yc��:W7�{r!�L^���9a!�Pv�4�v�u�\.]R���u�6�]�L��Zzs�4*�襰x�v��r	-�Q]�.o���t~�1�9>ְ�A��%��#I2���W����T�-9`�6��C�R8�r0s�Hݹ�G�s�	~_d��B�9���P�e�H.w�!�l�M��W��ٕ�9��T������Fy���ڕ���S�.�J�+����<��D��`���q��1���7��;X�mI^J?@7�I5�^�>� Gy�P����_p�ofM}dG�O8p��M�������)u�P/ܭ�ᗙ.��r�6�1�T�h�8�Q�#���]N�{��P�W��V�Ǵx�ȡ�, �̿D[�k��L:d���g��m�����?���k�-n�ܨ�� 	���=�Wc��0���aaq��
�$�M�&��Y,���V�S$��_�J�|�.���FA}��O>|&�GI�*����/�9�?w��ا��������J��r��zJ:���@&�)017�G6��Ƽ���9�/>����m���r<��qć7f���(>�r����bHs��5a��0	xi�(w�T�#_쟁�H�(HG}��e�2���R�zj��$I_��n��Ύ]S���g�#��+m$.����np�:�ܲ���P}ظ��;EF�c�,ds'>ڦ���,����u��+Sؤ2b�lg�z�*c
v�5�<Ƥ��(�?^F-A^ǆ��=7Q$�P+���[��ϸRr>.0��ER�:?7�~:�!��E�/r�D]�����ԭ���=�=�}�h�Q]3�?�
qu�'���5H��0��ȭ�&9JDT���|��Ȧf�	�����A��B�x��2�l�~*�������t�>�S�9}n��C�/����n�1�$��X�4������K1^�J�v�ɔ|�m�V�1s�br��6�J��7��7�dV�xL'w|�V�F�-��y�C�����*�_'9����+�]��Oh-ds�	*w]Z`��:4�7�kg2j�z,+�fΔ5��>@��ݵ<yc��$��=,m��+簝Z��؋F��� ~��UV>��g�S����ܭ��^瞪���$��0�d��26������8=!���=���d�g�z�,�>:����:8�*{YW���4��d켗���Y����
	[�C��L�H �R�J������]N���,�%k��PA����RVl����B��	�#n�b�_��w���Z�Y��є,A���9��4ko�����~s:����x�G"����Ö�Ɍ"L+cv �2�/~�v)���8i�2�H���G�����`-q���;� ��S��_x�-�FX
�+�|ctJR��w>(X�e2CLcL�ľ�1�.��k�,<�X�{���������U=}j�_��4������m���Q����<�V�|�I���	x��NP�I���'�9N��`h�o1�8�������Rf������p�� ��F�ܽ�K����n����S3K}�d�ey�?A2����'�T'��dR�t��j�Glݻ��:���b���u-z����m��!��ÔE'+*��]�����-�	�,>��?��s�Q�H�a◴���x.[�
rۻ�}Vo��QN�ΖԂw�$�'��^�s�h(u�d�Y�2G�h�;w��`��� c�E|��%��gsnYeD�bx����\[g1�� ��	|��V�L�Z���d#������A����P�X�hxI���N������'[�ᒒ
�o����Vpg�w^�!�Ąvd߮����%��"m{���Ӓ`W�W���X��ɧ.86�Z���Pq�#��3�DT+Q�����`q����	.#-�-�'�ĭ�i4sP	 >�
m�$=�UܮɎ�}`�nv���F�@�a�٭�.T���5R�7X`ݷн�1i�=V5AQ#��+^��O4^�--�Y���X��_<�Y��1$q��[y�ofV�6b�~���Ʊg�L*1�E�}�q�
���9z����5ʴ�kbL6����$$�u�ʕ��y��P�	:'��3\q��G��-p�ɶ�{hdw��/��Z�qOR�j�`W؆Ỳ���e��=8�h}��
K��V��B�Ə�D���׬�A��H�Ò�Hɏv7�H:P���g��I��pr���5��ytB�-)�R�j���Cj>W�3�o�p���)�ut��u���lϟR:>����!8qG�O8悍!p"ɵ��ܣ��D��8����][�0`x|0�d��3�?�3J�|���H��]����_2����`f��e��4W.�/9-uQ�cW緤���s��A��M��0&�4����\'��i��g���nT�F���3H�Nj@3t��^/A�3(W��EѾ=GU󁘏j(�A��}��"Tw�ta�J���)[�����o��7XV��J^J�4Z&H�y���y�ux�_i�Cg�aa�&����W���Ž��\hp�b3�AcU��!5bM�:�ML[��T�7�vy�D+���Ǩ�V�2�2���D�Jc�ϛ���#���Y�i���H翬��(��1K��vf%����������l"X�^q��L5�k�'����{�QT��x�$�*{�3�W��I%����u�&���he���N�x��E�zo#��m�+T}�ۇRh9l_�w�x���?��;_�ɬ��fdl8:s�?���_=�`V}ͥ����=�`WZOs�0�o�
W&�VR϶ԊXL$�fFjԙ����(�pSU�A�iju2��[�����,��8��^�W���`���5���=C��N�B=��v���>q�%QL�T%>W�����5�>f�/fD�M/>&8�����ݿy
�h��IP&��,T=��/�нT �������X��܆Y4:��.+�~t����J�&Gqz�T�2����C�P�)�֘N�{>���C�d��+���NT����_�i)�^DN�}4�$�r��y�-ΠI�Ņ��G���I������o� 九��j�����np��"
�P�e5�t��T	|4xw��8B8�Ee�N��@O���5#��m���TNW�d�!�O�l��ɼ�k�#%��`�q�� �h���y����v����hݼ�=�ʣ�sD9D����_���i�&��Ef?��U��H�Di�|)��M���/C�,3�Q�w�6��vF%n��$�د����M�ZM���! ��F�{7�u3��kO�Vso��ލ
a���d-��Ͻv�Ւ!ƈ�wc����ԍ�Y,wyv�Q�Aǈo,�+�6B�<���n�Ƥ��hT�ơhg�Ƕ�4Y�^݋9�)��Ƅ���ϭ�{~���TY��L��F���@ۛH'����y�����F�râ���6���/�q�$Ά�%��6ּ54#���`!�y69�v����3���;�\;�s5�
�L��%�����0#p4��':�����EQ��}�ԝ�`�z��U��r�nN�,ȻyYt�{{X���{J�x�\6ɷ����\�e@��,{�q�yKX�]�C�W��O)��%�ߴ��A�x�������: ��X>Sù �*u0vQTʕ���j�䜲B6�FB���f]P�;�A�z�*�$0��*�Ku�^n��e]\8]�FDf�➵��7��/復��=��a�JMm�<|��J�qpQba�I��x�?�&�QS�i��d�{�  &�H���G�1�	�7b	W��2�o���U�����N���W�A�2s�vl��ہ��@BQa�b%��D�|�l~E^z#N���~[.�:os>�7�����C�~յD7�a�|�p$l2��_�k�^�s�/�ْVd:�q��]�ϻ
q��qr���~S�m�vz6�Go�w)-���n��=t����#�U���K�"Qe��yE})�r��������=%��#9y�#f9�����y��x�{�U��<��+��&��`�C�h-�譡�Ҁ0z��^̽�j8K*_�XBq܉D9ʒ��N����w??�B�w�������ׂ뱿���[[����GPV���t���/ĉ�a���8 o| �i��gf��Z���g�I1Ak�Zh��E�׋�.�v�n�zWˤ!s����C������x�Le7�,S�K��GY����`�����t�t�9�����]1���ӊzcK���v��p��K��x���]�ۤa��g�hs��ܢA�5��T�Y��K5#�� ǝc�d��.
sQ���9����`O���6�Qi({�Mf-���2]��.���� ��k��4��EXn^���.������Zۈ.`\]��K̯�HD���e��_C=�p�I�8������a���*m����Ku�y��t�}��Zp�m�� ����	���4�B���(i�6>u,:Ig�}}��[��@���k[��jwd�"WB�������X.k
g�_.�k
�K'����G��ռM�˷c\�j�ÁcA�4�|����ba��ٸ��GH��0qi ?���^�M��r�L��b�6�P�u���<d�gضt�C&P������������#�m�<��KFWg|?�����C�O`T��-�_��;�Y���#��+@L%�=Ò��� ��n±F����|��*J�Fo��G�)^�ǉYE��R�D��G�����9��@�5�����13�c���,I��_�U�
��č��\�:^7��g�s	�V�Y{��#y��2 ެ��/5�*?t�d�_����������1�-i1L�L b���k<eU:7�h�W��Ol*ƪ8�*���#cB�H٨*UZ*D,�5&�\�;')�`獀�	O��W��Ǥ��L|��
��V�b�"3Y����b��n��gZ���ǟ��78]��#��~3��m�����є}��mYS��? \����:�����3{�����Y��uM�����?��k�qz��ŕ��g���(�؟5��a]wy�4v<�**ٳ;G��4#,�w@�JZS?%��/%��{���p�oA��B�c8���(�84q��ߜ9�Wv�N���H�ր�������:��+��L
H��J˿s�7(��u���_���~�bíәl��}3��=-�o�j���E"a�3�ܣ��ό��M�'
�D;��T��
B�,�������S�N%ۜ�q��F��@�?[>QHv٢�Ե1���U�HPĀC�&'L����V�<��.��2��|ӷT)�;��t��&�n&؄XA�C�E2�]!8�����^��@6F�
H�(.�J�i�D�N�N|S����U��c�H��|6�#��#K�6-�+�)�9��:�t?m��g)�"X��4O~�j�ʳH8ø�?�X���hec���,�,�(ot��!=+�%Է��8ءT������L��!Ӓd���!x����1Xl%�Έ"�5E[�#y"��vb�L�|�{2�S��Jķh����Um�Yq�6�g{;��jǑ����w\��J?\X�f��Fe5�x@R�W����C������ ��&� ���	��
P^:�d�� �Z-7�'&r;*'IO-"��/#������?�c���/�&ే�(9绎	�4�YC�W�~Oe1�7N�����?M�q2�,�)��Q��Y��`BUl��]��[
��(K��H�]�_` �+��2���)?�?�or?&p�h���wC��@���'?*�}HԖ P��ʥIu]y�;���N&�<�n�8�8g��]EF9Qcܪ*��b
Q�f�K�cc�Տ������e �����lz�|`3�Q#:1�rR�1v���u���S��}�Q-K�	�N�M-K�^G		�ڴ��L�N��׉�4+d�>}�c��y�D&�ʷ�%:%UiD�+�M���#�Dh�H��)��Έ۲�N�E�a5g�6.��+�+��k�D���w֊e=97�2�<$5Y�;5ȏ��ZM�8�ֱL�c�3$#u���rn��E!o=i��/���`*l���^ܼ�4�3��KM��gEd�cVs?^hUܼ��� d���@%��,�w�jf��q� 8�4ȑZ����6�}�|����A�an��e���b���=�4��{��1�:������U�^h:���mQ�x�}����]�K���q���{H+%�fve��.�8,����:H+�}��D��G����h:�.����5��;6rT��0y)����m�S3�'��l�� �l#FH��DQbOF�4�>��U��\�#��p���#2Dc������1�}��{jY���t�麶�\.}V�;վ��^3���^i���I�g�eH���	G�tɭ�C�'`Kzw��_�[͜�1��{���
4��)|y�ܗ�ߤ��b���R01�i\����5�W��d&Qߐ|h5x�(8���f��h�����5m]��pj���A>:�	eS�pl�ZeUq��A����V���D�D���~=����#4��|�Ź�l!;4̠��RWS��M	J��i��OG>���0�b���/\ �1��9�@��L�]�A�e3'�sg⁒�v�D�􌑙 RV����fڐkyF��h��B�n���SzA��e�Gv���W�jz|g����V�`ġ��ϰ�k-��� F�#g�ZҼ�d����>b���+*�'��3���fM�=���R;���L9φh�`�e��Md0Sx;L [�\G���D����I�6�e�RU$��C�~]���R?	!��'z���5#�k�?[�`�`�T|0��]@�d�0�^��G�k�V�:)C�S��s�����J��؟y��}j����(\��Qg��2���~���蔯r�7�'�jT��l�.����O�z�1ٟǭ}��	S����Ij�[��H�m��s�n#pxp��ī�Ē��nQ��u�$tvNku�>7d�N�3US6��jEN�.=����b���e��`HޗY}WC	4���t��6;V���/E�NU97|�{j2��i��Hu��_c>8�n��g!�g�����z�=�i����.�����;`�d����FBcĸ�2F��,��aw�V���׫R����:���˫9e����2��~.��6�y3n�r���L�X���D^Ie�]�аu:8 ��G�q
��6��B��<к�Y�1躈2��[Ͱ!
�-��v&7�7"�i3�3�L$��YOU2q%�o�Rxu	�{Lv�eQ��w{7�����ݓ.�VL���e�<���2��	%��y�X��������z�p4��x�yE�q�?����Rd�YgX�E9��4�1�1��Y�m����R��t����B���y�U��s�A�K���%U�9	!�����c ���=��Ky��y�V$O�b���
��8�,��j�x;�&[_z��V�O~�-���I]�wr�Vi��#qq�c6x�w9�Ҿ3�`B|��g�I%1n�
aηÒ�ִ,"�"I�� �[��}��=���w`�!��c��(.��Y�$7�|[t�A{��W�q?��ACf��b�� �"jк9��$��p�������V>{K�6���pA��nɽW�<L#���U���Nh
�Bo���u*���4!�xY���@-tpk�$a��������:o�����T���< ��J�Ǉ&9��w��1���Q���x��Y,c�+�l_`qZ�i�Șb�]{����`R$��,�L�`�/��#���3�T'g�hx�&	V�v��&-_B{�M�����S������.�1Õ���A�[�)!Y��8��ʷB��+������*	���$ '�2�����cd/�����Ҙ�����qV�,uQ�ֻ;� �]��38��`�̸��%�'Z��8�¥PF�t��.��`��y������9��ݦha�\��n��5��G����{��/	l8}˅q��<+لs	��\�>��%]����:��УԂr>���6�ȢH�����?(�K�3��a+�ڠ�)_�s���z�S���ی�hD�}"�K�A	D��r[Ȩ�"�D�|>�k��%�Ǐ�1�ܫ��#)š���f�	X���Ls7����$_�}�V�+�6}q/���?�2e�ο�	k0+X�цo؎�;��M�ё�}eK��J�Ć#�8S��:-�d��f�H����-J��\^��HR�ꮒ47�Q��Ty�ʏe���<#$d�Ì��u0��d*ԡlR��������c��Q)�MYr���~����1\KO��vzTo>�۪�J�MC�p�R��=����vV���l�%��[!��M�a�E��l����	)~�jk�A����\�c�{�mw'��T�xr����f�?*��_�|����4uL4d��2.G+�=}�ؒ��������7��Ά��Z4���Ӏ��\Nc��&؄�Igy�%�В�ZŲ̅���.K���b���;Θ��0�}�'v��Y]��M��t������<�-�JW�'z	���N�}WB�0V �4��L�x��7!栱����QL��ߣ?1�o:����P��缾؋�ي�r�`Jd�?�����E6=�ŷ[��(fl�R({��[v-.?�/�4ReR���L��K�!�M���?�u)߳��k��j��h���!:_��8�ܪyN)�ȋ��<i�Y+�s�ъ��j�]EݭNK��(b|�&��s��K���:z�5��[!�)5��������-P���)��U2D@���rfz�����b.����UT��~����b(�
�<��=9�ykx4w)M��q� ��*k_Ƽ��׺���e�253x�^�>����y|����8��û�~�zk����Q����x�x|���KD�(�[�ͧ���-c�e��-��`�㲽� �{�v9��e�HRU�W�{�پ�u�#��I�s�7�Rt�Q�����L����00�������f�KCi�h�e�;;n�1����|(�e���jL`B"h{T�l����.Y�4;3�2�����\����|GX�ٳ�#���P���I�f��|��-8	�E��"NO4��/$�!�`8Z[hC�A����y	q1�B�7��K�ɰ��M=Co��I�.,����������ݪV]��s�V�þ�3���]�2�	@7R���m.!��@H�1en��X���@7�~9G�a����z#/d�}�1O|~j�k�#WD�:+�"��*�R��fFD"�������4%������`i,��!M_[�T''��裸��hf�wtji2ܟ�/aLh�c-�sj��+����t�B�J�����bz++��6���xr���|ߓ�c�\G�g�1���I�P�˩�G�/����S`����GAilg��陛 ��?8恶D|#��=�� �9�H�$�
޲X~��� m\+Pc�6V����@n��Y�Bt���Pt?���Y��+������M�	�,���N�_��l����9�
�)o���5���\o"Uj1Yr�E��Л��
Y�7�*���	(�6M��^�-m��*��w"wY���IL�l�%�� Ϩ�D�sD-�f�8S�~��~��EЧ��Lz%���a
V�t��"	1�|\8L�k���V�Jq�퓃����R$�1����KԹJ���1ۗ��w�N�����vOȧK��g2����y=6%�ԑϣ�>>�[U]��e��B�@?t5�
����P�8��<0�s�|��2�Ƀs��l!��W�LE�t�M!�(�EPS
3`FЋB`�3+'��k��(���GK����oiMHX	5ݨ����	� ����Ϡ���)�i�ܜޝs��-�-֒>Hkҏ���UIX���7��:A ���Y����LY�%�������<��P"k���+�&���x�a��IZ�t�`��K��Z<flwvL��tH�7�U5G}�U�ٷ����K�=:��)���zE��B���H�"N�5Q3��[��\}�T��Gt�ځ��{�����+	��	��r����$0���+Wc��,Ukwn�G�_�Fu6��(M,�X�Y0���^i��&Zop%�9D����	|�U�)Τ~\��w-�T��.����CXW�R��#�ueo�d�.@�-�|>t{@R��E�%yt�V;��,������o�d�XF6~IL��4tr�!��C�����K���u3��Sۀ��j=t���T��!�y���p�v��j���1��|��<�@ݵ����@���r�6���7e��~m��������[}�bo}�g�M�m�)��z5��)�?�3���������YzP��e�X�!~.��'Q�@��{:M�ڕ���6h�� ���s�"}+���s�z�um3��Ι��"��{���Q&�j��t��{��H�#G�v&�G��?�hK�:8!8��R��b�������wȹ�1�
��3�C�]�_�X AUHF�ʏ�D� �0ŝj��Pˬ�C�/�;	 ��Ϛ��0��#��0��T'��n4(xZ�JK�c�s�|�2�y	�U�<�S�цg��$���_;�/�h�UiI$!�����|9H/:yuhhab�ȡ�:���N����3��o�L�5/5��T�Z�0I7|A1�6V��eI�����8���i�/��|��^ߴ��QDzϠ=�'p�D�/���I�c� (tܐ'
߿<�t���(���]%�y̿�d�ÝU�dš韶��GO��?yZ�)D��X�HW*d�j��2e�mǔ�L���}:pdd�z�)�O�A��������N���}�c���G���P{�x���܈������8�U��g����Q~`�'5o�(���U;���9�ڙM	c���4��M�NHҘ�/Hϟ�t�S9p��=�K�Ĥ�f��]l	f���,ЪC���b��yQ����0�LMdt&2M�Q(��׶�e�SHaC��Cm�m�Rq�Q5��0p���}�5�:=Gb���8��Я7Ձ�������$x�iYѵ`s��i*��D�D�f�G6�Z'�Ҫ]\;z��t*}m�귐����3�~%Ǌu�F|O
���k^8�8B���	���}�|9Q�#��A����#K��ث��e*H )I8h���m��\O�t:W
Hvm�8lX���<�[GI��D])S`��}������Z#���"_���5Y\�����kž�j��}�xA�`�2%y��w+���a�Y���4pH���%EY��j�뤼����b�|gk��ݡ�$���)64){^�5ȀM
:�Y���%��c�{�:
���8�F]]��SVk! <�鈝*��.
r�ql�R�_�BM�%ɦ
\P��V�7���c�њ���s~{@^�o��Rz��g�sv���r�(�(��B�� 3�T/u��k^�{��B��F�#aɺָ���A!seα�p�I�w���������T,�1� �T!�Q��e���F��+��/��R*{1A5G�jt�/�Mkg$���P�>Mz̴��z�)� y+Nz�+/�{�f���h�g�Y$~��S��./�)�g÷{NGM��Ծ Cj˱Ge����Ɍӏ�Ga�Wo��?֭�J�'�z�3I���h��:v��k�����2�Ժ�P���i��î�y�侘��� �"��p�<�)7�ڲfNt��+�(?j��3U�	,Sm���ږ��Q$=�ʰ~I-�z�;��-F;e8e����@��df �L�Lʄ/OfW�:2�����%�4"��G�0���m/����L"�0t*Cj��Q�a�����i�Xء7��h��_gP�:c��R?I�/#�KZ��땡4ᡓ��H�71xN��?�^,g���o8�w:����5�,m���+rS�WD褼� �I�Y] �C�^��#X�ϣ����,�G��ʛzS����]f����q) �"�W�Ei��Fy���f����"��V�.N�t�IQ�یh���e��-���S<���5����w���#�+�c90���f��u�6.:Ѭ�������Xsy+�4�7������1RY��c��%q%*\!��8dA4ޕs���!s�&�CUj_9���v
��yb���)/�غ�0,L��*:�u�/4���{c��k�z���KX�Y�53���z̑0 e�T�-YZ4!�U
�@tQY�k�T��x����F��i�8X��M�qOs�H{V�����Iw����t=�6�kh*��isW���$w����Ѕ��1.��-]� �6,C����P��&�ĀdBW��z��N��Ȣf�Y��%��}f0ܻ����c����b��05���!pa�*�WT�����+)1ƴ��@��?Fj��9F�XnR�Mf�<��άeg��ծ�ӹOkĝ�t��j�'���"}���{Nd<=���D�~tċ��-���7�� �rn�EH�oq��5��^B�6�薫��Ǭ.5��Ձ
u�&�Z1���ȊɣI��q�xEq���J����ɢԷ���.I�zƟ���5B�^�<�5n;����w�5�����Ws���B�P���t圤����9*����~��Q�������w��I;�M`Sw9�끧ru�S�E�?r��M����!�rl�JYÒx���m{��b"r�LU�����"Z݅s�|�B5�;i�׋�'���}T:�=���s����4%՞�Bkw�fT̎���P�5+��{��yL�=ar��/�4��.bn:�՝�~` �bJ3�8�)���Z�Fc�p>�5�<+Eb�)ۮ)��,'Õ�WrQ+0���&*ը�u���"��?S��0D>�O�7��xϞi�N��6ShF0]w���{B��L������5�z�$ϭ��PP�PF�ekVu�'�[���s&�=�`^�r�U�-�-���,�WaKKy�0�*v��x�$��f����LA��@��n�Eɍ����GF��{���'1G+���M\�9UJ�D4��
hL��YE𽂴ϩX�s���t����c�|hr�) �6�wal6��ݶ�I>�'����Xg�<<#��b��/�]ǰ7�p����
�;nD8�2�'�����9_��]-�P�9}��bM�N"gc۪��,����0����bor}��}LZ+����a��d]���3��v&ؤq�I�b�(:����hKT/�g��D�mF��4Ɗ�]T�: �_��.t� ݑ����{�m��ɵ9\Y�p�E����r�^��|ID����uq�����!ֻcl�̅<k��i�N��6��0�g��t�&f��/'A�h��HvO�Va��m$�}��Ƶk%�J��,�AB�陸�R?�)��W��6�;�苭��Y���х���r]�5�a4$�cg��]]���w��z�벧nj��v��<C��.��@M��󧯁ӥ?��yG��|?v.,lϏ�֍��T�'r�2 +dK����6٪��F�h�̀�	���f�Q6Nz�R�,D�S���l��Mis��E��������n�94����'1D�`�������N�Zq}A�Mh^�s)W��L��S-h�R$\��3��:2�:�M��P�xr�z*'���U�X�EeQ�ܐP�7e�q�R�w�ĶJ�"w	ق![����F�>	�wO��O`
�?R֍>4X8�?Dm�z<��!Kuľ_aT}}��w�����}k*\\���ģ�bˎ)QZ�C��6'�y4�Ē��B�(�zzr�"�QE��/�2�`�Q��֪uf�;~����"�EØoz�L�A�)�f�:�O�֋X�ݶ'�e�<��9�a}�%�E���_%�eI�!���ĵǭ&GT`f��&�0pۭp/ܩ][�nI��_Մ���%���rQr-��f0��'�؉����,ޭ0�!^9���U�{��,��.ړR���.EԌ�<ԞJ�u�R����Шsk�8�5Y	�u|���c�����L����Y�rLĐ��sq�"Ώ�(��4�Hi�I3�u,4�G{�(��;�J-/ڱ�T�}�XӍ�q�S��U�0�r.xLXRy�]*���w�T����˱�Z��(�9����D�ǹ�Fmbtc��߸�|@�n3n]��2�$M�1yMWB���g��\�E)���fwF^-�@dDh�A��'!�fX�pP�b)���'&³��4��v"�.`}�C�:$�[��L0�kd��	-�|�����;`�j��:�w�B�|�KYf�D~�~���RفeB�,f�k[��p�$3�	 wR.��\
v⎡���p�$�p�� �~�>��i�-�P'9�>���Sl�<��'����B��sﱯg�l�'�;!�[�D�@�h|����}�b<*�K�r������=��Kd��tJL��jے�[��	y@̬$Fz�Ǯ,�o�S*���K���Hk��̗o��͒A+�Z ���������-���^I���蜤��&Q;�OB��ҔA�fw`�~9�,�ʅ�bg$��:"��S��X�%����FN�H� C�.�P?�SCK4_��N�29�h�a����E$�6X9��/��w%�U$�ޤ���U�*Ke��B+罪h,;5����Τ�8�X:t��;��l��08
P"a�W����Q�O|��^�n�GՁDf�.�����ݏ_֊���]���pH�؂��UH��%�
�t3��"MrY_�0o��QYߊkZYϔ��;�>RAz�vIj,'������(���Ij�:��]x�\�!R;/�t��D?-|�f�"�p�k��;* �@���u��܅<��xEߖX��kǅk��pk�ѣ��CC�,��>QRn[�Ņq�K�<\3�%����+ǃ -�hD�(�$/_F��r�w���ޘ���KN����t�Q�)�H�õ��'B�q�����CS1�6�J�Y]|"�&�"���C�H>�ܗ����O�t<��&tr�z �Y̊����Sq�=��/IƶO+�[XBT'�Q}o�݂.��f�=ןɱ�f�����r&��c����?���E5%'�͈?m������q��$a��PEwr�O�omՁ��k���CX���{���x;�~�d��������$��S������l�!r��m����W��WSEY�u�b��9�,���AK��̳�sϥ{ド�L��BŜ���1	������5��
W1���z`n;�2|��pl�A��-���"�.���&G����˩�&d�7���8���+*�ט�N#���^Sy�h��JV3���g^o��ywG�!l��kNe����k���n�3Y�I���]���U+��2�<�Rm���6��.����F;�ɒ�1���u�\�[��j�;N(M�1-���\�-2�۾JRk����D�aW����F1����am�a�:��"�F>����H�.iM�$�Z�|'T�m�8�7��yסr[�ȷ3�0��?�=P������n�ϯU�U很��8X�>qz'%#�2Q�~	4i�Α\�f�O�����h2�|�� �sRCЀ����B-�_Pl�;_M���bM����%�&]0���]�c����=�<0�	�C�a{� Yw��y��C�'��W1��ށ��:�~�����9��2̔3��C��ݶ�G�o��Y�r���F��.}
�2޺�W�-�r�̴ ��tڣ8������[!�"n�%��o�ߥ9��M� �������`��ё*g��T���g��|d贍P�V�I{/|M,�SR,}��Gl׻�'v'��� �b�ucy�0��y�|C+�9q|
�Q��Yeo���=I"�}�d��F\�>�<9m��$y����C�j�7�ވ(�f���I�Z����a����MIX��,
��jY�ӌ����2@�ٳq�yκn+���s[�)�e͌�F�~�q�����)�J��:����s�6�#����_��،~Ա�z�;H��`5eLIa�����j.�3d�TM�P=��e	k�r$�Ilq`M��\�
f)�� ����?�Z70)=ƓL.�TM���G�_4��HCJx�ߒZy��ˣmڑ&�Р�n���2sr���	]:��=<�r�0&[7��C���&����ec�p͜����J��a�O���!	��u�I٭^��&�����C̳6o��G�h���������b���`��8�i�u��9�c�����_8�/�9�@�fxF�`���d��8��ī2�)�J���&��8�W�g�y� ��`�A��4����=��D�M���1�]B��QY3�Slv�.ym��0��8�@E*`K-�(`���)��>�I�'���� 6m4ʜJ�h�MV]#���r���b�#���b��X�,阨LBs��C6|����<!��;�Z"�������%V����9g����J+����1�̶��i�Y����0Fa�4�F�����l����9�i9�T�[����WЊ�ˏ'��(�)���C�C>rn�����M�B� z�,�p� �"�]�|���v݀�K�+�G0'� 
$�om���*���2���9�F�F8�����My��oR;�"�$%�r� �O�n����*�VRrG�~~� �[A����%��KRP��Õ\�\�ɽ�E�{��C���9�mR� p��I�C�ԩ�^R2:����jq��3U̷q�YW�v}�gŪ���#y���rFGAf��Z�G��Dک���N|�v�}J������l�?K{h�%�ٰ��v#1��c�;�W1�B��B����}��"�3�˦�	WOo��/\�et��2�q_���.��Ӛ�܎���2�,�+SJc�1=�׳��JA+u�ұY�J�5�#D�}�G�z�	HI�<�ϲk���̸���$oxF��
�;`��[��\]�=���e��m�,�?r��^����)�y��NQ�0u\|���9��	9*�[��{�yx�[������B������p�:��xݰ~�X�օOŻ@�g��I²^N�:��u 6����Q8�/9��S%{q��'`5��te��n�{�w�씇5����y�w�3�I)qrA�pd�F��E,�������&��L�rIF��y�4`NIa�P0����0F���sF�}�e��,ۊ�����EJ�z��S�K��[�gى�)�:���0��@��^9���E���:rI9x�J87�:�t``E7�.O3��Nw�x��HO����γ��k���p~@f�Y0fQ�Y/@{�?*��{���_%CoE��욗3Y�ܨy�Lr�d�#~w��-9�9p-�5���ݷ$�Ψ�.\�u��v���k����}��B�W��~�V��4�NkyT囜Fx�~��M��\�Yv�C{K���D��%�w7��^�m qF����rO.iQ��'��|��rs��ȉ��3��8|@�&�ͥ�#}["կz���5	:Bca/h��Bv×q�G�эMp8�@�m-�S�8��=]:�F�l*π�߬m
j�i��gV����u��#��<v<����]��t�Μ\I?Qȅ�lQ��r�����,�7��G���H��ъw�jB9+��f�$�7�������(�5/�NA��o���a�_Ҭ�$+��|��F���{1!8���Nz�	'�/@��|��-en͓aE( ����ۘ0����9��|q�������.���Ōd�9��\�s$�T���6��ܱ�:t59� k8i�l�J����͙�ǁ2�fn�N�/l��*r�Ka���!P�98Y�����~�ј-�}�ݡ��V���C�_��&B�>{�f�����F)�	�yؖ��/�\�,
��d�j���~��Ӂ	ƸI8�s������/u�C���cy���c6�4������ђ�U��� a���}����L�=��pܓ�h��3���_eFg�Z��|\8RNk��!AK�lg���2�4f���z��!�^tO�Z߻�ss�w�6QI��5�\G�%�I{��_
�R��\�����,�+š�u�-q�klp&���\�4�F]�Bg\���c�χ�8yѴ�;�{�F3��^�J��"�#�t���?��܏���ٔ����?_]�9�9|]�=+�m:PrŊT��
f�U�T�%�w�V�)���|���Hv'$x(�/�\1��i�R�X��R`y��s1Z 6�:��"ʑ����FŤ�����e���C�,ͫOV:��L,&�*��d{�J3|�]��7Q�+�RF�;��*x��Q���&������U�� �+F�����M�jk��J�iR�q�8x_'�;'��w�ܛ�`S��8�R<r���?S��uRgw-Ma�:Q�B��BSa�N��p��ߞ-Ѯx5�qW�m����lqǿj׉I��žW�
�"oFj�*�x
��kRȖj%�/����Y%'M߃ѼÿI4*b����]���MyE'�8�H��J"�h�9�K��R�?�p�zvort�qz<�n|*�׾R�9�F���>O{�������O&�P�lQ�E3���2��0@�>`K�`L�j���h�)�0��$4#����i�8e�,�r��\./�n� m��~����8���/�+�U*�g2�6ń/Ky����m
��;���1O�x�.P�G��BݹKR��Q���ȏ���)A�g����zl]����G�AxԠ��q5^���"����D����ݪGjU�C�w�LſW9���6�A=o�ЃP
���~W=��e��A�_'R)J!���x��N���V�`���u.G�i��R�u�X2�H���p�S��_���ۅ-�+�[>*1Ś^J�<�bo�6qx!_U�$�2�Ks����������XA#xrfه�̛�֖^A��	*��Å% oA�N��Ե�Z6:�Юa��{�%	�w�w���D�B;ogCm0�3S�� Ҍ1�������')ؐ�JI|�qKB�W4I4\����6.��"�7�8Q+��Aj�2j���uv��t�>������g�cF5�M����[���l���<n�X|r4\�q�-	=��+��o�?�"��#�t�����[�\�[N���Ǿi�:���;��y���؈��M���ƀ�	Ͷo���Cp�`�K����I������T@8	Vg�w���%��E�h��v �7U��HE�f$����$�/��}�^�8�#�K�m�{���r���k˟�`^W�O(��� )����W� �h�����kk�_⓳n:�����ͷR�*�
��*�Q?t�q�V\���TU���g��^l	ڦ�U�����[�h�z+���R.�-����t���Y5�u���E�@�h�Y�Q�0㰃Ԁrh�!�8#k�a}r�� �s[�z�>���4F^�ң�
7���:�o��4E����6"\�� 7�+�S;
ee����}��
��g�1"Һ�Cc�pk�O5_��:��j*�8�,�(WE�B(֪��N����`�jC�߹LO:�v|pX�/h�fN<�6�b܋�� �e<}���'A�;�,w��^BҶHw��C-c{3%t�	�/-��ȱ3���/��T�iP��R�۪H��yU��ۥm��vZēD�ri�(Z�*�w8eB�<v�n���"�2�@�gG�m+�y�q�;>�J�aK$�f����ɨ,y�IT�3]���1���	��_c��?h�{�I�-A�9�GzP�d���رSN��=��ބài�d�:��v����N�����C�Դ��g����!8Aw"��E=1�@�w�pL����^z�??��+/�+���
��������$����,��z�����t3�������Bέ��Ŀ>�#�#��(����
�[cS�<��� T����B��aJ�t�īF�F�K�1�����;Ơ��>��գ)�y����D=�ⵓf*қ�4ܝ�eGrF��!���J������0�V�w<�l0�>�iD�*��˹<�������(��W� $�g)ٽ��$fWԈ\@�,Jb<�z�4��,�3�J�핕��6��Fi� 0��޸�/1)n���̋f��[JS��I��p�����HWX�Wu��]�D(�6�ץ0VX0)O�ɇN����+�]z�}��*T���ހ�ȫ+7��d�� �yS�
��9�W���1yG�+$�h.D� ���U��L\�Vl{8��I���:���V�̦�rs�I1G�41.X���3Č�\U�+��otW�?���������
0�+ʦ^&�9<I/�v��Gr�V\SܵgxY�Dr�T�"��u8���[�����N���,�g&ل��*
9�z�DhWRp�k�όz�̠��V��u�r�d���n|���ի� �#11<W>��ߥ(X����񭗶�	�S�����8��O��{&.n+��D�_bzB�+�l1{B�a�d��8�[��#�^��}�ux��o��	��8�&	�\Hѿ��U)���B�W�P8KFM1שB�����X�L�C�c��d�?L�S�.�����w�k�\�&Є��D�-���Y_�^�{�XĶ,+��ߙkN�gbG�-�uDo3�~EUu`� B�h?ٗ�U�;�����-��BBTg8�
�>V�0�|��� �p4&9�Mu�ֹ~��)�H����X+��KD�C�e�Pl֔��J�M=�d�y�\5W�X����EA�"�(Z�NI��g<�Y�Ў�P���D��$y����3�$)����溄��-AW�Xkf���C0��XǺ��,C&��;�-���׳�c�X���/��V�u8�d��8%��_����pC�ޖ��,@9�3rZX��C#2!HT��Na�e:��T-W��ډ-h\�Zs�
�����	�5���G��۪cU]���=����m&-Yp)�Vm�-��sWU�i�3W���t_HC���Y�+O&�����Bg��� ����6�K����o���a	��k�]B�͏D<�UY(1�$%Ԙw��17$Bŵwq3�,��OO��g\���*$���:�lg��)����t���;�Q��G�Rj��P?W�~Mw�C�n�"��y���!���9�ĩc4���E��σ^���˞�3��T�+c�*!=��2:*p�A�T��p��E�Q����?���|�?�6���qыy�f_e����vT�@��mi&�	��)$ϖu�	l�_x�'=�}�&V0y���ɔ�TY1��� s��WE���<���`ܗ��"o�{�>[Q{OZ�� ����;�:D�tF����G�؉l?�@�\��ck�����b/ˍ=��^�yG՛&���'"7{�n�k��`�*�� D,�D��9c�k�d'���ݫ�xXC$�Yϻ�1���Ӻ���E���ؿr��ɻ;/��S���e�󮁣 R`�D�/���W��(�\��5 ���\�R�z��qe(���I��i��R��7��w�!�w��~�Կ��߫�w�����A�?�9�q�Y�̻8�����i�'��}j��l�U������O<u��s�Is3�`����ރL@P,s��i���R*��kq�j'�ѷtΓ� �҆B� K�H[�BE��x"z'��O�v�+��L�~��D��I��p�l-�h�$�>P��s�Ԩ/�����d�e-��7�� jSH������<��9���J{�Z+fBDh[�\t:��`{}ج��_�"���-�%U�
�NN��scZV$�*j~n��� %�,Cܳ}Yfw��.8-��R+K�/@�Xu�g������k���.���i�B1Lß%������诺D�-T��b�^�GX�e��'��ᓄ�H������w.��{2��b�.�e�nD.�8�xWz��+z�i���j�:��Ӽy�AI�*���F�^,}9%� ���@��X���F]y�񜧨4�{�ù�UH@b�V�@�]��:�_SA(e�X�]!)�1͛�^|�%_�t�x�7���x@��^*f��4�tW�j�5qg);�P��4e�� �����n�5|l�3���gc�J�i��>�spK�v㩀��B�_8�`�s�%}���D�g�9Ē`�\�oe���R����'֣��0P�3� N|�$��.c�V�_���
K&��Za������sy��n|l��{H�|D3ư�勚z	����yv�~�hR;˨���i�����'�R��\v�}$�'�-<��|�r���l��h�Ȧ��Ᶎ�ԣ|?ĉx1�[�"e��y�k SJڏ%$n�]��� �#��ho�Ja[HI劯�aKjRQi�ٺ��&��C���UZ�H�\'� ����u���Gd�\M9m�*l��g�ю��O���ǿI�)Tt�c4����d�\�=�>6J��̭���XT\���J(��of�`j�r��j�py�����@��Z���<Z为3z�}�p}���+����s嵣�2��`H�|p�`2�\�C�I��5����Ui���|�w�| ���ʲ�Y����^�:t1a$c��z�6�W�pT>�W5�7��|��JyߊE�J.��(�{X����ʢyWP����ɠ���#jT�9}�'�M=���j�H�-��o�9��Ŕ3{rna,3�NnP��U ��J!�2��Eʮ6n��=���[����@X��#��	�b���x
��@k�B��M>�4wz5K�C��8��O,oڳ҂'�����CБ����"4�?�$dOB�1�=`B�p9�[p�-&�#���\m�x�ͷB4��<⮨%.ܻ�IIg�S���[λ ���G��c��c���u���}�yq�&()��$y�u���n=��Z�a��}PʝP͍��ѓB1�E�X��n�U�:����\��G������w��Ft~	A�B ���m�x���Y�2Ӽ.�d��h���DǏN����,2c�q�|q|�Ր�u?(x�C���tSkG�i��R'�*X5�&{r!n|~m�|�(L�9���OLPx��4ų�����j�u���F+��7�����F������>���3 � ��!�gD�7��!�T��:ޠ��]��N*	<��`��ţ�J�O��MX���'�:�� ��e����^������î"{%7� �8�RX=�Oİ��~V� ��?���מ�
�����NU7�2�7y�#�ef��d�2��}:v"���1q���Q��k��#3�I�(����bB���LߤZ��~�h�RO����\��o��_]{���%���ݐ驀�^]��^F�xq]�h���2'��+��*Z�,[�uՅ�S4L+�?E����<���*�@p��Zcs�,bƷυke�$���D�)��S*|�Ib��Q��Kss)7�F�
Qv�-,N�}R�22|�M}BZj����>��5��"�/y~/�z�x����|�7?s��M�.�o�bm���Qq9�as"�����2�-T<�Rx6fI�s�E�(-��r=w��/cP!��a������� &8P�X��j���ӷ�M�U��[�!�k�A��b��,>�"x��3��p�j8����vk*�>JJZ�d�v�a���i6�.8����'�����v��fj8!<��["��p��~�0���`�Gu��Rx��%�m-I0�bok�#Lm(p�W�w��t����@b3cS7�0�p��4�oCהMQ�`��N��n0A�!ˈ�2/[U���+/�d�Sʑۣ��6�i���Y����~!(�gA���o����kr�j��2j�!=s�6Ն���,c���<a��������h�׶��E��E���t�+6ܭ0�����ח�~�W���~��e�n��F���}����? ��
ѐ��A|�HO��x>Jhqu-*|�?�E���S�t?س�x���8	aM�]��lWH` ���Sj��䄕Z�]�o*_qn�ڷ$�L�.�%���:� ?�����@J?]bg�7�"꒣Ҿ8�s9�d�������F��@�nrO��v�@^G�=��z����d�H1 ����`a$P��\��� <�FS%;� 37�/����#q���,&�c"@��Y�*EX4�!���e�L^j�u��B�A���l��_��X�ʺ���Z����/N�(�M��|��4P2\c�:����()I���I��}:v�j��������^�ӾV��T %�p�mCxu����$�z��HB�����[�m8���0W̠�z[�?Cz^bO�����޸F�&趟걝*���Ӗ���6i��K�����?A ax�qzk��p��Ӕ�:�(y �����{DQzA�}��4U庄ԇ֡o��H��D�2J;�L|pr���Tc}Ғb�֛�:�S�_2~^��,����z[�ǹ�9�޹�Z��_/(���/O����6`ɔ��a6M����>�����9F���� �+85Ka4]�>:>������\{&0Ƌ�<���lbܑ-��0��3�:�%H��晍\�R)�K�p��:�
����7��!��Mɂ��WLX�?/I��ʐ�zQQ�����~=�7PAi��絰u�
D������EToS�q���J\�UQC�f5Ԟ=Ȋ�����uRn��S���̢6�9���{��$U!e�'B`��O�L6��䣍���E����Qom�4��M��%lu�?�Lg� Q�t�����/M�-1���L�X��'����K"�A�4��HF)~Yh�5�B����W� k�KH�;Մc�/���l�x�뢫:w�}���A�jm�X��ndb�3��'�)Ȳ���	8���0�b7��TX�y[;���M�#8�
V���`U�<�O�]��+�]�~(}����\�#[r9{��\��V�� ��u�6~�Xe���e}:I�28&��e,z��H�-?�(���'�gGE�����􉢕���d�V!����9��;�4�-~��ܕʐ��ZꉿR7KBZb�|�P��u=)1���{٬�$��ێ���2k.~]I/�OT~f��_�lqR%� "G\�4���ϦLR���C)��0@�����ӽ��GX¯o�u0������A��R��5��v��nlr��(@�~�U�>z�F-|m�!F3�Ť�[ X<6-�b��QW�t�㽀K�xUĂw[�3�߉�	[�o�����eX/�g$�_Ӿ�J�Ჱֳ}�[���V�$V -.U%���+�
Ȉ�l(��K��/jX�, �oH��eC���8vi��h�����s9�y�̹��亰]�vc��U���g��,���*�UF�x��v1_�AĦ7º,z=�F��r�{I@�w�蝬���Nq���l5�H��3U����%yOp.h�� ѷb}Q �Q"�E���h���(��c�Ŧ�ltkd&�	u�@x@u��t��=:�+��oo�ށ�f[t�c\����V`KF����r�#�I:����P[�FT�h�� �����u?u�t濻x�M��1pݜ��j�I����2���`�ao�s�	m�d��� � �&-+#.P�c�m�9ޠ�g�0��S��EoV��\I¤�q�d��T�a���^;Z���p�\��έ}<�:]wg�Y���܊?D��D���ZCȵV^t��%h���֊9g-�j��� Q=�_c�⑓1h�Z�<�LŦ7c�d�a��`�B��V�ØL8�MP_�{~r`ȸ��xɖ�๟�`J|�Cz�z����XTk�r���on�.��:���!�P�u�	ko����^��Jz�kG�	�c�gf:�e�']i�,�k"����V��^R�Y��c�P�4C�IpC�	�r����������5�%�S���f���"�����C`z�*����a�B�.�-���֑J��u<t�Θ�o��dLc�G�ܵ�CYF����G'��4Q���8��D��P{9�������pg@�`�O{�$EE�-�%4*{��Vj��q��@�Mx�&�ᔔeD�a�e����f^�0ԉ���n�:߼�R��n��%%'���(�n7�Z�36��ے�Ӫ�_A�c���w��]H*z���}%`;S�;S�A��y������2wj�M�� �\D5�_�7չ0�^���+��Sy����̻�����=U���4�Z��%x#�`[�������1%sS�r޹Pߎ-�~M��T�s�/IxyT�7~�X��-<�ZT��tW1�p�I3���*���aO:3!E)թ���U����j0���c��O�u����wA�T�A�� �V|�H���/UF��giK#2�8o>�텊E��SZ{%1v#U�ۘ ����v���&�6}���=��Ŗդ��VM3Y�F;k.�������2�e�����8���1�oΚr9/�tُ��w1�v fZ u��g�c%����E\v�`>	w��o,���y7����FDR�#��
m�6��k���Y��W��Ӓ�X�N韃sA��^e�������8� �޵U�=~��nc��!%S�ic�P�x����������}{/�.�
yʼT-PN����c�X`E�%���PM�o�����ؘ�gg�Aɸ ��:٠)��6l�j��@�TWi�*�$�/�h+E����G�C �O�N�\[n�0��4�K�Ǘ������_P��;A���Eg� �3����K=�W?[�b��԰r����_�.{��S�F�n�r|�"�v%�?!_��
oyM�q'�hAJG�W?��Kf�_s�����{"�[����1\�g�@��`ǗTr��6��m�9��)y�c�ܛ��.p��[��3���pxaFSAͽ�g
�}�	Ĝe����cWv5���"�d?F�-�Q�A�r��-���=�f{� M�n�((e�fȍŠ�p@����������M��U<�l����M�s�.����Edg8�`�vfx&߮�[��_��+l#=Or�mҜ��v�2k��]��k�����c�(���;��m�]3�I�ѥ�R�Zs��2*����Us�1����%�h1���B����Ny�����E��@]��������|�wRw���-�&Aq���L�j/�T��ȹVL�k6q��_���Ep�3�6U�o�JZ��!��fBn.�Zs2��]&D5��D=�!�,�V�D7���<h�WkS֒8���x�G�⹮��:�2#���`���c�1֐��yq���i�F`��k��I{���z�ޠ��ڣ���Q����Ȩ��h�͛���"��O����
�2h��i `��X���e�h�CD��2�o��xV�����
�;tO4�>��'����$��.An��©2����g�t�Ё��?�o�7����Ƌ��#rW���_1�
�!ma�����.�W�W0��d��gI�38�Vg۩*ӆ��Ejg���ߣ���H���Z�����������U�ɃY����^ ��z���lP������s0RW?���|��U�_=�X9��xm��y� ��WgWW��Gd9=�����/�V=Zb%Z�LO���~+X���	�wI^f��S"��^C�̆�*e\���+���0�+3rQQ�Y�y�P��*�����>����V&����4��v1�A��������(.ԟnc{��-Q��a�{,�hs�h�
�e�Ǧ���m��\xJg����~����F\1>Hy���	���q�V�K�x1��T�Gn�~@�����D@��i��* ,( i&L���t>�"Tèۻ��|�8L����!B˦�φA�.rY<���k�ٰϟJ�u\�
MoW{����8�����Jw��5͍�A�ζ����{$�k�K%t�n���>��O���Դ�tI	I�F�S�%�a(�vp�,W
0�i��/O>��˗[ƹ^�V���H��\r�
��R9G�w�q��{��{o:q9�W���I󭁊Bc�91W΍rJG+��R'�Q�0M�2xly�͝�,=���9W����\�;OE�iKְ��=���/�+̈=��lK��� f�0L8�am�,��~���d����[	�s���g���	A�zj(Y3C?Ձ������a�h{���V-/;KX���ҞD��zcZ�榷UdL	�fP����Ϩo�v��n:���ň���r����C�7�Kf���KT���zt�S����3�v�����f���Qf�QU��T����>>�i3�r���e��a�X�vy�kmn�P�'ǟ��&�Y��Ds)��sS���c4R"�8Ƃb�!�W��E4p��cE��:�y�B�r�Q^���t��h(�ju/`��a����u�0W�����6n^֋Q����=��__�����S*29U�ފs����,f���J��+æ1RA�թLQ9�J�(N_y�>?1-.PAY�:0s�ƕG�e��/��]X4e(+$fݐMw� ���R��c���T'-!�*��6����6��!�,��3i�@��1YAQ�ǻs<��pj�1>� i�yg�i�0ʾ�so���?�s?"W":b)I;�7�1>[oXess��u�s.�_��0Ī/�Ѓo^�"$=��#)1� �j���$BKD��1�;wd�8�5�?A�Yg��n	붭o}�p�׿.��^:&D�^���Y� �u��7| ~ϑ
���!z�L'�o����S{�R�3��C��Z(�3?x��X� ��AV+�<�`q���W��S��I�'�E�MNI2����+���V�K읹i)�V���I;�>�aS�
� G��룔*���H�MhV綌�p�w�Z,z�����-6������ih���Pn�LL�h�hk����~�&�e�@�z���#��#��>fP�.T� �7'<`j�V
�u����q��O;^~'a����Or?�5�KQ�NL߲���{��h�߹?�r�՝��A%�w�R��w�O�*�\e��+��a]�4Q�w���FRFV{�y�g��q�a�L~�[ylT+D���@b8�mC�����k-_M��t�ACϲ�@�l�8rEq ��`7����g�)�f�4N����v�P�XD���;�p�!�o΅ɠM�����T��w�,0�@����{w�|KyKc4�;ĸ�۵����+��=�U̳8�	Y��Z���*���s漸�sl�D��6˩�{-:^H�4�=�o�J���x^0�T��Kf��O�uAa=�~���=ʲ�Z�C� �㓓ϲ-M�CL:�����o����1�a:���/yW��T�U��t����+���`�4��?o2^���,)"b�}�����d�z&�W�e���3�^�G��e�,�/����_�M��_ �KP�T�LH�0��ֈ~H�ILR �P�bR��ꃋ:b�]qt�tI��i�um{��bn��[�g4k|�>��Q�]6DJ�wP��6�C$)�;}���{���(r5� ��L3L;7�?@O��c�\�����-ۖ���pI�2�=BA�$m�?vE5�]$�����f�������L��iX�M�P����RRO�X[�'^c9���u%F�����F�}� ��b
��Ky8g�<�bp�6h�~��&/	�D�h_,x�Q���D�g�O�0�Ypx-x�����GKN��(���G�#Ur
��g;{�E��F�n�9�'6^�� �L��&�b��Pꭘ�v�+ɧw����+=v��n�X�%Zx��AK�I�מ`�H�_j���Q99��dHv�E3F����E|���R��T����Js�G�oT /=,�Ȗq�-�s�7�Sy���-Uh�o��0��m&O���A�N����D23�EM�_Ĵ]��n�f�'�u�"Qᅍ�H�#��H����f��}7n&b;U�1�������ag/3�G�S����a�-��m��٫�yO
�=b+�������i�J\#�����(J��<F�E��ϝ#�m�NG|O��řuFe�t|�x��i�,�!��t�ÿ�S�+[՟Xӽ�cM~���Ck�U�f��.�}Υ�L�׬p��SN���Ec�*׭I����P�� ���p�Ќ��������I���~E������X뎥+o�����[��]�PE��2w��=o>�(Y�i�R�H�L��p�r�2�&��eC.0u/A��l�g�6�j��t5������a{�ѯ����t8�T��fE4��s�(P�N�*���F��?�S�j[n����k��UF�U�NL���Ӊ(��j��j��.f�ͥ���ޢ����Gw5)�/��+@\.�Xw���t�AF�����a��-[�BD��-��?R��S����.�z�d�����&<Qy��ܞ����`?oO�YX��p[jx�<�(�'��9L�+F�s��rv��wZu��`K�f�+��}Aˢ̾�9%@��\����泑���d.%���Yiè���Fh�hMu��ԡ�z�_�tJeW�m�_H��dwX�ڹ,X �N鷽t�$�h���k6�V�����ENՙ�R�9��FcmTz �s�����c����ͨ�IaM���z"@OE���^G�j��<Jl<04�Q��T9WI��M�Y"|��*�դ�������Ш2���MKF���t�y�-Ң{9���<[���K�-h�Z	��YL�(0P`t�h�&YzɁ�3�)�e��O��d���e��}Ql~�Z��}K���u��o��(��H휅�S�u�D��m˴<�S<���ڬB�T;��-Y:����G/q�JJ&ߠ a�	F�=Д�#]c����9e�������=$��Φ(UW7c$�h��m��w����H�S'Xv�/Ѓ��C�+��}��3]R.�V����)?��y���lC��$�ɪ8 ��#⺠�c�����r��83�;�=Z2GK/��C��I-�I,�`Pw���9I%�~���������Z1�0d�7�I�u��H�+s&���Qx؅���PKK��Z�:��"��}a�����gw���鶒�m��w���_J{�ciz���ޯ �
�����D�t��Ƨg~Z�g��l��ލzV��2a��`>sl�4< ��w2��a@܆U�#h� �٩B�e:H2�;�*��"7UxR������pX� _4v��PBX4�/��b�m�`��D��m#3��ț~4���L%���/�����T6S�PI�7{���n��VTX/���a~��`���k(C�-�L���w��_�Lj�y
�6}+�u�=�ř�F��Mk|bN�{f���N�"�1H��ۯ3���k�9�S>I��9��p*��2dG�$�� 3�,̭9��Q!�; �>v�;�ӋD���Q�)�	��,��)��[�OR��Q�~uH~H��MX���������ǆ�ss�;�s5>p������d^f�g�Z�s��5�Ŕ�i�DH�!7�:��6:w5R�J\Ir��5瘐E��-���!��wx����`	�k1�0ɫ�O[U� ��)��$װe�������.r�K���lz�t-!��.��Ɵ�gԺ�@��1��'@$�-�#"�bM��ż�~X[���r��~IO�`Sb���i\r��E0'H*����8�,c�7�]#�ǂlc��%6W!^i��{6�!1��4��*>K������`���	#;�c��$}���t��'�fB@�uQ�5|�?O�7Nu���=��26�ஂ;Zʉf�'2^0'���kH:��d�>���=9:-�,	ן S��� 0�>���]��$q���4*��}r�-S��2d���n���2�oD�z�h�s��X�W/��ɼ��R�UHiEYO�j�u>���UH�h,;��$�y)��Kgm��f@�Q\s�%��VC��3����KM4�l�:eVb���M�i�O=�4�zs$���<�ZTN��� ��dHVW�g�3���i�<�bMT�t���	Em�ok��SFJ�5����4���/���1J�����t��H��kv#�-{�qU�������e$��K6.ߎ�`�?F��� ���1��=�Y�Q�ti�wǱ��hQ���֙ ����=P�A�Nt\�w6����q�9-�^�n��s���t��{EpC-��(?��wfYѯ�r���y����ع�}��i̊d:�U*�U�)�2��-!�:��a��a
�?W_�)�R(e��[hܽ�U�|0P�ϣ�����������;���lH� �4c'���VS½~�+n�|�SECo30���2��X�aj_�-n�x����	��u �� B� C̚=<���i�Wd~N'��;Cm+V`�b�hѽ7��
)�"��R�C���i�J���āV�J�'�b�F;����Dj3t82������N�h���N�\�+�sD�D�!9�����I�9.��4q��p�ݢ�1��p���}���9�>r���&o���y��ҺxmxL�������/EE��@$,g�)@�/j��.�j��}�
I7� ����fu��3�*�/��`u0{�k�̔.� �v'w�n�.�(s�;SB���	��oڀ_���Y�4��mj�`���~\a�������X\�y<�y�(L_���rx�?��Ŵw���b�n���Ӊj�X�b9�q����U�y�������;Hru�q
�2��e34�@Y�8^<�'Z�	�|m��
�c85�mĚ�'λ�; �H�,,��p���<�V��:5��3{k��� �<W�(>��g�e�#�{DM��O/�H�����. �,��B"�)Х��#�K��o��WfZ�����Z灸�􉀲�E�j���qѴ�Dd�����=z;�`ro�w���*���ɩ��|�#WK�T�?+��	I���[�x{l��z�H�Z��M'g2N�K\��;d���	���*�5f���L   �] ,]��������8�:)��rB��m��)I(��?!��:b(�/��Q_a���#zrb��"Y���:�^�;�:kG����K �-�[�r����o'}�c���f-K�X�jD��J�wh��ʬFuo��%�~}�8D!�� 5(�����
�ڕ��c�!��Um��bD�j�FǬ�+�Z�S�ћ{��m������'�j�e�v<>LR��/�e����uo-�xl�c��Qߋ׽��N��2gQ�~3s��0GZ����9�Y�c��A�e���P/�5+"$�+ֶ7oʉ���?duU|�Fg��Xmi������L�:�O
O"	�_W�.�(�9>��0|x2��icn���D�hY��D?�'�x�B<.����̤3���$ą<�8I�T��|��9�$���"����og��**�J��$�R����)�?u>lΤ���2)͡�ް0mHI����L�E�ǰ�|��w��l��4���L`'��m�0V1;�d_���z2�����_�'��.~nGב��{#�+�.G�]��')���+j���A�vo�r�6���p7?������5���-�`ѣDi?"Y�!�lHY�^��#��B<�Z4�A;���GW~��>e;��J%�`��?�$\�#M0,�O��N�-A��v�%��\����#�N�&�.�w�d8�!�E�Xec��� �����ۮ�s?�<�2��I�(�$ �h�ڂ�oGig���S��%nQ{�����|���$�:��	���Z7UH^TV�=������y�5Mw�n��L���o��*P<��L�tP�̡&@�����C�M@��2�1��P>���LԞJG�]�������o�V>}�3֎J�Y���1��+A�l�2�r\���`%�]o�"�G2.o�J\H�驣o�b�/��w$jV�n�a���{~�I�S��3��2ҨzV�ws9��Yy�\��=���c!���'[����L��
�`F����;#�/W.���K�Mq�5Uwf�V��h�4�B�w�%ֿ�!#�&
�N'����$��6B�)M,�`�o��9UP0F�N�!{P{9��İLk�G4�|��n�U���~ai��F]@!c�o�;�dˏ�ac-ܛ�҄��W����@%l��ߙ������>��J����3����a�.�B�)�H6M��J7����]�u8H�͵�Dr��ć���3{�����?�fe}��g9�B�Ȁ�r���2:��$�]�</;+����yJ�幘�>��0|�̣M��OΈ�~�D�O�\��<k]@��&;/�ҿF��d����$l�j6�	�;iիE����CaC���ھ�OB��}%������F��#�*2��BmhX���f?��h`���Z6�{���G�(��
��<k?��WZ��Y�=|�~��,����-_�K���'O�'>��&���c�5��L�e%��0t/�C���Z����cJ�1���:
�YO�iC^>��"9%���{\8��S��#�E �sO�G+�x~x3������`Ȇc�&����b�_<,=��c:\���m���z����<�,�q�ZB+:�TK�^ �K$���v`��2V4�\D�?T��\�k��ڪ��P�#�Q��*3�G���a��-N��T�I6�
��y	r.&P��'H�Ʉ�G�@�m�3�7���ξ(CP>L���L+�f\�Ȼ'��/~5Pawo�J�*�����n�.-@�|߳*Ę�7*��3��$y���SS�ڑLt SO��b�|��Y Z	�x�
�K�2UmP8q�ŝ�Y݌0
\��h�e%�G�ha����g4��.�G�=agB�p��ًm{Z*�0�ku�}0>��q�����09
(��%�<_?�{�������C��ݙA͌�'�����I�� {)S׶�2jb�4���H���n5W-���w�@=NQ$"�IJ}�x�������� 7>6�VS�L3�+!I���ɶ<��U�
>Z���ha��r�砤CLw8?6uٹ� 7�/�S�;�� �ԑ���Հw��y8��8]K���fV�!����W��;]��	���/�HO@p��$�����#�.��s�hq"�L��F��)t�G��͚��_l/)2�Ϊ�au)yڅ7�ڼs5]��9k/������}����#dzc�;@�����t{������\H��v�Xsv��H�j>7`����������PS�W��9!��B�~�@3nt�� B�h���P�&t���g$4,+z-��VR:R���8ɂ��d}�~g�_�/n�Z�d�/�&�+��/�/���'~�vKI/[��.��}jrfTGR�+{w�RO�(���0��Y��? ��x��DRt�d%yC,IK��\��)-���Dn�mX�[��O>pR�0�_�Uw�r�	=�V3u,��g���_9�%j}��-�J������XB��Z�6�tR�U�����gupS:zm�S^=F#���6��d�n)Z���Y�O
��g#��^���U�4��X���0�9e�)}I�f^������i��TPL̤.�QZ�^�\�B}9�m�p"�Oti��$��f�����۾����ْ�z��K�F�5��.M|!0:��uF	��MF[�x��ʻ���uU>Y�М�ç��|"�݂�P��`V����w>s���B�\�+�
x�B��S��}�@�6ţ.�-���n2��&�Ÿח=L�lĘ����$��ɦ3=�3=:kI5<@H������U�o��C���ƔD�������-�[ �RlM-0JS�����l�㩒0>�&)C�Vze9Ԧ]�g���E�
�TCs�
�Z�H��'ڙ뽦E�q�#��dVq�y�E���P�)���MU̐��GKUpi�$����T�"��C�{p�QN���O��)/d���'���A?[Z��QQ�3j��}a��5��N�&i��="d �hM�_���|�� �-R����(v�`��*��� ���C������Ի@�����V�,�K{$St�&4ۏ� '��P��D���P�Z�#�p6e�Q����7Q��w�B=��K���Aw�5MYY�b�\.9/�W��`��Id>#�J�/�ݤz]��^�����e9�@>�Y�Z���W6��b�J����M
&��Z|���c�(c#�c�C(�3X=]gf@v�E���j�"�L��;����/q�����p�J���S�H��&���v�g,a+9��9!�z�\��G����l�
��9�`h����f������~E�Nd� �����.7��a�0�(���M�w�F)��6�O�!+wS���Dn�	�PӁO�lDo+��"�N�6�&�r�*iD��Aw� xޣ�����=)����G'����oc�T���f�)�R�U�C�~�����
%��}[>HKHO"S߬A�I_���.[�#e�[=�,c~��2�m:�!����J�|&
z'U�@�I�"eo�Wg�C���6�8 �׎�x.�p *��'��B"��t"%Ԫt��.�n�ARX����@�f�r��5���^�ש���Ⱥ��gqp��|'��K"m]I�-��yB!2�vS�<`I��N@srP������v�[����$��1���M^�B��U�$L�Ae)���k�z��J��{�~�33���k�gU�i��v�8�������GY4�ox�ܙ�׈��Y��IS��tIi
4N
 I�:�����ZV��@�M��d ���lj���3�� r�d�����Ds��hް����b���2/��O��>P�=5Ӛn�^�xTS���h�����	�4[���s�y[�dT�8(�q�:�w~����E;`yΕ��3b�0����<��쟃��YT]�U-s2�iU��?n�����'�	�!Lc�Q
�~�z�V�˅��`�y��c����\|녡56'�R�Z�uY�]q��|(S"K����~ ��W�Ӱ��ð��-(p��������.�8���~�i �g�W�Y� �j\�B���B9�R�Wlݕ/EW�HU���=�o]�?2�<�݌�S�K���~��u�^�5ZW�� &���٤�e�4j�!vc�8��8BE��8�0���|k��j8�wr��Rќk��5g\�UB��f����ފXg.���1?�3�F�GJ�+n����V�ɰ3�2J���T��V��p���
�N�����s�9��2v!w�]��Kdd�!SvC*e�1��7�����×r`ۢ�G�y
����V�wu�x����� ֝�֎�a����^�S�txo�3��(�K+�6��bPG�.��e����M��q����>k�=jsR��O����uW�Dݽ��KQ�6�B��I���\1y���#x��~]_�s�����_� ���aM�a�$Ao� }Gbl`4�>�\��#��w<��#t��3��H��eK���zÿ��}Xr�z�w�,F��SwI�'�臠����(�e���@�D�)z'"7q�O;�qA�4MA�� ����N��KL=�*L���!ĬI^�O�Ů|Zr_!e-�r�&���4(���x�|���Ml�yy4��&�/�՟~=��D�.�z����'�F���$n�anP���������y'ϓI?����\"�-ӣ�ӵ��d{��-����K��Ѝr��xk��#	w�#���fK{杉R���[�4��)���%[�IESaٿ�a_��|����~savk�������f�J>
�F@]��tC����kM�տ�񫉞��4��C�˦j5	%��"6��>�|`l�\�l��}.,�ʿI'��1��]|0RG�\�7I�O��`�R�����b��Ԛ�*�T��do��]E���ӿ�)��e��Ʀ �f����b�x��"��dca�Rԃb�LZ��Y�4�0q�-\���P��Z��}�<&I���aR�iEޖb��e����8s���b��?��� ����.}"0c��{5�xK�y͟��ᠻԮ��fwn�����D��I��z�xU� n�T���ޚ%�q�Mu��i�6�bz�a�{O������pze�������.�^M�>�i�Y�z��o2޴
�.ҽ!������;��m��D$�U�܍⎹f*\�p����78i���t\C�j�-l�l�އl�(��:����ޥ'3��s6-$�{��\�α��_���r���uC� Wɟ��F��r�(%���'�W��hj�SM�lr�����s\dښ��J�DGg�;��9^k��^X?��'����rU�8�2=�-�Iڅ�V����ޕ�G����k�?�yj�1�c�ݓ�~�S+���������ka�T$q�'�´Nn���i���f>kBs�`u���V�N�6+�����4n?��K)��=����q�tf}|���߀a�V`���n��`�[6?26q1��#h�ҭ�x�T ~�����;����噍+/�_`����	O(�|{!l���o�~v7�j��Q�ua��\W�J����y���B�[Z@5�XX���é���
L��8r��^;�Bl����b���Jw�d8p_\��c*�e�b�ÔW����8����U�^��r{j�>�5��)X������^����%$� �����fg�Y4��:�	īf��y!�ݯi�ڐ�X����ݲ^�+�Kb�}�UX,�>��Ҫ�"�Q�p)^<�a�4P	�o
b�T�c�Ȫ"�8�z<�����M���^��NLG�wS2�r{�]���"|ď??c����"n�ӎ��|���;�R�L��a`fr�q(h��Z}gQ�N�bW'*=�~���T��@|��v��-�1�fK{, k�Ż hS	�eU<X��Fe�} �&a�b�	duZ�p�	/��f�@���!"��P� p�ed8��e�ZNY�w�u���R�k�qԡ}����� �??������ѕ	��/�1����as6Ǒ������f�u��s�'-�:ϦF�!�`1no���gfsg���P��#A��-'��%��r �D(��<S�.�9,	}���j+C^��5����֮U�T�m���1O(㧿���܄��M��3T��� ��\�Ϝ/��׭�U�@\���x�d&Q���;e�e�;�{��rF��n|�_�(HF5��� �:�����Ӫ7@I[$�T�J\�W�x9��cB���FD�>���RdN1�e�p�	?Ү�s����ˎo�Qò�"�ܺ":v����M
�������焫 �H��cy5�j�l���p�������7�eŇ���+M�Ah����b#��u�L��;���ꨡV��ry���k�X��;Ō`^�"���q�'n<�;��g��w����$͏.M�o$���-c��d������}jJȐ��΅Y�ͩ?�]ZSa��X5X�s|����Bbf�Jx������Fmȇ=�;�v0=�~�&��اb��	�Y!�ۙ Qf2��k(PY�g	�$|<G~}KkOD��[��%7"�V��ʲ��w �7Ǖ��cnTH�^�H��G�S��}�}@n�ֵ��c �2�vO�.z_���	���H�xv3i�����&i���5u�~������T=L`�yn�(� ��Q���>g�<��p������� ��h��5L����y �J���E^���(U,�	�vQ2.��5(g>�T�_s2�v�O�-ۤ��:��K5�C����=`�
�ٴ�U��������k?9���3mt�)���/\I +�h؏��<�$9*�n.ˁZ⦨�Խ@��K+���6U�M�}��ⲓ����n&$� pJK�Ѭ��-$d��m��pi�t�	A��`;��a_��a����4��T��ת�P���WBd��Z)'(%D�M��{S?��QA�O�W{1AE)�n}@Be��&MRg2VM$��ڐ�z�Sz�LH�K.9�m�����F��)�ҚRގ�Z.�6'N�Q�9��_FUL?��Z�V��f��=f��P��/��w��j7p����U���K<y�����db)��^pvT?Q��A#Q�>p�������R¸���Y�rL)�(O	��b�H�'�%�����?+�\X��n/� G;N��d�R%`�#
Y�K�^)��E��?a+�6�jW���,Aj�C_X���l���G��B�r�|�\1/p�O�F� ��	-��Ŧy�(��������1x��b����d�[�/�܀ٽ;
K�!�&\J1�Kۨm��rm��v�q���=No�h�k^y��}����?��vR��Fɳ�'����������,}��p�1�,;{'J�PҨ�I������6m�Va?�v��w�q�֡��wL���tI��id�p#��=�L�Q��f[��J+�/ �d��q���9؇�Ӧ� �cd��۪�Ȉ���]?�BJ����-p~�ф������_6�?�f�D�Bw��O tl�A����c�{�HOz �u����󟕓�{��l�NQ�y/ݷ��в��k�(�Cg����:.z�F��/�t���D���$Eh���`�ۼ=x�)��16����������`�xp�7ER10X����ѣ���
�<�S���e�9"]U��ĵ8��ES�����3�
tQ[���ZK駯���Hc��t�ǒ�em8�H�Ѐk�^���J𶜭���6�g��1�F1T�jÃ�V���#*o����Ԫ:��x�,do� c�q�U�cN��#���t�IG�!�����7�:m��~�$�B|G{��:/��7-�[��.��<
z�I.a;��q�"�;��q*�0�MP��t����g�W�x���ڀh�.��5�/����;9,�e~�9���G�0�W�׏�(�s�H��e�XC����<u�NH��-��Dr�4u��DV���=Ԣ�� �.��/~��I�&���K���-���Wt���9:�.h֡N�P��(G���9�<�;����;_N�()݈�3�P�f���vJ_L��v���q�UZh�~�v;0�;if����M9���eғ��G4oy�-���3�t��j�ă��u����҈�P����&�8�f p��#\=](�r/*���HxM�>W5����K�j��-�W���J���'�
�]ah�x��_�K��O��0�����ۏ�	���UJB�W^H��jk��/ I9��:V>P�b�?:�a����,\�	��:�O�79'6���5��)«�%ϊ��T�N�b����Ŗ����洦���A<*4p�Y'�pY�W���+��/C���G�����ٯ}�iE�5NI��Y&p�5�n��dJ��m�u� �t�$H<֪�����i������j?�չo�U��(�8\UtA5(�d����+(任�)�+K"]c��*���GQ���9�r��cvA^�%���g���h�/A�)۷He������x\�.���N��	��w��ph�"�������8l�m�^/�� &p����m60 ������/�`s��K���%��*�p��c�f-��C"�(�X�S�B�ύ�Umw#o�d��{�?����>(�T
�K���@���5:��(�h��cLf��� ���L��#E�����
�Y��������	��p�~���������m��2�N'�,��嗽#I��������=E�z}� 8��g����6~��)��������*��w���T9�P_����wg�9:���>�z���!}Ȅ�SSN^����Ŷ����Q7HGo�I�}�CJ�9��ݚ���{�d���Fu�	�9���	�d�  ZP������`��/Y0j���>G�'C��\�Zx�p﷩q���&��Ƹn��qh'�}#X��*Qy'T���o�eF���T�#a�k�RHʾ%���U52UnL�8��i�f�3/�2��?����|���
���wa���Mz�ǈ��أ��4�uZX�����r}�{����Y�^���FW�m�0V�m��.厇a�s��I4t(O�91>f�Nmu!I���^����"���<��x���a��ڗ0!� U�E�g&"g�W��ψFw����%l3ր�V:�~�M�����42�I#��b�Wy��.o��{d��0��\��x�t�xoh��P� �l�O��!)z,!HhG�6���p��ǨәR�he��(�;U���b�����?Z�QI��^#D�RZEƎ�e|�`5nZ�>�3'�9Ou�i(9�՛����]�-�5Ѐ
G���ď��y�E�ޕoO��K�WK�U�\���Z��g h5<�Sgx`w�JۓKy�)͋W&��٦�����e^1�U���c]�@1��n[p���(�'_$kC���H��t�_Ƿ� 9������=�/t2�G���f��#������ʱ�W-�G�oI�ow�����Wv��/�9}ݏ��!�[���G��2��{�yk��Ί�>�`���<���!�d�n��g��ƙcu�rU���o�Lk˗H:VN:�w-�A�ZɎx���1�ժ�
43�g�����d�>�Ed&
 �6z\�\��T\�9�!�����d��r����~ ����=��s?�8 �y�U�N�0m��1կ���#V��X��J�����g6�읻~^�;j�@�3��!��.��:���V�.*�?�7��I��:��۫�Y�ж�#�� �eqJV����r�%��x�� ��v?a"�f�ξ�$#y���Mi��i�Ut6�ʆV�Fo�c�G��G�8��O�a�g%mb�T@���������FfL�����Ʀ���T{����?��� �7>>W��]���������RF��%�3�[��1�K�ߛۍ:��>w�tNk�Md5�{��w��Y���b�&�f���ڰj�4��v	� +��ٻx��_��2��z!��5��%��2��9ʍ�fq�a��,�m�y�, Y�*���˃�4����7���(��/�>3�vPA�4X�{*f��A*��e�#�ͭP�̇
\�D�'�g�۝� ���`����5��ӑ}�5���n�!��`4A�^�k�M����9��~�ɬ_�䯰ꆥS��24���Q߿E��Iؽ��:d5�Q4_�����2^���q�#�es�U��l�0�?_���v�L8��oTmo(7�b�˙\Vy�WN�K�`�l���B��pH۠�"G�2�Gk��rv��
U���t��\�vl���
g�KeN�Ӟؚ����ᡌrv�>~�4��P*�`�gQ4�n�B�E�-���)��q
&\f[=����F��c9s궸�5�U�G�Yy,ܣ�L�X=k�����Oc�7KJab��3��n�`��l&H�kܚ�Ƌ|��
v>/�%�ޤ���vg��P\M����#�D�F��c�=����p5g'A+:_@8�Z���"犰�DALK��9;����܁n��Q,OMm:m?퇿�2��φ9�AR�W�����}��CfE�{2�< B�J�\%���\�v���
"-q=�~(P��p�7���'X?��>>��C]I%И8�#�������.��#@ۚ�֤ע�̭>���D,�L#����Z(�n�����ufӜDo��T�LX��w`�;��v:&�z.�z�CIГ������2�/��L)�RH瑗2BXk���Kx�՛�H�fz��Mp�wEW�6|������
EE#J��jŉD��P˚��?)d/�t�)w�u,������Kz�ļ�ٞ ,t�D�������JϾ�d�@�ƂJ`���ZZrt��>��/������1��ʽ[�h�`�s��o�>&��5��%߯��<�
���8`	?�m$�m?�д���'�n ���[�R�;���t�����R0Ely������*�+�=�0���`����'�].bHq��Oz(�F'�Q�(���C�=��n�%�Dtz(>��ua� fT-ކB��~��#ws!�i�A�g8��4=�ˀ��.����G�(�!`�!I�7nP��O��B9���n�)Qh�;;G����YNܛ2}.Z�'`�Tо7'�����9pv�;� '=]J�c����,(6�$ XQ��#�ǸײADW�56�̊V���w����Fa��d ̏\	2�n��TF,PS���eT�ԃK����=OH׊$?�F�|��!�T����'7����<��8�_�fJl���`���r2�X)�g�VMBe9�S�X������Uqφܞ߯\=&,]�E::���F����u
��Kx����&�J��J��.��2��螖h}7��\h��E�J���tG�d�nR)���L�n��0*�ۜV%2	��K)�8�N�U)��x�v����ş]���ݠ�'2Ya@	3}?/����5�ʦ����,	�cE�L�xCs��EW�zj��b������<�5��ㇹP�3F�O����l�ߢkb>�����^]Asd�c�$�K��1�(����4���~�����Q��nB�w\
�����:ӧ����6�ґ"����n��ٙ|�W��%^c�6_���|�CW���&w�f�3�(Ry;L�l�3�u�6�'����R���D��͟%�䣴��g�m�>>�RD<0H�~��\�s�.��K�H>u��4�;�Mrz(����{�61F�m��í��������!bQ7,���n=Ϭ����������ܕ�e�qO��E�AWW�am���p���7�d��i=֎X6��SH $�[�^��^�d�������!��2���]����l�G[�|"-���Ʊm�D�����G3��A��J�w���-�
Y!� pQ���Fݲ���5^���� D���d=`��xyU�Ƕ�dMVA�R������6�ֲ�'�����<g4�eݠ�6�̆�jE:0���C }J�#�j�!�kt����hz�[�f�Q��A
S�!"�	 4��t\:�y��u�Vυ��ށ����Ӗ�1�}����oYv���ک�E�2���@�r�tt	��C�i��z��i�}�3��
Pu>e���v�G��0��9�p�����b���R�>�"���'���=�{nf�6��*[��(�q��w`�}�8��#�$%y��=��Aֆd*� �0���c���cU����;�]����(� 5%q\���?�J<$�Uoϲ�����q�	�8��ǌ/e��b3�e�33JW��^��~k�/?��@��7�'��y�F���JF@�P��dx������-������ e2-�����V��>�g;����Y����VA�&~6�lT	�	�*$���Nod�`F��b{��!?]=�����B�m�����R-��D��G��aĆ:J����\���O��d�
麁<m��X�%[�2��%�ݗL��̌ �~����\rͺ���&�h{c�L�a"�h��;Z�{z��jf�n3YrS:p�N��Hx5O�񱼇I�:��u��^�YiKK��exF�THWҷ=(����D�R߿��������ו5ٞ�z5V[@�b.�y�G��Y���ZR�u(���e��[TL��'.�����C��TmA�K�W����c8�=����PO����^i�����^Ui��	�۱��e�I��Q��n.^�\�c�j,�Y��U�0|�D\Bvr����.�^��	����i�3$u $�{����V�'��@�F�( ��Ǟ0�j����t��>�s���LZ��_�@�����la:*VV���s5S8�����Rw� ��_2�\�\R��Y��*)�J���ɹg=�H�r\{�:�׆T	��
�R>W�=H��]BT,�`�3�|��k̼�捯V��)�m�����G�����^�ֹz��W\�u?o�����,�����.�-թ.:+�����/�64��`:й�Im��_���>yE���Ët� b��Kؤ��C?Ec5?5�����
n��_1�qCb����%�F��Ͻ�qx7��]��^�����f؆m�L�}��ʘw�)��g�ڌ���ݢ=��%���`ZG�O��t!tc� �9m�_�Kn��`O����~�S�h��Ԫ�﷿�ȂR�{<���:�m���u��$���	���Vd�M+,K�c<����~��+�j�T��d��c�@�oQ���h�:�-��+2D�\ȉ(H�>w!������/����BOMB��ٻM�M�mFpd�W�s��s2�e��H�AVe�Xm���������o|]=����m��U�t������e���g�~����fAl�Y� �Y��f���
(u�"��)R�{^|uKܧNp{ө����ߧx�^.M�;�"!ݩ�/��z� 	�4�ܛ��ŕ}$
q���@D&5T�\�ě9��������X|]�FXY���.W�'EƘ:�d���I�"�fϦ@Ǿ�U�����mҲTث6\jsdi�c����i�xd,�(- j�nqK#�N�� �דf �.UT����6�1j�ng5*�h'׮�g>��Kd�k��h�A/"@����KK:���_w@���]k����e�婣�^����>ұ��z���JmZ'�&��AT�a���Q�G�awS��c�R)��j�~4�������|ڬ����Ȍ�P4�W�d0�U�Ws;�X�y�U0GZa(��K�}�,�9o+��{��1Q�Û"�.�Ņ���E"g�m��@@�Q�eB���lIVwzN��V��(��C� �:��?X\T�%u`&��R���TO�e�#9����i~:o��4�p�2[-v Y)P�p���m����?�}�����K3g�zJ:9��|�}��8W�m��]�����Լ�O�xʥ��z��~9))q�8j�B�-�sϞ�o��9���Y�f���`	��܎+�s�����哈�� '���w��f�1�W��`��C�ً�L��*��=�s|3H���+��)B��|�%��ظ!���4���<������e(�<�.���|.��gxJ��[���6��byҁf�9Y��2���d,�1��bp����WY7�!]��hmG���R"G��q�T��K�<(]�r@Ed%>�T�h���f�u-q{�M7'��{��	D�hl�)%�Ҷ��5G."UpR�� ��A����#��+T��!E���.�͕b��~qr�t��ZWg�)�r�=H"��zЌi�Q�
����%��(�a����g��]5�PC�U1�'7�촔�@)IOpQ_I�$
'O��IN��hPkxJ���q�oVr��׌&�O��H�(�NR��GMֶ�		�F����dJh��3u($U��o�:5Q�����:@h���eZ�����mT�O��?�����)��z'%Ϟm��C��	�;�v�M����e�J0޲�u����P��巕O�7��W5"��*��kF.x�?g�NB'�)��$�`f{I�/���u;V�?M�*�xSA�jJ�#��P���L
������,��TR���ؾ��kU��ׅ�n�v&�j�G,{�²�HL�Д?:��3�%D� ��G�;(�#�e��ʒ��&Ԓ�&葉���b��R�<�+��y=��VPKܔ������Rl����S���CP�~Zr٦���wSB8�(��{|q���ѧ�Ta�~.iI�gH]���T��wyo��:�l�ύ�^�x�fe|L5�׆Lk�� +2H�%����r��%p����$�ؠa5{o��0���~ �w��%������Ffʗ��/��P#�����&�J�\�#y�V���I��ź�1��ec����?�#�	Jk1�5�6:�[��1�^�	]m��,.���	e���3~�w�13���۱��3�W����<��z��w���a����kɹ�V��A��8�shJ����k�4�Y�y�Al��~4?kl���륏a!S���k íQNΓ�Xu������{Q��]��I4ׯ%/�4��|�ui�B	?�<����WV�m�}+�VYǎ6'j˄��o�a�EB��
��Q�$��2�`9rz�2�Ш���{ƕ�l��_B-{3�ެݬ�dA�dL��u�Q~ͤ�3�ä��A�>^�gQPKH#��jJR&H)������wF��Xm$�wI�j%�_
84=��	�&��c�\�[z��Q�=r+`�)�~Dji�H��#��z���ʨH �nْu�Hl��e�*S@��c9��	�9���E6�M��H5�Y*���C��rҴ|u��Tr�|?�|oc�@���O��/|Ղ�|�Ai��(Ǒ�ˡ����������ʪ�"���Hn���_0`��E@���B�c� dC�Gh}ɇ�C
r�1�z
w����n$o�@9�Ҕ/�Gl,M��fB�4��� ��ݟ��@֩��dV�����yObcW��F=��i9{+�:mX�(� qŊF��]J��궳D�"�l%>��i\k�������ɬ��X�D�a`6l�e����Kt�m{��Y��_���������)��P�.�7��O��8���#;�-�Bi��yy�/�IWnm}N�-�RW5bt�s	��$�o�g^��{�*A�.C=�U�'%���V�Q�8��U���ڜ��<c������pj'tR8y�/��虣�|`B3��c1fK���?�9��Z�`5���y]�xA�����.��Vj�$��3D�J)u���K@��LSqQ�Fn�C�5��A�������(|��,uF�S�*۬k�&���s��ɛr��AuM,���L�@�~Y+�2ΠX�D�@w�]�]��r���׺�?:��j�ςR�X�SV�n|��o`��e\;^ߪ��4%"�n5�"`Z��2�ީmʰ�*3g��$�1��v�D����LQ'��"��\tۧ��;uي������}
�.[2���+���[5=�#�ؗ���L�BAz\Le�WZ�s�f����3���X��4��C��(/y���
N*�}�EH۴Yf'����"=��H�^��6ԁ"�D�c)�dH�+Qπ'y-JM �J��a-�)�����0�4o�^/�朴�֔6%o�m�TߐTsU�����g���+���G��B�(��f���'g���c�ꣵ�^mhN䌹������o���c����?�`G6(m���u��\���e���X1O�C<�!4��8.L#�NϫS.=�0�:��G����f��E94��jq�!����-{�����C��G�6����J�@��ܼ\"�J�2�7�D�)(�'e�qߔ�O��1h����C�OyH#
S��D)D�j��,����o����21��%ˮ\D~/-W\I�I}[ȝ���DX(�����\a�H�՛���hk]-��$��~��6.�U��NF� 6
���L�w7�Q$�1~U��#�� ��_*�n��[>�bUE*fyj����	41���ؽ�9���e���hv��ɽg���#>�-����nO�s�$1M	D��)qY58�����y�La���.��d���+��$��}�pap�&�~���~�i$�O̟Y+@�F�v3{L������ͨ������d�Wk.=�����yP謇*����#�z��@��G�  b�3˚R3
B�X�TӦp+�>��ބ��.�O�>z �3�E��� ���mb�X~��v��$E���X��ۛ��E)<���͂G8,�q4vih�ɤD���fJ"[�J��E)K�d��|��<m񢜚�`��OM��A��ț��e�`A�㡉Qv�����*�M}uFv9�#A���)ᷴc���i�B?𽬻���%��.�	�#q�f�&���/%�PI1T�b)���Uhg��엠͢��
}��ڄJ�}���晲��� *�3cճ=�dm�Hy� �����QQ�F�
�,�y�
dy'��?��wlf�!�3�������OE�Zx��}CP�J�l&���j?eQu�k�]E���y�.j�9�6�cI
�ȱ�[&�j���]�?`�\V9�xN��k�pjÌ������z�d��Q;��ʕ��J�7����\���O�&^�,-�P? {]~q��k��<ð=�g3YK�p�P�_*5�b��#bH������W&5�<Z�%{��X$�u�0-{���}���A���$�Fbx������y��ٔ�W�S�S�V5z��e��4{�i��{}1��Ռ���m��EieJ1~0"�*�83�N|����rW;G�4O���C�ĉ#;�:��<���%R�������@ 7af-ҖR>3�e�z'DK���rz ��An�fz�ή��������z*iD���v�ʞl�L�����ڦq���U�S\1q���=T�BwtG(�JjHI��şK���a��9sQI�g̪�L.��>;t��ё%�W���\b�]�]?%݉"^��li��?z�<���)�!�s����'
��94�v��z��ʮ�Y�tx�p�U,��_�pT;�ez�*���D�+,�jJk}ǭ�N�x��[�� �t�C!�D�.Mx�����҉��yJ��z�\=�(�n3E��Ē_D"��ELx��@NFcGH/P4�r�����]4i;����w[�|��LTm�^�f�vY����w�_��|˟��8L�2��`l
��2�qjqp�Ɗ��B������ )01�D�E�z5�/Hd�|
���|B��@������ݑU�/�G�ve��:��S��r��f&�l.�ua��e�x��_Ӧ�~��!��n���l��B8��.��݀l}��O���&�������Qo]&�7�d(�h9s�X ���=�t��CͮxQ����F�Y��T'��EK
Go�"�`S�	���ZP�+C~l� �%1Oxq�^�{?e0��D�,�)�n�4�[uoe�M3l�`(���κ��J�i�W�����d��>��N �4��)���#���3vXJ0�����C\�I�V�';A��7�3*�X�?���ʶ�Y*�q�\W��C�����Q�WF��@)��ӣ� ED�j{�o�,�������jʅ7A\���c�$M��"��0`�u�ה5�ǋ=7���!��ԗR��)ۨ���I���������"d�BIN�@o���ʵ��B0 �1���)��?��8�_G��īf!t�b_5��.�i������l:mU9(9,��:��[]�����^��]�ӓ�A�g�慰̫�y"�%�Z�T��p#A��>�u�XSZW�^`Mo�w��1F��A١��R6��T�D�.YoqN(� 6ہ��㑍�8)8��F��p�0��T�!�@h�����|u���`Z����zv�[��L�H��0��*)nAv��l8���Y�A�i�[o�cs��ú��r�z��Q�Z�n�J`٨Ќ�u}�G����������#�;"9�м�r>�H�>o���e(>I��wq�ʴ��ơ�3��A������7>.�d8�t�����3�^�ܩ�h�;�J��L<?��+0x�֛Uϑ����T}V�5:����{Sb�	i����۾t�ꁞ+Gv�aFc��z��[�ػ*��ɱ����Ԇ��`�6�r^:(�V��q)�u���؄8s��ֈ9����9��f}�	cƧJVp�����0ܶ�������x r��s&��6y�o\��6�-y����w������]t{�o�����~�x��2��BeC�*,7tC�C�?J�+O}�O�o #�Ӕ��=\�\H���Qc����.��p�I䛅my��p��RD�@?�μ����l[Y,�ߙW�b0�@2�Pr�y��{��w���{��˴e.�G�K�G��hc)/"ط�pT]˾����)��]�2ǌ{.0�]���SC0!��lh�n��|�PQ�N�I�z�Q�Q��`��h���p�3LDB�Y��~���V�z����*?e��`��g��]Ǽ	�VȀ����T����3�q��߮��C7�@����
m�Z�Cք�̊��4ˡ�dO�N6O�w�F��̇�q����?����7�7�D\+jK�R#�Xu`�ݰ)6B�N�̷�:UyZ����5��B����]D�d�ے�X�$��K`ߗ�7o[���?��R2�~�>�۰Ox��皧�b���7'ˌ���);�$�v��i�+)
m�H��QO�ƹ dv7�g �uhD���s�9��B[Y�@ǔ7m�n�}Ș�m�3��>,bZ�gv�I��1Ln�LsP����jGx}��t���̑YlJ����bط|^~j��-zp^�o�>W���4��ڢWH��vz��v�2���L=�g��8����1�
~��(����+����3xEYk�5�k����Q�����=��DG��<��:���,�<�]����q1�<B:�N��w�p�>S[��\����1�"�JO��j�Q���k�:0�)p��g��0ş�F	�譟&�r��2I�D�����#����������C0�8_:����Nǒr͠�O:�n�=��b�����NKX���I'����R�:���;�_��*c�A�(�����>8�P�蝍�\���.ʕ�t�k�4�~J�b��MP��N�Ms0/��TGx �LIʢ�#m�L��ڤ�e�T]��E����f�Ho��m5��w��LH��-4~7���P�����c*�v��˷AN)N�ja�p~��`@�����6�eq��l�K��	�[���wȞ��E����'�]#E '�y?O'"�m�gx.�~G�o����w���q�q���\1�7(�	ld�	<��uV�e���Z�/��󾂫S����LKJ�<�Q����:����#�ZB�BQ���[��H�z��Aj�\��i~h��߉���p-�&���>+�&���Ųx��7�Bc�"N�@��*�/07*��R6����	�o�����z��u\#���b�}�����8#�ʨy��$}�+?�y�O������,+_.������2�m���Tu���Q�@0���O�!Si�$��ټg�ZO^Ѽ�#z�b��`�t��SI�X ��{�T�cN����~�S7z�z�R��x�8n��Nm�=pM�+�ix�Ȗ��e��q�\�~(�/�J�7�R"�*kd�{V�g�{Gf���f燣��6�r�<�ɿ�U"�F>�'4���NRƙV��%����(o��N�O,���yOX^�a�Վ"d�YK��-�)�{�cC*��h���d�sY_��H"k� n�����i��>-���VҵCBԈ�T���"���[@����-eB�G���O�1%�@8#/��#��;�Uc�n�+y�}�K��mĂ��Lȯ�r�C��)��#����`�F��~xk��h��^�㸯J�u�˸f�#aV9 �e7�o�I ����I��G�u�&ܩU~&�*b�˟�Uᒝ{�tgp~����j��3J��؝�1���7Иu��N��ug��:c�:*:����@�'��	�.��# ������k$��T������N"r%f�����b1_�F6|��w�]�Ep);p�(�jsc�j����d2�W-#
�r���o���Ryw��^� ���+�]A���V���G=���gކC�>�V1����ܫV�岣D�h�Z�<S!8��w���9�"G�Gqx�`�����vi��1��ac�D	T.��JT	�`D���gb�R\���4�O���:�SV����(r�a$��!�7�*.Gʟ�X��l�='���׃��=d���MK�G�.�
])~/�G�Ǎ��4ߵ^��N6�Js1p��H�@�%j��������� ��z��ǯB��R�g9�䭃��(8�E/z�G��ɩm	�)����N<eܣs��{R!鋪�5k�<\�}�w�B/!(hƋl�|g+�|C�. ����F�f�Z�>�7��U�PqxB܌�ƹ��@3i�Ɏ6��?	�_;��)�q�G��p*�(Zf|���-|>Xӯ���Yi�h��xX���q���k��g>�Mt��IMw"�¡餝���ĩ_�^.Dڕ9yο�X��`
�~/䮿L�C4�JwK������}:�"���*���>����^��P��+�ū��/Lkr�����a�ӑW0��ުo� ZbSX����Bp��T���_t�d� �]�<b9����/���k��q���*�c/��8��ֳpGa�~�Y�&��֬r,m�2~�`�;$'yZ�����!P�������:�:�'�.X_�l�vPg��������S�ə-X�Uahލ`�n ^V˾9@�U.����96zAz=��>9�j��Ey�/��i��ej�Q(�*�k���D�K��X�H�p�<b��w�B\?׼B��k%�l�)���t%��5l?	�q+��zC���ҽ����7�ҧ����^
mޤ`�}�K8iY�.tgq ������#�u&��G�{��@������hkq�����%V#�z�s�%-F��"��o*:�۶�W��� ����"�{0�*�/a�cn��Ѿ�cڰ��Üf*]Y��-6!k|B���^�Y��6ok*��l�(�%,\:�B�� |?>+��𨉉�R��{��P�pa�z��k�=�Q��Ƭ-t;�E;Y�{��?#f0�ۜ{��_o/}ƹ�aTd99�}��ɺ�(
�������6H�LX�{O|T�R��F�}0�j�Jae�vî���������a��[��8�gֿ���j�H��e�?VU����,"{9��E��U�ԩ���M�
�JX�NzC�o���*/G&o[�����Ş#��Ĺnt�2�>J��|k��r1��8b)s,�\Z�W�����P�cS�:��:3bI��zh}�F��);"������@iz��@�p��$�{�3�[�fn��˽I���~D�c}���K���Q դ��(����U�������!L���_�2�zį�l~�<��7r��/1+2�|��Pjϋ���F=
d��&El��ԄFx�?W�y/uDJ��=�ʔ-�JA�A����F�[��%:ܑ��H��'W�$N�V]���2��6.���J�]�`�_�%ʳ{�����5�������0��(�Q٪0�i2�|8��ª�,�0�m��$����ܥu����Ƚ�h���s\���13�(����-3����g��X�R����Y���'V��p �����*2���$�Ԗ/��M�M�Ѥ;��V���B�ڸ̿�c�!�� �V�Ď8g�8��Ko�5-`	���ף:�_dr'��xx�6,	&pd��P�˄N�#A���SF�Uc�t=�겾���m�4����gd�'/�)�5�2��=N}#7F\Y���x&P���:��$�ia����|V@����1�SwD�o	�3!�.O���s=;�ģGa�\Z:~D�3 0��sI,�@��B�r����(-ʏ2y!��w������4?����ұ���F��L�Wh�6`��ۈ��^�b�[���>����n��E�&�Ӣ�Uj�x����+Ļ&��~k�&���nҬ�9?��q�G2Ax�Y��u^o4�>��OM��f�ԏ
��}x���@i����9���zy�DYcK�]-d6}�x:�zD�-X͚�kJ-J(ӛ/<��������A��D�{@b!�W���AQ�U%+Q)�IR��,o���'h�;��2��à�!S��=�$ڕܟT�g�(@v�zR.*�Һ���4c�[���#W�
'�n�f/����<��h�oE�lʠ�o�&)�aa3E[��ؒ6�<�)�V,�C0���j�hL˳� z5����~�Xz+�E�Ŵ kcfb�&���o!8#m�}K��3��!.>s&�)�$��?�X8bCv�m������:��T�:,��n_��Z��t)�:.mG-�V��⃓��r�<����.y���9+���t�"����\�u�_f���D;���9S|������}6m��(a���x��цڐc_7y�A洡�����]�)�<�Yȑ�.ª���=h�5!mX�PD�l~ �ad{���'�{������ ,��W�4z�~���(��2\j�ͫ�%��T�k�S����ZN�����HD�3���}	w������ՄQ�/������;�'����ɖo
��X�=p��1�L9de+�Q�`ǘݽ54�_�
X�o��Bܴ�N��E��Z5 3M�K�k��A����E����:��He�t��|"s�8��8�nB�){G���U�Qit\��k��v;$���2;�l�_ba��q����֞n>:/�EcW-�Ԉ��DA�;[��b픻�U0�A���g�z��>��P���a	JCq#)w��.G���.=51,$�H8��F�{���nA�&��y'���l8�^D�)���C�����u{u��j����et��2�T�1����M��n�;a��R(�����\ɱs�"��n ��9�tuZ#(�/�%���vv�-hN���X�`K��S���jo�䯯u˦LB����h뫪����)q}:�'�%�g=��O��{:g��<!قM�Aoj��sI�Qr�qq�c�^�fjow~���֯k�T�{K�l��^{ϔ?����Ч�w+)q%�̜z���8�$Q�B�
��ץ!��r�������F��o�;��_$��4��_����Mow�J�-���\�۷-�]�g ���I8�/���T��_R J⳹�F��`1>��{~�Mw>Z�lC��a?���·���ә�,� #���q.nӲ�_���8�a�Δ�;���F�QR�eN�����z]J�OE$�7����Ѩ�K�������;�ff�N�q�wyo�S�d,�e��i۹����+"�GE,�#Y���)��7����<�5v���*�8�� ��X-#��S-o�����5�Ƥ�=��48D�D����UE(>�[�-�	�\��B�h�βq�@�4��L��u��W�ΔǬZ归2��B���Bs���'Z|&Q�F}Q�wyJ�N�vη^��vP{��a���~�?&7��� ���\����� ȩ�4�XG|ޭ�Z\��eޒ]��<jk�B�t{�+�L�����Bs��舽��-�~�Pl��?Yp�,+U�wG�[��<�[��Z7���zO]�區��a���A�\E2xUS�v������^U��)���^'�'$��V`�m�0�H��om���r�m�[��v��D��vP}-z i����^Ii��3\|<�J��^P\,��w����n�sP�,]�w#��%�����\\p2EY�������:s-u��mA15���X`�Zτ���:L_��k䭰�M|�4w�[�S���z���]���}�ʙE��ɲz�]�歽�ޫev؍�� �A$�n4x��bR��2� ���޾�&���ȹ, #�[���eż�-��X���>�=y��j�k�cP<����v��KL/�y O��pZPQh @.Y��b8� ���ߙ��
W��2�mlz����ҥ��\I�˗���`Nv�<U'<*�t�]"��]��T��~v�}� �q�5C!��,��0)AE�V�{���3``����N� \�w���;�b#ʹS��lі��=J5F�)6R�t>�-�؜H�fIFK�����3���'��x�|��i��%)�!�pX��먷Mn���e�~Zm�\��G�d%�(��X6�b�l��CF�+��;˒��\�������z�E�.�Z�A�s�\���L,!9�2��L����bӺ0�t-=��j��:���2`�7w�4fx`���R��ٶ&���0�0���*w�J�1�VT��@��vr�ZL����h�&C^��ˑ�&���GF;n��T	7����%�)��V}������"Daury���R����������e/bL�$��#i�=�%�D�!ˡ_�sYL<#3c���LM�e,�'�k�D�?6�$E�K��*��D�(gu&�Z���a�(��Ǒ�����Ln)Z�(��]T_y�F?�.���|��5uE|�Yp��3�l)�L3N �8��r���$ʜ��v���5$��A��"�}O�t��<Ԫ�j�*&@��_�.z7.�Z��J�d��!�,�'��d>�4�����A��D�W$d��<6�Y`2ٹa�������8�)t�Ād�ip�n3\�a�3Y<`a�#x/l�r*l�^ppM�6j�8��5o��pN�@�#�y^u� ����Q��?<o���EU�N�)_y�f4�I�)��V-%$^��43DuJA_s7��q���j��k�o���9��, ȅ O�e�jY�y+}<Xd(X�P�C���ba�V#Z�R��.ik��P�.Q�*C�⯂��y�`�ʥr����|��fE��tP��0�N���[F�_���:�q0ۍX�m��{��Y�����Đ����c�])u�$�s���N�C@{�)��e���4$����Gq�^���,�u�Ʊkyq�dJ�e+���gƇ/0�7$ ��U�X����x/��5aI똦����fْa���V�5 2�=/��}���ߝ!�G8I������񞊍��e���~�
��fr�$ݨ��p,L����d��#�8��8���J�q�04�~����u���[f�����z���C��1N+h�X��"(䘣�YԢ���:���asz���~'ǅ�Q޴0,T8�%�S�s#c��Y&�z��J��z3;ƭ�@��?����a , ���&É�^���l4����d��C���s�^�<5�=Zt^�\�?#ȳ�E���6�a��0Y
�}���W��p���C�-(�}�\�J̡+��u�
}�H��i�������#S��Ə��+���;e��Sg���t&--�^�
ey�^�5Ѓ��bT��a6�5B���4�s1/0%o��&�g�քWJ�B�ΝA#<�)�fž/a�Y�����ĶD>���-�ƃ���;��")����`9t��".�}pC��OO���>���ޡ�"�X�B���Dh��Z�����3�$�<����k	̰��L��Z1E,�����/��� ������Xo�x�$���s��%������TeW�#l �� ��PL�M�����X��?����^k_,ۢ-	�%=�5P���=)Κ�t�44ݾ���tdKD̯g[���>�c�N0���M�f�x�V�����<[�9��@�1�-#�'�C���GQ�k�����
r�qsw��2��mY���WB��[+�'��N1�
M�O�O����+��?�]�P�Q��tF8"�� ������P�Y���$�j���ܣс�B��UIɹ�v���v�ࣨ�{H!\���aW�#�f�l3`��T�|�\uV$�9N<Vܘg��A��c7@�M�}�2��d8����@�[�"�Š������R#��I�	me�?Uw��t ���\%�T`��Ĺű"-�E�.���`�VR�eik�V_	y���ka��7F�2�%���4�
9{��C���j6g�3�f�O./����I���Q�`Q~�p�ejlܛztHɻ%ZÌrF! Q����O��<���ǂ���4�{�h �.)����"��U�~�z�6?`bK-�Z	�LS��9�,���湑���>ջ[���X���|�"w$q�4bPdU%dw{�= �D�0b%�5%ߝz�f�zFv�/�]��I� ��`ٸ�h����y&X�<e� ������� R���y=(V� �ثhM��j�����B��c�$��%�V��)b|��J*�zs"J�����b	�]oս:t�nK�Jߪ�P^_Qm�m�^~hU�$%��cf�^f2�~�0*��藆+���V�:#�S�-e�jh)ԆcՌ�p%�?�wއ&R�[��G�4�wR�\�s��8=�n������������L7� 6�%dK�A�]��Y)�k��;�WҺ��~A!�����ǯ��+e���_SK<]
�o��lC�?�8��~��&SS0�;�DV� ��g�(.Y{f�,�1��)�$/��w�|i#'�S�*n��PpB)T�3�����%��U�=Q;��7+�M��R@�w[�����kv�cgE�@��w��͑.����~ �h�}����W1� ܾ�M06m?Ʌ�c��Tj�c�3!x�S-J�ڙ:�����?�<�>�fT��}IR���y�P]��x�}ˡ+��}�Y=r� &����k����,�x�kg6��5i��闐Ph�p�G �o�q<;�k��o������'��d�7)C̋^}��8:���,�i�7��!+��)ݟ>~�����Q^����Y��"N��V�	��,���b8/r��`�;P�5Z<��Fր-�P���kN�Vctk� �O����ah6iy���=�NB#��z�����c佥8���lPXn��} �R��}+�H�R�.g{t_�C1��m?M*�N�u�9�G���T��GaD�D�a�xG�&��f(�S��@'�Y��e���2�@�� �Q� ?�z[�>�S���E��9G��5���%TUre���(hM�k�l|5�ic�h܅ex{�ig���P7�����_��e�~1��,��7�mw[�,�T7BÅ����
9���
nv0[�ehM�	����'���	:��Rƫ��o�]Ax�^j�6*7���X�≊��莇����UO*A�rc3��9]�7s�v��M�F7����b��J(�g~�PG4�+�DPE��$�{�zMY��*�U5o�r`M�׶ٞ]����(`z"cN��  �x�Ǝ!�������xzIL��Ҵ����w����%��Q�?���V�?�>���u�<U�t���I�f��Q�%%����J�
i��'B� c��2�ֿ�<T3�b4p�Օ��H��a�O��I�������ǭ�ڑ�z�f3����h�s��Bt\�zn��qLؿQՊ�^�Z<c}�ߐ6PpS��B^Uj��[*Z.�e��_�Ͷ��Nt��*����t�?�O�sʕ�,������u�7��ȠYi�jX�w�S�ӤH�*�j�lB��±��!.~�>�w=Q?:����[j� ������rc�t��v�]�OXΕ rj�4S��u�K�CA���R���Ʌen�>qu����#a;�(�bٟ��pUM�ɺ������!��m�P�i��(��Y�!����M�q��"��=�P���%�����U$���[K��Y�adP���Z���ѓ��M��&�3���lM���m���ĵNG^)�Is8�^L�s�<�YE�B.ݲ��1�`�y�fY�ܿ��p����$��\0�l%j�b�mp�l�[D<z ��iz�����o��7#��r�i4�J,d/�|���B�
�|\���)Dv>�^r�/˗n�)ݝ�8��}����u�G��P�!L}�v6�f��F���/�q���>6Ϋ�-�b_y���c|���h��md���[��&��/��Xt������H���\�8w�v�e� �B�t���u"F�Z�G+1�3���mx�J�	���[S?W�c^c`�O"LH+�1��|F�̯{\��C���d��ۣ��Q��9`� ���?�؍uaE������\r1VG��+	w�us�ԥ�ML\X�í�w�������	Q�9n=����i��]V^�����q�(9��I�t�r�gu���]F#��F,M|��ZQ��w���^|��@�L�M>����a���y�y���Z�W��d}�PM�҂aaAV��Vy����)�r�s���"&�����
֡y���M9������KF���E��PpJܒ���P�O�9�\Ɩ@�cm��~)"��TG�q�R�����^i��^h4s��D�J!����S��P|���j���w�^�9�<�3�N1��k:��K�N	.ޤ�����Qͩ��s�=�N'�_�f�ޞbT,�0+<?���G���
���#�r+�e:��=ݚ}EFV>l�i@�AV�tW���_{G&*�K%\����#��SĀl��DG��i��E��ǋI�9�Xx�����w�i������xBĐ^�n'~�#���Z�����}�����+�q��Fp~�@��I����#��]�8������k-`�0���X�c��H}i,��7Ω�"�a�u��B���趄��\�'#37'���j֧��f�yN����_N�yn#����@��zܾߌq߬F�(B�cO���"�3�38�U�B��,������Boց�����xM�a a�2 I��X�)�R��<wǾ�XtL(�8↵�ڨ�$;��e��'�,S�B����}���?��L[���Jr�D�[�qCrW�ۂ�=���WY��������C=� 	�ߣ��*����5m�̹�"x�y�\[�w�e�P.U\X0�]Z07&̢AiY�[�E���Z�V�2��zGB��2�Ŷ�*�^�=Z�+|�)I+����'y�^g�HX���a��Y˲+u浂�$�xT�k�ҿ��g6��z��Q�i���g���Z=�mM{�Il)�j�<(���)�u]�'XO�ϩ����������x���V;�P^r0<�� �P��{�����~m�4�c�۫�OwnVg�RO$n�l� �+��~"I#7*�u�Y�K�^�K���[f/��A49��� `��a�vyB�x��2zA�9$nܣ�-�C��]�a،Ta���0M���Rp�1�gڌ�\�_��y�姚����U:�)�l��"��|�?�Z�~�R��pU
��A�*6�!��@����0Y������A�R�i��/���h}�"���5�5�K�sd�F)�w��0�%*��w:��C sO�Y��J��i���,��%?Z��SaO�A�o֌n��"[Bˌ�h1Я�X.´z٠��Ǌ2G,#����:� LA�Yr��Խ�� ���ӈ)ͷ����OQ9J��l�.V3�������sǮ��x���ן�'=96��-��0�L{&�ǡy t�vOr������`��+�喹(�SV�(B�h��a}�Y)R��8�b�>8��}��zw��N���\�)ΛJ��1r?0r��xOM�=-θq��7իTQ���C���/N�*K�E*X^8r4���M�2�������;�kc�(@�k�!]]w!^C��`{N�^�+��&sh���b+��}i������#�X�l�C�~��wj�1��C�D����su/���|�D�s��Z��9W�$C�� ������ ��
}_ox<���"�L��mr��N����E�a���Ü|���'�Ans;�x�)Ex�]�_�xH��I<3�0����B0��Z2��ɽ������u?�%��ׇeG�����n �L���h�vV'v�p��r��N<�B��N��h;X��z�yu��2��j����٤���c�8��X���E랁��=�����¢l�Dv���8=ƝH$�F���P~��P�͖����/�Djm�I�-�0J^�I��j)�4��>EAg����v��vZZ��Ť[��Փ�:JM;c��m	�誌��`s�nk�&y��7S\��0��&��j
��V(������2|f��wT��b���쇔԰rG�b ��ݛ�ހ�I������C�G��3^�����?���ϥb���-(
(��v�+.�ͯ��(�9w�K�����4ʶ�A3�T����hY�\�U��\�i�J�cey��K^:�_��b��%�7���*ˠ�܂�b��F��M���@����x���]���������M'E8�P�-��M�<]=�ly0�0-zL��:`|����-Tv-�C��(p�����-�2a�"}��ꌋ/u'
�C��իP��W�N��q<Hv�i���uӹ7@:�C ��$ҏ��H�4
PhBoF��ŉ;����!^O\\��@�� *�RI8����T���r�$$����~�hn�W�9o�(_G6XIп�4޲��T>��h|�i�S��1"<]\���K���tc����Vֽ~[	�ʱ��'�,!8|ʇi��0ܶs�O��H�ٸ�ҴK���%�l�a{�������}p�x�`���壵�`6��M1a���h����|:���õ�wpmT=]q�����D5�� �����wa����đ��'c%�X�5�<��.G�)!W����OK���T�`%N��.�Q���jO}�f1�����ӆI�ہn[
�/G�f�!Xo�Gd}�ZZze����b+�;��D�4�"�-�47��X)4��q$�_}i�+�49~4ز�D�h�$m�.����?N
�阱�"Z��5���CؗjF�N�����5q�k�O�֒�����8��/\z�:�2���r�Ns��M�hJ��9��>��XbwIB��#o�ʳo��N�n�y���TE��DJ��}	Н�U9�H�@��_��6X�$0KW|��H=C�9F�o�=)�w�Ll�T�kO�^�@U��b����
.:�G6�H�Qw�K'��f�CS����;H��I�A��Y��Wk����.�z���Q N�x�:?�Q��RSWE%�D1��!�cp���tD����"����ǂ/��w�g�w:��zT�$�>_���"N��gU�'��Y�S��$����']�Fv�/��}\�m_�S�����1�J�����|��K�(/O�D�m��������nW��kq��.�P���U4�X�x�u�s��FNG�3�^��}��K�m!0����ƍ�YX���Xv���[|Cr��S���XO,@&�@�H:�|ůś���"�;��z�r"b��>p{Ⱥ�tRU�^��y^i+`
��w��s/ZtWBm�5'����GН�����0��A��d���^��=?��.d�8p~��Qp�k6�Ym�\U}ӑ��}�&�As��nR�uܩ-��ߑ=&�X�r�J��L/�Dg�)*I{��P��N�{No��y&�1E�o�&�a�+Wv̥\��ٵ��w.6�#�^�q�FϷČƚ�wWj3#�@�c��A��o�!w��쭇 ���3�;�Yvt�C�,ϟ[y��|&����VIE~lyfr�E\��]��TQ跟L6���$73��ø�bo��)^�l������~�Ȩ\�?𶧫�8�~���ۆP�Ws��\�&	��r�� ��Ө#�]q�bL�;���Q(2����2>&ި��H�|��\n��\(�D�GV�` *e�E���,��D��wJor$^EBRBG�ӫ訩Ԋ�J��Axc�F<:�W3�/?���0׵}�0?��cZ�}G͈�.�E�u���(*�5Pj��Av��4C�),�L�Y�\9�c����ma��|ir�x5f��b��gVZy�U�2mDe[xz��sdS���'\{�s��E��l�X��q�E9}�t��Z���=�[@p�_�#��v=x���%v���&�*��F�Ւ{�2B��s$�xvoz�� �54��5��4�QRqIͨ\��n��!�+I�	�2BLV���F�'���T�z�3���͌�S��N0$�E��2uH���a�2%b��)ӷ|u�����{���DP�9�gn��J)Õk6M�JK������ņ����uO������^ݷb�Ims��{SB��/@@h��_ߜ�Ǘ�Z	܋�Pɡ;e�9Y- �����Z�Z��o!���.�wC��GLˠc��a�<L>�{W�8q�J�Φɉ/��Y��^��3�ԝ�y'J������Ԭ��K��S�^�>o&QƠ�%�.L3�PH�x")h�r�Fqj�Y����bڃ{ɦ��IA?� [c&����?*\<J̛�.��/�n�Պ,�H�X�Ͷ4@��6]u�q����Hl���l����)�{����Ė&��:OV�wJ��Ѕ��N�So�Q/O=���;����,�!t��oD`�|xz����rnC�
�K��,�LΉz������r>��@��� � w�i��E(g~��ջ�?e��ŀ�����ő�B���#ϹL��ˎhԒ�]�v�k�N�{ފ1f�TozVXٯ�IG�������!o���:Yc��`/=�F8
҇�[/��w�Es�T�E[In��P!��͢�,�c!Ԁ0p�<������ǔ{��8p�4�f
�x���7v>Q�����Amz�<_CCȊ{<'���-����5�.m�j�Sk���T9_/���b�zJ�h��S)^��t{a�/����dV1ɋ�IM�%�	��k=�jrw�=8cUI��~���2����Q_N����6��E�{��o�r}�P$%��l|�G��0����c8t�-�>���:�%_��c�ŕ���E�#-�����P��9�g���M�wO}c�T��1�4;�s
��KV�MU���.�'YX���gTɚg�F�'�4��dHP��P��w��c��9��6s942\>����'Xk�y�k��x�]��Q��c�#b&� ����o�&ֹ|�N2���9^��DV�N&�Ѯ�����=+�!���� �ugGg�}@���g�ᚨ��7�s6��r��oe1�k9�t4c7O�ʪ�����xe�$�-����`�9?ܭ�-
=	O��D�i��2��tx�O|�����j�����0��_їU,A^�DHC�y�|dxZ*m�~e:ݐ�_�'�j�]y�P��DO������O���{YE����y������J�_<��@0�B�
j2��0�n{_���;rQ�Hn�'��n��f� O:"�"��
�L�Z��D(��2�/8�O���7�n��U�G������_�QaN4ޫ�`��֋��v��� ������Ab:��k�Yn����%.!����k��ow�c����7���C���6�Q sMe��є�>@�7�!`��\�.;��N�� o��\�۲$��/7a����0�Q|av�	.�d���7��A�1��4j�'�!�$r�ÆQ"w}���FC��G_�����;1�P�	���E�ފz8ռ]63�$ �SJ⵭�{�O��Z�����J��#�D~�� ��o�l�O�Q+_]P=tĞq���I�:�l/KM=}KY��|�fG�2}
��Q�V���|Z+/��^�S|ԁ�)�z�K�0���x�Ջa9�W�Ç-��(�kt�/��y�UO9������N��W�t�.��]�������z[Ȱ��шΗ�����y�ۏ̟��r2n3�PZ/5＀+)}��h�gh��E;�}�����R�$	[����#�v�-�܁��*��Ihx�2V��~֪�}n�(~R��l$*����s��(_����󌅫��`t��z7��56h�'zH����x@�ͳ�wl������l<���x�#�㙼	�/n���!����#�>��� �{Her��9
���l�У��8wv���-�ZQ���-�� my��I��_�8ӌu8�&�a8a:��ĝ�著!�\�P�0��I�A�rS�/�4�g�@����b�K��b����1X!�f��X
��t�˻�݋-��.y�1P��HG���٘Qn�~[��ި�!%� ���VNE�y��\���<V(�C��#Q�Fi�21L$��!`�ەջ����� �������r��N��fZ�|Ƴ�Z���y��b���9I� I��t�ճ
�ރn�X�A�ܤ�ߑ�Lx˺��ʠc;�^2�L��3���kI�e�w�b[��H�]o��rT�e�
D�Ks����um��7���R�Uu����E�dR���	�,�o[I�i�C���+��z�C�з�d�c��7��Y\�T�y���*E����Ii�3{��*�k�]�
g~&�.A���&�M��+�O����P'����qC8<��M`Ƙ�4�]Q&~&>��&b�r]�*|��H�Y1�88�<��%�m���IZ����k,M �e3�.��;A��^����90}',�g��^���� 2�4�����o�4��Y�S������=V�8|M�2�������_:�|al�4�=�^�)�Z,;�����������#٘v�.��a�٥�B�8?��!Y����W db8���8V2T/dJTV�������Fs��,I&D�=�i�G�w�*U��^\����E�W!M��"� �f���i��E;Z���d��4]�	�G��`^2Q�8��o�:̦wiƅ��$�*tx \O��R�B�pp2�H�bO�Lr�64���Gƴf%�WE3N��u�Y���a�z���<v�LѠ�"����0P(�oF�h���s�Z׶N~��Y$��� jV��_���V�&J���:�)xl��
_-���P9�kǥL����u{(c=��h�Ԑ�|urc"�J�+,�<jqi xTLA��wY'Ԣ=/�v���*��F�B`�J'�{��U��@����xH�h��͆ڌ��!N�dA�Vu/K���N�Y��T�@J�^��/�³.|ð�l'D<��I�&�0�7�SшT���FG����l�X�!�� dw�/je��Da�@��p&��o����@��ِb1\$^��za�ֆ��V�[�x2B�"�q��"�@����c֡��y18�΄l����dU���Y��2e�o�h����.k�z��:�A�-W���w�{\��g� \�Y"T�j������zk���&���*e�9
x�f_ԉ�R���ϱo���-�������k=o#P��
dZ*��d6��	?�@>m�-�>�׌f^+r"�J��Z���Sܶ~xƭ����J��w��T�����P�G�tq�F�xA �!�r�&/��7��L'@���L�t��^:�^�[��g����"2�|��<$Y���G�oq-sM�/����3D��}FƗ�Fӆ����6��'�m���.z?\�_����J{�)���V���&���`�H�ٽ4�e��j�V���T"��R���8a�w���,@9��͝3ƌ�~fߊ-�HU����qSPjԪ)��@�kY��J|���SzL�)#�ɃN;�S�am:\�&<�|ɵO��O��:���Nʪ���DP��.Dx$L/���l��������Q,��[����Y'R)�:8Q��GA���:�bi�
�x�ȼ�ՏH�oV������7�˓�QB#�i�@���֚�����|�u�#�ʉמ�dK+�����|��N���AC0`S	,�A��s��-0��q���m����J���$��ƞ�+���������ҡУ�פ��J��J'�~�w�%k!��+쐭G�Qf�g���j�^�A��NK3�H��_�/}���O�0�`�7�D���p<I���b�5���ٱ�U8V�b+���k��d��SLֽǂ�^�uuy%���Q�Ù8
�k2�q}Vlm�P���tF|�Y{��*�.cU���Q�$����j�A�]��fP��H���spk�:4���Ø�
��Qf���7[�X���S>���iN�v�g�0E�� 2�5�fe��	i�d���n��0�I$?��0&h�X�x/�`Z�H�+t:�E^�ޏ� ��\k�-ҵ�,V��yYS�Fm�w�>�nI��=�㜨)��4E�DUV&��y4x�}�7R.;	�=�q3�&���_����^f
�K�p4�5O�p:e��������Mn$=�I%<��]}���t\t5�z��Y���I�R|ʘ�I�P�����BH�!�:iY�0Jv,��=(T��r~s��i3��@��i@M̛\!Pw<
Y�G��� ����!�i�/{�&~)������[��8.������p'��:q0� W�����S�O/��Pm� �ݢ�i�G�J��p��4�M�EDwm����Bhw�}��"�Xk:h!�;X�n��A��]���TN����N$�b��=<'��.�����=��>,W�2O���'	������Wr�����	ۡ��|�U�8N��k�
wU �����T�u�5�h����-��x���d�h��������3�s��^qW�zRTf3�a�ҧ�JtzC�}z�0�e띾Y�.6�i�Ӄ�2�-�՜��>�)�Q%o;��1d�9��GB��ʵl8u���PS6,}EC��n�I�w��z�NP�9*���#i1��}����R�����'���#F<���lB۲�g!���Ǹ�3�:N�nG^���y�G���q}�-�K@o��:L���C]�:�V�o�-'8�2�l��`.�-hHˮƗ-���h�>��a�Z�y�`�1������I端����P�&N���S�IzV�����7���gU.�ՌoKj�,F��yH��{��� ��������O����;��Vx=;\Gܽs���r�>��|å��_ �Y,#�
�	o���<}w�d�]1��t�0bD �ܩ��XnJ(�{K���w���*�%Rv蕩4ar�<�ʁ|�E�CQ�U6�iA��m"h�k`#�31s{]l��%7[��e,��R��X+�
h7��i78_�!���eN���]���T�Vb�Qb|��f��J�6{�ם Qz���;�xL�sx�q7Rvq�6�_������v>�Z��p�{�]�.ac �Ε�5��|������ �bM�6�u|�ڸA��>4�$}Y�e�3h�kכ��{����WZ����7� eվB�������L��W���i�������T�~9�â/��c�6��@�$xR�\�G��̆TM���hL�����T����Y���Ϝ]'���҆�v��>�xM�_�»F�֍�1A�T)�{=�H��2�%-�����hn$Q"����U,G�]l��ɒ{�ӯ�߼ïU��5�U��{�+�Jz>\H�ͨp2������#���IRMެQ�+�c�Lb�.PB]�ta\1~!�m/�uo�-���E�]ݘ��U��,yT3��ό�����V"+�+/�(��%n�G]%���,�2C!Z�Z�kB�5�
?�疫֨i���P���.c�k x����̴c< ƼU��n�����oL�z㳍$?�^�dܧy\�[>�dy&�h��&���ͪ2F3|n�� �W�d���󔌟��5�hN֠��!�ٛU�uл6�G��kbG����79��_�Dĳ�G7�%�Q�K����-��������yU��jn�6���Jr�"J�(��\��?'J����n���!x������u�p[D�-M�
��>'8*,4�/lmG�\��i�2�FC��V�gG���i5}��Z|��S
g`�,��:O��~[J8j��b��i2D���W�����҈��8�s c%�W��Z�QoG���"�;�b\S�J��ڊ@f�M��ԇG����X���k��� w��Q���V���/��c�κ1M|hՆN��b퍡nsVm�H�^��Q[ )}�±7E�h���E.��`�����aw[CT�Z:����j���y��!�N�]`&��`5 �\�!w���ڔ�voB����N�
�ɮ��QQo�o�{�}�(�0���P�%��I��Z副�X�%���J���Lu�Lk�e�T1�ܧ~2��V�ZO��Sm���R_����%�~ c�Qpf����4�9�x��R��뢣N�?4��Uߝ��ww_X�aKY˧i�s�X��od���Q�e
������jZ�?���l���	*ٜ�4�lA�]1�q�A;���%|���Q^~�CYw"���;���G3@(ۗ�4Oآ�H-Al���Bf3���Di��D���GK�"���kfzy-r�������:�7�!���y�&g���E��z?w��W7m�X-�&�S4��]
��)���F��^Y��ߴdG��ޝ�Q:���Ε%Q�� oj�5y���(��>��.D���>2����r�/S2�ѩ>������B�_A�0p��`���o9�oszv;����eG��Ș?�x��Ǩ�8����a�'P�����d�
U���6?�uWCƸ���LY��Jp��=R���^"�( ���pЇ��:�=Y��b�R)���q����tQ��c�%ߜ���X9����۩>W8���G�^2?����k��B�-�����~t͏j�:�jC��;xaf%���'8�zX�zo�m��rEk�"���?��.b���r�-A<��a����DKD�2{żUݗ���δ��(B�(�;RT,�/��q*!���F��\�T�I=@6( ����h5c�P:����VL�.�����%��Я���'�5ywg3g0�ka�
��[�z�߀Y
����)clS�ȴ`�	6��=�o��'�~�e�LÕ�^���5q�[/5!��T��p��(�\�z�Ob�d2�~���AC���v��4s�q��,�Y�8�_�^v������<��2(@�����P 5���qD�4�;�$!�S��p��_)�i����h�30���fă[ӑ���@��m@�����m��C_�~�3�Hd;��r_�.��A_�>s%)�	߉*��k��qЀ���.Eŕ08�I"���f uYՈ�%�y^:^z�t����A��|�O��pb:3� ���-\L�R��TA�na����~��.�Zy��]��KO?��[zW����E`
�P�9ȭ y�������M.�>v:(UD�v�_���o�ϥ��م0�CT0t%�=t�%}G��j���N1ÁT0ն�M�e��RO�yv\H�{x/���!���.畃<�T=_~��ľVb�Uw�5�\If~��|L��o�i���^��B�K0Ţ͐���;�o�Љ��+�i����o�h��#	f���?aSj���+����&fC1Fž�g-@�RGu��ٌv�6U���^��6,�����䱩��|^U+�R�o6Z#���b���_�����'��ڲ9����u!b�wVP8�p����"�vJT����l`]��
�rU!hMk�Z��4�㶇ۤ�Z��-�=���|���q��B�@�h�?NSd�������51���'n�p
�1ӊ�I:�����Fǀ`gG�� @�"��mf����A�%��9���)��
�L�@bi�E?&`/a��C����Wr��j ���w�D����O�%�$>��49����dPt���.�(?N�i떫�zv�a����{b=�?�b���i@n��v��_�U���L�a~Y�-)(��&:�Q�x�"�D���Q�f��D4�.[[nK�J;V[�|�']/B#�$_�#}H�qr�N�Q������|5! �E+�U��ԇՑ5/p�w	{��d�w�p:�.J&r6�Vl;�/��4B�ojZ�oJ�~D;�� T5�}&O�hQ� �G�C����b��jgu�af��T�Ho����y����ƾ����C�T���w�bK ��P-��>1>H�Le���y߯�R�W��L�%�(��
�1tPX;�Kˮ��=3�4L�êR?��?�s��p� cD�f�eP��$ͿY��cS��$��<�v&٦��wm��A�b ������2tj	$��}SC��oN���_*� yH0Z��:���a�/���2QzX��o��[7:�r�Q.��<��}K��5�T@�Tq��v\+��3���-4����RQyj�$�V��=>���ɶ�3bI����V��c4�4O1�d�ڢq%ÑM|y]j�ɿ\C��jS'�Dɭ\0pR��
K`%'� ݢI�V �����x�"����ϗ|���S�"=�3ʜ�xT����K?���Ѯ� �|�叛�4�$r�� 4k�q;�_����/�_���r������JN)�Af�+-qb��7�.�1��ugt�l�!�BHyU�k��P����^2M��2)�\���F7�<�>啥=�Q6�b�S{��Y��\Q鑨�4'�ciZ��7/���^P�	��$p�#bHNy(���ׁ���U�A���(�p»a�x�K���{D�}4u:�2�Z|M����H�	��-&�L@`[��V�m �a-���W�Ule�9�[%�\�t�;������1+�c�A�r�T�����;p MH���j��v�b��Z��^0�'��\j�4L鵸n�Mh�3\��oK ۠�P��8R��V/��2�(Ћ�0�@�~I�#� pvd]0LF��h1P�� TK�|�ē�k�m
�xo��u>�2y��Ksh���"��,>�Z�@�H!�h3�׬o�+�37��h�y�r�
�Zp]��\�����T��I�aq�K$�.@y�Ʒ�Ź��'���O�C�G*�;ڢy���-�"��]��_"x�m1U7Ei���Q�$��q�����c�j%���,����s6�����%�'F�i�d��f�Q}緲IAjA���X�nP�\|/ޢsc����ae�������°!Tk���x^�4^|�s�p��5r:X0C����y�%�yZ<�Y\��c�l����,W�p�	�L�.k��of�Yf	�cm͒���=��:0����R��X��K;$��SӮ��	Y�.�a|��6M�O������d�{���lP�V|~�:��`)�ӏ��4�p�?��?�>B��A"�$0����b�$6mj���Y@��N*-@'�ӕ���.��4�+ֵ����g����� ���jn�)E�X
��h��%�La���&�y���[m��F
�ߞ�k�i����8�2��ɄS�ƕ���ǥ���x��3�>�+'s.`
^y	��2],��� ��х��I��ɰO��C��̟9^�����������5��x�+z~z�^a��u��Ķ.*����7�
gd�Vm�m
cĴq^˯n���(��<����I(=��P��P�y����휨���NK�w�������}Ì�q�9�w���E�+a� �g`�v�/b�yY袨��1\G����bSj�=q�ӳce Z��[��g���1��,r���Q���5������oQ����ʽ��1Cľ�� ��+�:@[�:b�������,W����=��8e���!@t�<���Hv :R"�&~-(��`'k��6��[  4%�Rg'#����˔
/T�N�_0@�c(���y`:sϬ:f��>�����C�Cu�:�*�t�,U�(��hy`������L$�y����r�!�aF����h���啩U����z�3K�`>Q��w�ɽ�$)qt���v�~��`g���
��R�Ss��.�G���6�S�P¢��J�	�a�@L\$\��U��p�'୔e�N۩i�����2yP\k�!�2��B�H�7���9��Dl��r��(y���*�	%�/�O�!������֮f7a�Jb;��Zr���$.��S��c����[�>~��=�z��f��gcJ��5��֜O�/lЛoqrwvW��~�rk�d �YVQ�-�ٚ�x���bZ$XYL�،E�F�j}g�Z��h܆V��shJ�2.�؆�����ն!e��c���)�t���@V�e�4A��/+�h_;1%x�4�>��� ����:�zԈ���˩�_0��g���~a�Y�j/O}_Xz�����"Ś^�S`�����7=l��k׫�~L����<F~K� <_L�h��+�﮸mFFNy�p�t0v��
���������M���"�'Ӣ�Y��N�6$}Q	�Q';�e�������j��ۄ��N��UoH!ۘB�2\���r�����ևY5��U�K��(�Z	�6���>&T��<�8����3S7�p��e����G$��ǟ>\���M��EI�"�TO���R��P��qw+�]��1���JNΖ�	ӥ.Z�j�2[ ���To 8�l�1�ٳ ��q���G�;j�6^�#��b�g�g9hΌ�x<f����X6`�����.��3��Qϴ8údǽ,q �U{HP[��x��;�qn�c����iF]$v9
?-H��st6��FL��]x��
�� sJ[�8grC>�O��![���ǯ��Y�4P��J��fDC<��H�8l�
�9��S��&ZM��Am�1��_��;�Z�g�����+�*��r�/���fbr��g���#
��s��h���	䥇DM�fLl��Z�)�^��u�&���Y\ӎE ���*L��⩥ǒnB| �t��T�`����x ���[��ʃ.�����#TPڡ�Nj�������5�=���z�C�ɔd�cQ�J���1�+��0cB\ H��M�M�u^H�obo�-�<�c�Ӊ\á,؂q���:xD��ᐙi�$.�w&��m�� ����l�	_Y�i�r��1��O�;���~+K���	t�.�G5����X]D�-Ւ�{3'�H��'�L?A�e��N����&A��0vg�1ʉ.�)�?/��w�_��&��~/��|�����w�
�#���6���ASx�I֙�Ơ�����A�&OÊ��y�3Aֶ R���䣊O�7#�t��}�ίJ��Ň��F^��<�Xt�1���������&���8�l�uSǓ��,9=��5ұFΠWc�[.���?�2�ǭB�� a~�(�.���C�
|����B����'�xDp9��1���\�7A�ɥ�Oe*�!��)@��q27�b��n%��w7������ics�����S�Sؔ�<*4��p0e�2�ul�\JbK#�͹�>�\z�ft�#��l��bL������2M�ɡ���W\�jo���,�Z��9��=�v���2/B� 49tE]b�/�t;�bG�Q�jB/�е��Z�� 89�e�:�:U�A�O#j:�_S*�7�� E�'���i�����- �ĉ�/��<qGt�5�C.�~w���s$�G����W�a����U7P�A.r���+���)9��K�&��u���D�	G�k�X-�Rծ�)���"���ڜI4mm���<<�~��(�i$z��r)�<ٰ��BC�P|�Yf��%�J���p�e��+qO�C�s�,}X�k���� m��S�@	�F�l����
��P�����L��&�D#8~��ݑ��o�?�-�8x�.Z?���g�08����5!]�����Y�(v�Nü������� A�R���Vcb�=tL贒�����8��8���2��S�6�9����ӗ����+�H��{�b'�
?6+��<����~��;�)[��k�%-;b��$V�	��ຽ>�mO%:5���-F@��p�1�p���y�!ʁ���3��I:���IC?.!�:G���)T��H1���QGc�Q�:C��<��vm�]o�Om�M�"�.�ʑHݍN�%��/�����â�[��z6â]Nd��r��N�;��n��( ���N
1���	|�t�=-��2����N��%<B#K�c�����4���5������zCrZ�������Г*����o�����Q]����J��ƚz8�2��@�BF�Wc�W����P�h�3�=�M�He����)%��.I֖vO�ߑ��)����@�G�M��6��ֻt�L�:mKE���p1(��CX�_��t���:�y�lڊ��Px�o:B��n����Hp����%��F%���tB{��Y�^o�o�uO�m��8d[�>���}Ƒ���F��I�n�8D�L�gS}X51�eO�����;H�3�P�BE� -�9JX �tq�[�_�q��B�O�T�q>Wty��ao������4L[{�(q��w��n_w�y�nEn�����KQt����6�̅l_�N-����0�xC�/We���xe���0Psc9�<�Þ �2�f�|�v��t�����;F�D&�f�Sk��Ӹ�_�bY����0��TL�a5���u8o��] �goi%#H<ӭѪ#��̷z�B�n�W�m����j����Z�����_���7T��{z"�a�I�(�>�w�AfkBN��{x%<G�f+p�9Y��b(y�oS���*�z٤�bm�Uь�De"$�;|������4���*�8#������	پdR-ox2iL}�D|�ޡ�e����ET�i�y"p)�����VoKcᲦN����/�� ��Z�e�n�7*�������dE1�����(T�=�HBT���Z� �}�-����/S�)����2�|�E,0��:᪅Ni��$M�l� ��VV�7�+�U��h�3.�{:LBE���wV���p��o�t@��/s���/א~�]޲���/�,#/��e��*]�-�ekZN%_�>�&��0�(�ɋ�@����}�?�K^E#e���j<�䪤I�������Qp��� �}����\d���H��Ƶ^��T�G)��{��%��
R�V k�Feܞu��zVX%��Z�nKZk��}��������+Q��ێ����f%*�
���nQ����)�n��Y�l{����vZtۡHw���(18�'��lA��s8�^��#�7��_�&2�_T�JQ�*�x&$�*a��xEb���4��'����n�4>��W�=ל��}�67����������%��d@��L>C٘(�[���Vf� �ޫE��O��7��2�hq�!8��,] ���P2�������|+p��z<zｉ�0�_�r�1�^?�blJ��>��dȎ�i����,<&�F�	G��}��:9Ț�t��o�t|a�C,�m��\�7�U�1� �;q�-X9���^�[94��Ga%���i7�n˰�`�S�^�dh��L/�CMCs�8��:�wք�g*��v�B�&x��Ӥ�����t?N��w��w1�}Y���R�dy�e�����˘�+=���:FN�Yv���:��˖ӑ����j��e�b{ <�O�v�q.?ݠ�]��u`Y��[L��P�a��{{����+"i� ��#�h� @�q������E�V�Q:7^��_���s-�e�U��i(�N��B���Y&�d��o��0SE�+�a�7Q4x�����⋲dv�֊T�_avǆ���YS�����̖dƅʯ�ߜ��?h�����:��E;��-?����ҵO�H[IDɬL�M�ߦ�khYͭ�"��c��,�&����ٶ�r���N(�%0���vR��?�m%���B�=�}�ȼ�aB.e�ο[M��Pw ����^�-�Z
<�8D/���JO�ǜ齫[B�rS}�7�*�_��2� :���;_phˡ��.�l;��|
�D��E��P����2��� ;�7}�(��P��u�8�RH�@�q(ۨ	��D���'���\�x
*㔊����~�. bTA.�`������8�إ}��r��舥�1��,j�A'�S-�t���H���omﲮ����١�`�Jt9�z��)��9}I�J��uI,0��F�$":]����Eb��'�'@JB�oҴ���{Ja��짥�x��%d�hn�$�QF,�ʌ��]�D$��;fK���&�-ni2!#��sB+�ʠ9�o�)�Q�r(!�ۣ����0&��dfW	�<m��}�����w����]��̊0�Y�ޭy��R�R�
����8� ����q7��=\8�f�t��\QO/�p�1�mo�i,]�^���gۋƐp{,��x@���*$^�A�D���+�R8n<�*1��b#�k�̔���fl�r�"m�X@��D8�N� r礳1�o@*�j���%	]o�#+���,Qk�4n��.��K^�3f�:l��;0j
]��]%��cnyQ��G9@4���AT�S��kC0q��Nᩱ.������#1?빵�MU���t�#��O
�*w\I�W�>4�tA���~�֬��/A��s���n��/M89GT�b��Հ%��PF�D��n�1m�KV�jɓ�&�Z�*� �:����*��������B:�}��f���n,�V�R����R�j�`�Z��<��C��~�O�����]ΛXUO�}�����`V�^,�
���a��D�� �$��ҕq?���O��v�-��J�\�Κ��j�i�}�_Hf�˳$*`>$�Kqc�yCc��\Y*Q�0:�1G����q��|��9�>���x�(m����&p���I'7���Ф��y=��Ǵf0�������UB,ѩ���á"�]�q��	D�[L淂����.��2r8�Cu���"O+d��Ö���!k�3`?������Jm��7io:�t,�h���ʁ��^��6Ȅ�l�(XAr�=ʡ8�K<q*����	����>TeH�>B[��;���j�@٬ rT�Bn<�Vv��_<uH��M8���L�|#�m9�m��#%
�{��'����YEP���$G�6�_X��������/Wޤ�]C�`#��^i;L[QQ�Ȕ'�F[���7�i�+���Q@m{��%�M����h5WƗ��8
&��,��A`c����*e����FڨZi�5%|[�)1g��k��8Y�$,���-]�K�=�y.*S��@��/��e�OH��*�)D�A9�&�fZ�^35B����ٵH��@.k$���a��F�]H.9��l9���_߶gpc8�#r#�6;J�P�� /��sB����n��_krG΃�-���kiB`Y\r(��[�������M�=j����V��0��� 3V̈z���o
R��4����a�!M�8�1��25�y���j:`olDT��&�����g*_wQ���-��wn�u&39'���#��5H�3�Vk�%�0��b|9�P�_3g�1��~U��O��ۦ�k�tg�$�~ ��C����{.(%�˙�O:�<o�{_"����1���ρn|U�I��J�ō��K�8�m�¢�>��*j���vK�U&�Պt�z����M�d!��J����� ���6AJ�I�[�J]�#�]�V������`�3��ΠUGW��O���3�86�¨?����hd9��߽7WQg\�Xz��K �8� �QN�c�.&���(�b�_�\M"��6L�����Ҏ�˧�E�m��2~zzu�kc�p��p\�u��Ec��9�{)�q:�o���?[f��_��n��
�P�VF	~0�jr|ނ|Y�3iQ�<����:�k���ߡl�:.{�%{�'q��z`�7 �uf�������hN�=QM�sT�;=�M�yUXu��.6�ԩJ���������f��3|j�+}�3ކG�"rV�|� -�^�;dd���&ћ�B����Uyb/i�a�ðR�w��9:SOc�?�~\<}�U���(��e�+˪��>�n�x�������3�ei�{b�k���6�=�2��f���:{��z�I�§l;.mW:�_$zFFUe 5���A��-�1�\/w��	_�jX�g��}ɜ���^��{}�3�=Uw�u���x��H�!�ezrA�Y��`��5��"9��"ވf�qU�gu�fW��� ۉ�j#�}�L���wWfJ
D3��ڮ9D��#�M�f�%ȵ+F��ȯ�;��{`�W�ME-�U,1u��"^v߶o3�M=ԴN�<�����Wc>��pd{�7�6ws��uJ�-=�B�����;?h�"O�)f��$���}�����Z`�m�B��jW9$�PS܉�
Djf��n�˚�1�aҮ��w���4��R�����BǼ矻��%c�op�7�%�ו���K���:|��I�B(д�{�"^�hh3��23�)�71��y�osGt"�%4S��� _ad61V�J�!Ԅ$�-�\Zj�E&M�랑�f��l�ƴ0��"�-]=]�x�Tߗ���DtAZ�wQ�|�B�r���'�j�:��o_�����^�˛�ӌ�K�W��
϶��e ��wT�:S�ܽW[MV@�]��U�D2x��`�d��c���+�e{r���Qlf($�4|ꚾo��5d�>q��?tF�+b��W\��O�*i�yB*�g.1{?B�,d%^��*N�K37�r�rj��H�_�U|��<D�<M$A\�+���B+Y�q���	��L�Y��:�(��'�����^���9��fcEBom�H�5��)�Pz��4M����/�VM;r��0$�w��K
F����ż�	0���+�e��~�`�v	6��+�.�����q-r��R��^] ��	0~�L��(�z�����e�[� |�e����y�)X.Yܩ�F`jl���ct��R��z�ɘ�uxF���pcW�W�TZ-7������&m��(�v6����
��w�ޜ����8�ŚO&苺l�r���8$���#��B=݀�����$����j��j���	,/�-��d���`�U�[gz/�l��v��]xFw�,�y�(���Gx?��g�	�R�z��Z�1m���E��K	c���*��#�卨� �BG~�t��+��������:9ȗ
!�n�dP�v�]c���4@�1��)s ���ű�a�`Pn�]N�(�t��jD��0�w1ASr�4��e����c5���������^.鶆��n���?(�7���䶑���Y�3kB��?��e��ޏ�S"OJmt����I�+�GCv���)�j�����3TP�'1�5��g},��ƟrT��`���a�Q�K ��Ԯ����1�ܭ�3�b��V��{�5�YڂN�e>]�<�l&Q�8���������^�&ty���bS9D��k�P�.T1
8WyIݍo|�m�i�@7�.M���od����P��.�$S�����N�I=�����F�F��J�[��N ��qm�F��T�p#�>3��"(9�n|#ښ�:��G��:<&�����Ţpn ǣ#������R�YQ�Z<%��)kH`��
�xk�-�1�)?��v�������<"���(_�P�T(������\�a����!��ft0d0�n�ʐ�T�r����E�E�<�=��r�8),��0�/a`il8��J2��˓C���6>�(���uZA�"��g�we}�W��5+eD�᪳�v��Ѓ�-q���q6C,I஬�ѐ � �7�Ӡ��+κ�3F{R�IG8�?F��t�C�+��IK���SȈ�)p�)����6l��!��?�j����������l3cU��[R �c3�3��1O��.rb�z96p���J\��6���g�HT��`�[Ka���n�3T�}�_<��pA�YSMA��CIn�
<�!G������Ify�1U`,�Ff���˪�q� �^�3
x4�@�^6��l�h𼼧*6���p��=lU����C�|�KSwKkx�B��E/�@����jǨ&�6H8+��dMz�Q�C���>>�@��i�5��а�,:_�T��ƼO��@쎌�G%�����N�:`��sm֧��
G��9�O����z��4M\��Y��~�_�Ak�M߾HAͺ��?�Ȧ��}���U�>��/?�dH�ke�U/��Kɵ�ձ�C��cn��uQ�K��חX%���D�?���r��޹���SG��(jo��WX�Sn|�;=���9������}���G��R���b�Q�on0e�^�;I���e˔�ks���k���o��<�y��\r���׶R�����,o��G��; J 
F��x��G>��/G���j/�Bt��k�b�´��<$=��r��P��b	y��~�z?���ŻV�t .xuV3L8��Lgf����	��<��H�4�%��OUb��^�J3��r`�K����=KP����t���%��@��(����K�@6O/=�Zz{����gMW��s$�LQ�r ����~�p�3ܫ*8��n$b#����Mw#���]����(c�vq����@� +��G���c�_i:���聞y'��G��4�ő.�(�nU���	�v�eל�h{�X^7ꗕN����T�q��)N_�.�C{.r���0��Dof���9����۰|�-�����%S��w,S�A�����aG��*t��`ŀ��O��&�[s�y��6<[^�D.{��,��ڌ8�+���~>���S�DP9�ӎw6S�U�6S��6�� ��,S��P��X�ٵ��w>�I�tZ�=������� ?c�'@�a��,:�\�_��֖�>��;�=G�Kv����4fV�j�ݬ���7�K*u���J���o�� y���Q*a���
/�����1U�A��wB�<����'^��@J�uD4�צ��]��`[,d������O��8��V�rM�;�9�9�G�z�H��y�h�=�����|j�f9@�`���Q�G�(^#q��7�RcmKí>eqE�Q�ԥ)�s'�/�%����~y��-5M&&[�)-���(e�tit�� �e.T�uD�5K�1��8ʙ�cC�1���<xa+&x�i�=m+�>�`�}ks��Y�27��l<�]6"��#j��M�![�$β�-��}[�~����W8�֙��\<����xi�_7��s�@K���I�N8�����n.�(��z]���� KX����J���\��/a{��?��/\�ؗ�� ���}j�w4�>ΩK�t�].D�&-y�ƃ���ܽ(�	�.���M�W~̻w(�n\R7�O%��ӯ��^�K���Lϫ�6Ź�!�3�DE
��M�#�R, ~����/*����W5�o|N�x�G͕�j���g}H��ĳ
�]x�l��[U	L�^�Z�ڳ��	�P������F>���4��ȋb���G�T�hoSVk
:�G���P��yC���|5���q�Z�ٍ�[v����u�3O�_�yU(��N�_w�L(Z�W��Axd�D���c��)��'1����9�5l�hQj��ک4�4��x�h����m�q�
]�|�F fS�K�)��̚����PzҶ�\��2�zv��Y�7�����'J��UT�չ�`f����o��8[
�P�]]"�ID]���UE�h�`s�&a��·ގ� խ�H����CA����(�/gE�ql�7�鎱_�TS� +�B������t��"̼�:�:0�uYA>0�H����h`����@s�KY.�b�s�ǣ�4��ލ�K�LC��jڔT�gK���u%j�&t�6�߅�$>�z߿I��$��Llna��v�jih�i�2�I����8��[;���`��f��X��m�wr��Z�����_�\��<!�!ḛ����vR��~��j� �s�(�{w,P�_�#�3��B
�K�Nޤ	��{��΋k�w~v��������x��ب�
)�	��붦��3��8cdC�}��p��T�7J���] �7�Ak�fAV�Z������mS����"1�^y�i���N�#&����Lւ����� ���?����H8p�c�!����.Z;��PRfܴg9�2�k����y���yL?ǂ5�[GB���<��[%�o����mRHTQz%��Vncr�H$g�p�G� _���6�L4��ьI:���S����S1��֪J�FҔ���^��"P��劄��x�N��^�7��K�q���&��G:i�!�7z��� V�ޛ���5��ܺ���Os�u�߹ޕ�_��0O�~(�Իi�?�A��D4c�/���nӿ�0�`TXD(!P1>{ȉQ�H˲�tW^�X��L���x��\pk�1$�O�ތ��F���;�Q"�IX��kk9��A封>zW@g�*H���y�_�׭פ���Bg�J��w{v�-��_��
�]�5�6�Ȳ��O���Q��ͨI,#��HVZ��Wdm�T��͖��6�Ǝ����F@妪r�$V�5��ǽ���������g&��?�1.�.�%�q8T�zU63�6�?].^�)�ᔤ.�F[��u�h� <F�Q��`4b�tx����F�g�Ė8�v��=.��5��#g���J��P�����c)l̬yvʴ�7��3�&$G3<S5��4~ ��)�&y1�E��=O��7O�p}N<���=zo�d�9����&j��V K$N�la,�ǁ�5��!0j�"8��߃~��Ȫw�0����ŗn��!CZ�_�c	�Ř��Ǒ}�V��L���J	-���?q� �p{6 3��-1�1'/�M�K폔A{N�
���-�3��<Л�K#��9�h �~>�R�q��\E�+��_�QIx�܂@����� ֿ��!�ni�7���'��"����~�JrD���A�X�T�׍���G�Fғ�7G�����BC}�������U�a�J�x�H������w�ǐ����a4�K�B�D����9������R��;��T�@��,��}�Rse_������ �1H�/{��;K��|{oQJ���Pv�뷰+�0\�ẫ1|��hްT"�!�6���C�t���"���'U�H�@�/b�(1��Y�r�o��H��Z���ƪ�C��^�@)նqA�<�i��/�4�����k�#ix����,k�Ԁ��B�Oku�>	�{Xk���f�ݤ��F��Y���V��vk��ZS
h� 9Z_K�ߎ�-T�����+��V��><��W�]��D��
`�-�2b\t&�d�`�m�ڭ�<Ӟ�5؅��[�f�gT[}
	W����<%�?���7�?����$|{��!�~5@%�)�"��QH��$��m$�T%M���H�����U�'�(D��Ko���uO�{@�H�=�ߞ�,¼����JGI��c��Z �G7mS�LrI��9��W�tv܂�]���TM��[
����zC�
o���ߍ��@�-�P��S�;C�1�g4��G Xs��:6��o�L��$ ^��Q�x_!�_�aN�U����>�hKJUz������$+��M�p�����g{'�I���R�/�W��<�l����U�:�6�蔞����p@���e��r(���1��@�M��^9w�(>#gb6��k��!���z�0����b�Lb���N�ѕ	��w�_�y,<�NDOm�|Y�C����k�f�jg.�	i�S�3�w����F��|
ޑ\C�y ����R�w�4W\���&L�E�?�t&���2����vv�a",�؟	��!�51(�J��Ѻ��3��l���<�K����~�O��7+Z��g��}��͵u0�ن���U2�pLs\�c�Z84�ikj-*��F6U�h�fט�ĥ�ذ��4���/�0�El(6�����S�8D��M'�z��?�F=D)���1�
%zAgS�E�����c��XRi�F�Y��ȁ�ǖe��Lq����=߽%7�:�V��^��Sz��Ħ�����T$QD��&spC�|���y~�}t	I:8����U���+n��*��ԉ��\%FJU�h>��z���h[�@�_i��/aDj��>�g�8��:�@�{*(	�Yʍ����w���s��G���<�PB��cp.p�/�F0��xƕ��G|�
'�ʙ��,X�2��8�wx���Ҳ����;p�d�{m��6��"_�JU�R�& {����'Ĕw>��>�l�!�*^ v7}�ǆ=�fx�A���ͦ bv�ޅY}9��8Y	.�<���W�Ǟ��h� s�.��a�������6�w��7t5�Zb�G1b��En:�3'�s�N��+��.����Y�~SVYB��㏯��U\	��l�S ����v�I}2罧���'H������b��p�m���ۚ��乆f�#���Ɏ�"��M(���X-^I���:�%���9��p�~/D�p�Ђ��ׅ/���u���gcs�ܓ��|F�$��1�׌��v�<iUh@����Lki�������4���'�5��fY��:.iJ���)��:�� w\�܋�����W�a���*W�u�������N8OԔ�'�v�v���:FG��sY�G����\)��1��Z-@E��􎄼���3�75�G3�����T8з7}o4%��,P�� 9
|�)[}��C݌��x�G	�-j�|��ծ�K�@[>j����=a^:�TPu[��>ï�=\gi C�Z3�}?�a���8�\=�@ClW#�z�x��
?�ܶ輺ɥ����nr���j<��watu��`p���
�bl�rކK0��b��(�	_����w)�)�I����N�SFmc���
;��mU��]{��x_�wx3�>�L��'��	l�ۅ��T�
��&|��B@�:�/�h�mR@�"��Z�b�Дa�瘕"v�_k�_J\B����{�!���	ߴ��Y����8�k��`%�R� ^F��J�3:�0y̧@������ۄK��,(�9���iEb�f�]��mL�؂Z(������!��2y2P�Y�۳"kx��f�i�Cx�#2c�v��кc���,Ʉc-�/�W�ǹ��Z��	��� �]%�ߢ#�0�AB�5��c�!�����Nٰ��j�c��(9Wa"����#3^�ܧr�2��h���;٨P�|k�8I�вٙ�?ٱ	��
��<�tQꖹ,>�cg� ��|aV0A�<FdV�w)e�mRϼ��Y}!X;���$D�ˍq�83#�?N��6q('�Kl3�ͬk�?R���~�^�[y���Y,)#u�Г���&���9%�}E�_M�QO�ǩ���{eх�F�1�G��78�3|@�=흻�gP|��I^� Y�c�<�&V�Հ�cw~b�\������ɬH��e�A�@A��Vr�_h�/�+�>�g]�7;i ��kd��|k��'��E���ɽ�+j�[3 ��M�u
+Y'�R>Q!d��l��h��6Y��|1���O����]%{���[>r){�.��x�?u�3�����犟%^���n�>`�Uu:�|"�D'��Z���{�������o�Gj��F�Q;�;b#k,nz����F��A�s�X�ҷ�:_�'�{��`�ݬ�Y#ݿ'��)Z���������N��!2�!�����������6_��ڹ��T���	k·_V����U�)����V�ރE������e�:W���fTr��ɫf�C �s���R����Z�zz�t~U˔zG
)�Np����y6'�|)�EO��w��H#������_7����+l3Ϻ��ZG��x��5����.�,|XU�!��9<�%[Á��>%Y��Ε�"�T<
4��-����*�/�M}���f�DHUE
��U���$I/n��d�/�@���v�G�zl
M�:��s�l���T����+��S�da�ci;F�ߞ\
�T���<��GSսZp��;fę��(4Z'�H|��s)�=k��,�	P�e���R	���9U��L���_��ZB���S�T=G+�M\	$j;䤌����{x[��-W/�K�e��\�FfqggH��C����\.9����s�
�#�"��Gh��-v���^	����M�����[*���0T���iR�L{Џ�뾜M$����v��ٞ�-�}��-$�*a����]e��t�|�ә�E>6��)�|T��ݽ`��9�����B�>���a�����@;e\�D�[�I\k�ˤe%��d!�GBru��O�뇛# =;k��c�v,8����Dr�?����x��	c#>�dl!#�rnz�s��Ꮏ�A�_@-�<��DgQ��dsZ�}�$䍂�mE�8��(��v|���(.3W��c)(���˓�!(�y�v���7{���P�����G�/I�.�I���e��@�E� ��_ %��q�Yc���ӿ��-���j����>�$��Zt���)ϤmP�mw $��=l$h2����
�.�R�)��l��@�P]~:��&�o&��;���X�8�Q1��d�~y�_ˮ�# 7��~"6�jS��D Y_c,=���^����2�&���M>� ���9_�A���s�Ĝҿ+�&x�Ƿ[�<`E�_GDJ��[�A*���M-js����a�U��/}��*�Y�Oqnp����L�r�1J����T��]�ڢs|�%ܬφUW����z��o ��n_jl�L�����R�ѽ�u�!���h�5���Sq� o�3�ZL}�|��;(1���}(a�Pn΁e#Ѻ���~�4���k�1u*Xj�
!�pv�S��a�f� ��9E��f�Y�K�T�7�`P��H�/Z�lx�\9�_�φ�i��Z�R#��B��;y �~�q�{�rJ��[GBJE��w1���F��{�g1!5f}��qLX���12�fO�{�w[�+1�����0�]�s�z�x��S��S�c���pJЌf����$�8� 3!�o1�d��c�4�Q?�{�1Ex`
�/)�MK��Vq1��VD�ĝk��4��h��H��BzA��q��r�Z�Ǝ)f.&V�>f�U%.�%nZYZV�����Zzz�'�J`��#Hv�@/YT�j[�`H}*���Ǡ+��+��
��W<�Ky����hd�d�K�$��������|�z��C�<i���<Ur�\%i#��ڹ�+�D;ga��P>e������b������O�3�j.䂞�;�E��5	�!��l�d��~�*�leV��s�0��o��f9���m帲[=/*A�ZI6�3����
5W�8	�p��4��4���Fm�8�>fVB��o�cg�alK�`�V��!�5-�ʗ;3�6�I'G�y�q���桾*;D�
L\��P��C]3By'1B�� �91���\�������i.�.&+�iB������ّ���'<��!.����xuA���L�3a�%TM���썍b�c�����ȫw�*�[^�7qw��-M]����`�XT*ɴ�
��v.is�O�$M	,vqg)�ٴ�a���Eu��cr$ߕ��(٪W��ǔ܎�FB:p׉Ӈ��/�M���x�$�g��{6�U�RF�D���C���}NNf�j��	�|x�u	+�{��୵8ڄ�|%�݄#Ǥ��=��0^��
�̕��2��z�M8�\�tm�Vh���N;�@6��mh)���t��֭��uvC��v̌��7\tg�ѥr��� ,�4)���t���|r�N���hy��Xt�z�4B8�;ʵb���t��6\�'�Med������庣�-s��#r�bz��A������:ܙh.��qI��_����8�09�'�1���:��F?���]��Rr�1��1:T��	�I߷��Y�l�B*X_���a�T+b]ڨ~�VE�M�t\��B�^2��O��Qw��prT9�;Z��A�2+eح^�wh^���=����w�á��@�t$-
Z�sz�Ke��&��"]!�J#$`<�����I���5��(Ģ}�b�=��]u���P6)iЎ��4e�
㉓P��@�)L8��H��YW>��;�r�tjo>�p��K2ER�i��@3��_�yv[5����R��Q�;=��(1{ߎI�L���u����wyP��D�����Z�e�:<�>�"����@?�a?<n��:zȌ�`���2�K~�����nb)y����S�/��<�fpՒ��g����K�R����'���_�W��?�#K]���|�a�Ͳ65VM�S�9�Q�{"�P�3ʵ�5�7N��"K�Y��L�B�v TV� h�B���5�R�a.{��l;��.�F]��f��K�_�5���t�^�g�]�^��w,��y��&��U�?)/! 2��*M����7��*nڍ_�j;(�[�����$d@��`R�V�S=�n���[��z�o���A/}���Z1�*!�wU��~��^mf><��T�������Q�3x�\S�2*bФ�7�^�W;ޒ���`��=3�o������_�6\�E���Y�ؠY�K���H�{:�ڎ��f��)�8"t��@f�������?��am �z$SJ�9�S&~�/����]�t-�G9п_�pF�!w�b�sU�g�퀏��i��-	����_}�ޮ%`��?`�NKx�Ͻ.O\F��z�gQe�e��f��O���-��}&;�����S��p�$||Q;Ia_�5�� ط��9j�18/r�#D��fp�R^?(*��m�J��#F7�����Yq_��4��k�%c��R�ӉQb�U�3[/
'�xd�.٥u���1\:�����$p���qQ�Τ��\t���X j.��뤗��?W��� �d�\84�c1ikz�	�����U�j�5r�o&�%Q�����j���J�<�DFcCS6gj�ܖ���^�5�3-����N�ctj�
���7/�
�oUO2J���ax�Xaш����]C�m%lJ�2ݼۨu.�.;�=G���&��ًS٧�7����,�V�>ݕr)I>�Q���ӡU�@�HZU�����c����e�4��ʯ�㗛�7r���e-��;����"H�{c�^z88*�'7N� �yʁV�����wa;�ɲZ������ױ}��sX3���sǴ�)Ч��Ϙ��Tk�!�:B��S���+D�Z}�5tg��`g�W�Cߤ�[E��,V�o�\�:��%^�����CY��=��+���Hߗ��q�s�Y�'A��A��e~��et�.�[[�:���N�>��O��M_����pbvK��}�d�Cc�"�B���wv���l��z��1:����"�1	��>"�J�Iס3iu��(3��X�Tx��"9֢a�/�=�h6�d{Ogn�~�����	�i��> ��y˜�e^Bj�y�/�Il͞�V?�}�{��|߷�w�D�9����q�9|uj&_g@�b�1~�0ٙ�g�wiS	�]���5�KB�K��kDf�!�ڍ�!i��_c��!�����l���ļ<���e`� Q5R�{@uTP��Y폭K��F�����LJj[K+Cg��L;ߕ�-���J������w���D�W��$�0	�G\ޒ�,`9%�(���a^�7ٞu]� ��� ��n0��t�<Q[��򤹖���`�F�1���[^Q��:+�<?��}4��<������� �x}��>��`�|.�U�玌}<O���%MY�wY�v����l�p�H��?n	i��ŪR)�>��Su�E�c���(/DVq�Hc����l
�����z���8U@t��(��?��3`�πWi����}�B�oŊ96�/Ò��:�Z̃���b�wޡ�QC�|��ue0�4ň~:9`����^!t)���*M�1������8��4shה�^��:m���v�q�����ī�������|/�%IX;U(�>�];Ǻ��h1�T�W��>+�(M�EA�8��04j�rR�%�^&sY�[�An):��������Q�ab�FN`*1��^w�I�Y`���X���&�-dĪ�e���iE�7�K��,f��<���4�
)�o��}Sr�u��@Q��8B�vZ�xa��<�Cw�%�0��Og۷H������P^�k �<�aN�f�x�T��H�[�%kS1S!	s[�.���T��R�����u�~�\�	���y���nR���i,��Uz��AB�C:8�Y��GLC���~̢�z��3�)9�Bk��J���8�v�2:�e�E)��t�����Z�\Ʃˤ)F޼��4�]��!��+n��҄�E��"@�Om��kT
]������Q�mA�u�Ho�@��Y���Q������<��&��9���6=��B?�w�_X&j���[2ρ�I`����Oz���>-I��¢��Y�rrd��-jL�զZ�#����ʰ�{+�R����v�1L���ջ@��*�g�\#��5�=&ÙB���s�0�V����������w��Щ�eo����\�0MD���j�OH�F���U��c�R�?Jyq��c戒���l�o�s愈m:j;�LI�4��Wޠ�dYJ�С"� ӮS����Q�K�q� I����2��� �e:	�>����f1�^�����I�Yr��(1uR����=oWN�Zl�wo����u��]Z��*�"x��vn���g�?a�W��u����K��f;�[
H���XO��>&��y�x,yp�s��U�A�7� �']Nvd�-���	 R�IԈ�db�����Di���l��8��C9�#G4v�������[�ts>
�"�y_�����b�
���N߂u�r���י��	AZƻa@�ei���ƨ�(�+[�V���9�(e��}�����GjƳ����c���Cu<����ȕ*���G����FF?H1�ٖw��Caf�ϭ�(u�������i������h��5�S%b "w�����cDLC>J}��o	z��h�H���>�G�ꡄZ`ߖ��M�t;(��ݟ��WY��E�X>r��Y������B�:cw�E~]_���X�9Q�JJ_(�D�j��V��WZ� )�T'q^Y��=Gۦc�{OU��ڲ:����^���eb���t�~<�{T���G�4
Ϸ�$�w�z�a�"]FON]�N�0�XX�w-������7��#M}�|���qy��}Қ7�+ö��6�R��5�)�����GP���
J<⢑�����;���2Hj��g�0������L�zppn��1A:�<g��\�yqv7�x(���>:��KjU˥�*:F��7�뼼��7�����@T�����(��;{�#tt;~�>���u8�w֢^�}� �2"X�6a�"z�����U$���]�_�����`7fɅX��3ۈ����[J�2�zB����ź���H�%3V��y+���2/���B�b=	(��_�L.�]UM畎�>-
adO�p��f\�p�?Pl���v���^�/�S��\:��Z��m�w&[r�nj���*]��D���ئ��=�ԢDR���=mҰSg����M�3ׄ��rgv�Z�z�ֲ3_���\�2��zѹ�E���$m}�3��?~��<��L��_S���5����x�����:�!���=jKч��*3�hQ�Gm����W��,ȁ,�W�*z�s�*�Y��%k������d�S!`0LW��5˄n�
X;q����t;/�.*[2(���2��u5fB=z/�S��;����N�`��O ����p�-��t��d7[��l��Y��,S�S�r6&4�o)s6�I�^�� F=�:�4A+�;���qJ�S����Ŏ��j��&��֜�~�kX��݋Q�� c�.o�t���s��N�09!7���_��%P����� "�������2����CA������ġ
��������ej�T3���� �C*W��T�C��zݍSԑŧE��6V�:i���97��c���S%Q*1A��hE_����X��� ��{��˼g��e�7�,���?gpÛMU˲ڶ:46����,��'���hYB�e�A���y�w�ݡy�ғ�۠i*��-=h�'����2���W@}_pL�d$�i�p��O�ȳV� CO�qgPڿ5�ZO��p�� ��D��$B(��vl%�uV
N�nQy׸�>��Ў��w�JEP!R�TC�����$><j�>�
�?{�pg����	E�
�����e���Q��� ����mOpst6�OPLr�p{�Z���/�q�V����Ô4]�Ĵ}U�!wZ� �(�R^�q����(˳���Qxz=r ���K�J��ox���m��`D���D�B�qQ:��=B�B#�;d'����y~1N砙��/q��l]��m5���0��nx�c�ܜj¤����ƴԺ�.�4��:�7X2=Î��{�,�"M�S���'��I�+yU(%�W7���)��1~y�����,�J��oc!�d���ԉz�ž�@�|���S��If���{�Î@p��ǰ{���0�]�;t�r+�9*���蕣v�j�)���u��.kU����Qdd���YB�Dd�����W�%�d�� �?ܮ�\������a����"����� �@2�P��)��6��4���>A:5srX��?1��d�۾y��`���ƒ�/E���t�N��c���2I*p,C�q=��N|��:j�{p�eV����`�j,x�,З^���+����
�����.O�׹ml��?#~K��5!I�U.2�U����f3�%�4����Y]����#I0���Pn��O���h�~�D��fǙ���s���G����=3g+��5�TX��r��^Z�(�3���+�,�3xa�2����Pn{L�vse�����e}�ɛ��g��w/
#�8�6�����n+��/�8X�����s�����P-�kȱ��>IL��n\�
5aD��'�c7��	�B��t��c0���(���Q� �����eR�1je"p�1_����`���|��n�!%<�CGT����o���2�gE	o�e+��t��漢'�<�Jl��t %;]E�܅@D�O��\�)=����=G\I.)0���0
mi��Tܸa�¦��F;���3�(����QT�8�^�?'�ͧE��t����&���l^��H��x�	W�^�'ư�o=�XL����4��h� )Vb�Y��g�uÓ<�!E�H{� k�g'��K�=�_��!��ǲ��Օ,��?�x���uA��J��`떲����U���Z�1�(M��M��q�$:�5G��L�F���Ⱥ2`<�ΚY�<��HxG�C4q�<�J�ӱ��m���C*}��08��GUc$�f�Gי�V��^�}�: �jS�7�5K,��BD��MTưnL����6����z�n>-?��|�~�z������W�ԧ�X?�y�/4i�x�KA��/����c�<�O�:/UBT��(�NҐA�-i�u_�� �u�:g��%�����lVFQ��fw�^)�� �UL]Ӥ��`�k���Xr��Oz�󉲏E����R��q��kV���p)r�Y���6JP��J�_��ҏ%/�Ir]�G6v�G�7HU%���uQ;L�3aȯ�'�2�;�֛�6aMI��=}d��x�Zz���n$�g���R��Ŗ�������̗���6_�l⥋�د�7�å��������D9�*�z� ��!V ����֠#.�/�'��p��cӈi�\�Q{X��?f�"���<r��"��Z��I27���y�Lp��U�.T��V���)O�)��wz�ꖥQ.�u�an��* m�L��JTėP�%�N��L���&�� ;�����=#9Q�b�dY��5聳0����b��b+PW�W-��b�[}���gԗt^'B�`�g�nT�3-`5�P;���:f���&���FLiXɼ8VW������ٷqz�Od>J:��G�c���0��\~"��Y�C�rCH��'0&�7��������Z��e 
��x��<+[��|^�-�p�������ȶt�!��]��}|��A*L�bK��aϕ&3����w�.WY��|�I�H\�$�^���&�����1�,�2�dh�>����y'��͘�n���t�0`\�p�Ġ	�
($�w�Y����a�g��;� )6]�1r@��
k7L�J�_b�	���}�D�>�a�j֌i'�b��0��:ĵ7����Q �DC8�\� ��vShq���*,鐋l��W�� �xξs��T�X9����gr��5)M�"[�IQ������L+��)�g9-���J�bw�t`����_Ҏ��B?�Ԏ��^��pU`�PƘ��q��_mA��*N}��`��T	[�\�֟ʴ>�k�W��E���婌�#8B��-�nV��\S@���S�G��>΀��Wq?�.d$� 猦܃��p��dLT
����9�e5ͨ&�(4:o�0�9e�V4��k��:�B}�S�nn��/����r{�b��TO�0��W�E�{�M0k���Zq�$`�Oآ�9w�NM�o8�ʢ+v'���u@��G��<�yp]ʮ�I�R��ݳg�[x!�l#�3X�j@Zct�,*uP{���d���� o׮��!%���U��Ej�}��^ D���\�g����OCh��"(yy;�q	�����8v��.���X�G�ĸ���p�����d�#��d�'��'��p���*M4�5�Fx�$�!����	[)����O�]�6��Ң~$��S��6	�ě�$�6[��|�/��6������;��d���٨�ӓ�ieY�[.12�F��Ҙ���7	�s%�F%�1ǀ)<�qm�!M��#�n��Ǿa�v�����h$��J�ٳ���*�}F�
���
��y��_<{�R���L�?Y0�\a��B���%_w(#'�~�8��Z;�j���<���(	�D8��F�
��9�̛o��}�Ùf)R'pq��\e&�]��?ɵ�1���|���ֶ��y -��*8�l(׀{:^������P�P����w��AXL��J�� ���ܻM�E��O�Ugi�:_}�9e�O,I��֗���.q�:Xy����=퐯"ޱ��ք߲Bʣ߂��B���=�أ��NV��K�Sx��RȾ���;s_4׮&@h����k"j�`�}���u��2ﶶ�yy�H&ϓŽ�H�0�&=F�zY��t��B7�gh���N���p�&�\S{\��B�v����ԣ����G���%j��ג��������Ǒ�K~7�T���z�@�i����/ u��[�=ԮGp��&!*O�gi�R.;�ƇO/��$���H�� �:��=�r�G� �Ho[�>;�g^{��ŏ�*�N����f����^��hu�f��ֽ.�F��Ҁ4VOs���y���oz��f�] ���OD7i$�8F�+�Y��a�'��6miƷϧK��vd���%�=��	Rb<*�3��j2͈;A��.Y��/?w��}�υI�LvCw�6m d'�I	;|�K�H�R����$��hA�P�!˲w��l��*.?�IG���,Y�2����O�w���3*sz�Go�ѿ��!�Eh������k`\�D��k^���;��Q?����Z�l��(8C" �-�Q ���#���ɛ����MG�@ n)i��uN� ��&���������r�~���@	�V��op���¥G�;}6�}~�[ٝ�9M���;ӟ!��Q4)��"�C��Sl[{�`� ﳺF���:��]�\��{��40*@F����!N	8�2���>ZwVX;A�Q�~�EǇ[����_��%� �C��g�h6C�D��j�-8������3�ڸ<�2�¸���0�<�)#��$�"h�ϻml!������H��.H�̂o��`2�s�ɨ�]D��I��!F�"���Y�����N�3�m�~bc^-Y|�O`S}	��f�$� h#PB�W�o�ڐ�����)��	c
�j��6�*�'���B�G��f�����nad�(�'��Cy:_��V
����H�U�����J��O﩯��/!�%�*��G��J�:%ܤl�~"q�����I�x��������R,���>����1�[�wU��_N�/�(6S٭n�D�'�W#(?_�{��� _ϸ�8��_Y�{�n�zL�8�|y�*�������T,�HӴ����u�����x#}�s�%硤�+K���3%��5�a��v!����3��*l�L�uz4�+� ��!�@� �s��%w�e�:nmJ\1겓��4�S���BU���N�-�!�!��OP R�6s�6HF)䥨��:�[�:��Z�Ũ;����N%����`�b�1�O܂�]w���wӒ]�7I8_g�^��ʲ�s-ev���*A�xl_l��[��[�t����穹��
���.�3͛�c�sW�M�������f{xiPM�q>WZ��/F΄��Ɵ[�O4f�Q��P�v�s�b�I�}�@'�:��7�t��BM�t��>���G�Է�V9�S�3Or<Ķ�A#��.��w�a���9K�#�(�ת�a��Q7W�ώvn�VxMJ���n|����|S�?Kj�4�a���!_އ�u`����`�2Sm;>�K���l��;^�X�Mԙ!��=�au�Yq\� ([�"�E��*�#�֔��s"�q#������O���H�Y�X�X�#_DB(9�rN��$�*���.� �D�m�&Ɋ���[�}�A�}Z"�Q�r%gZbP���G��Ø�y^}oq0��V�Y�"�,k�6��*����PAGVs�Zpl1��i�5:{��z�W��h��h1��o�#|l�y2�0D��o���><�\��1ڑ�y�{�zƸ�t�,%Ǽ������(��uI��,10�T��y>��\�D���ŧ����^�^T:D�Q��67�E�0ƻ�6x[��\��2Uvϔ9ux��%�@��X�ۣqZ�l�	a~[�y��c>�'�=�=��~JT+qG�r���O�K���ȣ���`��Zv���3��IZ��8w�:78y���&8��BS����%���U>-_S�4��#z�$���8ū�,'�
���ș*�b�l�}u��������e�|�0�H���v���w����G���KS�ڈO���g��}�q���2*��x௅��V���L�r�N�fuK�������Eh��@E }06G��A���~Z��D�~(0Lm���2ٚ�z�P%%g?ٻ�{��L��^���J��`۶GqC,L�%�:�g1t�"�s;��������`�N:v͑���_��CF��c6�-��*q
��d�؉��N�%F��X���%�7b��=�_TnqK/�OF�nrs�'��H���Ȓ|����-�4�*���.�~�%���3+rd�*��6v�8����'ܛ��0�:�1� �Y�P��X~"n��+ ���9g��wuGO��L�ӿH�d�HU�Ė,Mp���#'I)X���i:���8��V���E��ut�	Wh�^�Z��Vk>�͊g=s�R��'��A���R���F�a�_���Q�|�h�n�FzH�;�$M�7?42_�����4$Ռb+������)C}´v^��<��Z�W6�E�p�pI�JY���#��%v0�ހ��$�g`G��ߚMu]|W4!$���r��.�VS�_��ߚ�`{����qh�R6�L�nf�X�Q,J�������C�Q����i}Z�8�ڋ��q95pjR�A��.�6��'�$�e	#Z�|��R� daRS�ځ_3�U�P�G.	��v$��;��W����#�$Ar>|g�Y!HU�E��	��bς�[t3ͷ��wnrx��`<�������
�_|�(	�E�ڗW-��nB'��È�ٶ#��~��±�5Ϧq�"T�L����2[��Uks�"����ۇx��-]�(���`�"t�F�1�}?��q`0I�4 �5;�U��u�%���i��i�˩�pr܊0ZU�'"!�%g�=����ycR�d[�\�:	�YKb�}��*跿[���=�P�^0p�v�r�b��bo%��Bļ�C�,R�l��d�8q��oM+�[�g/v�s?�Hs�v��C�5Gsv*�M�7�	�-�2�h�ªq{ ԛ���v��V^p}.�go�Ԁ;����OW�˚u$�4���er��"�9Ө?z�=8����o�7���̺&1�\��a��_�H��7�3̄�Uǌuά��UCM����X�/������z�kg���=XwP�����������r/GD��2��O��Ka�s0��W?��6������PO�t�Dʣ����6I_Nɖ�ӵ#�[N���N�č�:����>�(�'���cz{�oh��b����uɫI}��z�b�Ih�[M�Lf�./�ڑ,hEFKy�;�����ZG�JGEr�\��Yې��K�lذ�N-��j(����f�%�=@�.�O՗��lJ����Uz���~�+�:�"�΅u~��A���Ip�,��kaQ(����KA�8��\ćw'nrނ�����Q��2�~��?���*&�GSFn6��I.��:���%��ͤ���>.�<�|��d��+���?~D I�,�����hv.^������M5��'vޡ�S6��&�ڌ��׵��c��Я�
�!2��H܇g�A�,��u:'+� �?ֹ�{k���C��#ō5K���
�#�1/PN�X���3>]����Y�bQ�#���VK����qÞ��v�K�2k���2�	$�Ę]P̚B�!���v7��I=5�vAE�'?I���5�d ���������W��mGr��ML�gvf��!�Mm�8=5��R�ÈK��(j�/g������
�ك+�x<����Aҋ���s�44��ѥ��P��T��$�>�e��ݢ��Ğ{�f��3A¼�E�ɂ���'&=m�7cp����1o���;��	�����$v��n��P�����Y�eufUs7\T�a�fC�=	̄R��Yd#����#�b�� |䖱�c�r΢��iDBW����w �H�}�+��W7	E��8].?�f�����2��#��BGs4j)̴|BF�K$�H��Z���z[M��BP%R(�I9Q���~���O��k��B����TGԳ�ظ[�\��X�ŭ��9�
#(�T�[��k$=n'�S{�BV�NQKM�/q!O�z")���A|E�o��i��}ԧ��pZܝp'[ ��.eO����5��P]m
!�1�d;��z�qE���V���ҡ�T�7P^�Ue�̚u��6/�Я���=���rp���^ �<���pq�V+�`*{yh���/J�78�h>
v��F��KD�e�TD'�w�w�֝j���\�s���3�?h�Yфo�O��fb�@3pI��Yt�6��M[�~�ʏ+!aJ����Yʳk6�K���1�L�З�����a,�ٸ�������W��j3]�*�hDg��_�0`C�+-4
|8�,�/�r,
p_~�̵��\짬$z�.�\+!aN{��H���q����E�,h�Ƴ�h�Yٓ���b��o,�9<�*U�L�SZ?��9�[��Ө 
ܙ����]�+!oI 'N���������}�-5�i� k��"�5O0:��'��_�1�	������3N<�ω�ҊM�.ߜ��n�vfN�����r����*�3ե� B�fQ�oZv~l=�ZZ��4�y��\
�E�,9�svhg�۸�V�#w�m4��ƚ�G"�KTN�֒���9Ą1h5yU	����w����ݞ�\��l�'�M���	��!��o&�**3�)0�F�4|a�uy���̂���cGh�PE��o�x�/~��U�h�a)"���$�V�3	��ʺ�)��Jd[�s�s�����_�l͖nh!u>��uh���x���3X��VL��Y�J~uJ2�=���XBB8'K�������S>�O&:��Wx��L�F��b�Ӓ��(3��^���+���G-5^�oG����dm�+E�ѹ���'�#����sw�Pg��;�U�^�8ڋ���W������n�oI�����!�vm�������Qgi	\ֆ�2;5�?��Ȗ�kk@�z���YѶZEك���̛�ӷy�;j,!��DtlRԺ�R�:�?�>�d�ަy���^��V��ǚq?�H~�1�c(�M'O
���qbih��ɍϲ^Ղj�l1M	�(�}�ǯ<�8�1S��y��ř���^خ��{�"A�Ws�K���~��2h�������L7��4�7�O�����C'C��[�����&0p�kqM�Q�'� �<�[��$�+�>�&B;����k� �4!��2��)�vg�SG�'�P�2�:�C2X�Y���kY�J� ��}�nzW������
��X]XU�~�|O����V^�1
�G��iT����]-&��ژ�r"�4������K��r�̂�4��Z��*a[H���φ����6��q�2� e��~����7��T���Ɔ��l^���MO>����ndHȁ�4YP��Z���e�>����(�-�\'����	�IJ)E��3"��xP��ʨD��k�y�lmFå����F_#�l��nv��%�p5�4�\Xj�eZ�����:e\��"�1�Y�y����йS�|�B�&6�Ȏm�K10&��~�kF��0Ik1��}(��x�b '&�GHmT'�l#F��)�P�i�Xy\��>��_�"s�ٯW��ƾ�q�t�!6G����,���ƥ�ɦ�ܮm���3��3T-y�/��N�o�~���w��&f!�s�\�B8Q����uX��*�Q�g�y�L�ὑ֚�X�vTl��}>\H�����D<;lm�-�{^�K�%��З�F��}j�y��I=����J��[o]F �UO�	n���ѿ��ւw�����[[�9U�O��9�k�vn'�	�)=4�V�E�i���Q�z��$�vå�9�ǻ�o����� �-jށN� ���$>y��B��ݨ/�q)#$��d��Wo�Fju7���?�l+6_Qw�+&tA���-�����#h���!aV=�	7"ʌ���7�}��5�y����������J��W���nS���d�%�#%;��s:���4��$<i��]ET�3�(�����N1
��2�2���-7oQ��ƶ5��0�	kF�+�3M"ϝ�� |�}��XP�NgI�=0FsR��n�*h��y<���?"���@��j8�y9y[�z';��{c�Gk|ҰC���6V��5G����6�a��)�r�gK��9�G���Ha_Ӟ�şC��ӝ#؅b��'č
�|�s��V�e��!��a/�J�pd�h>WV '�s[>��;��d�����2R�����Ci;�H/����Rl�%Sz��c�<1�ԡwH������T���|pT/�?C�Q�`�lnOs�"����2o�7���{�B�����NS��}�¶-V�rk�zi�r5��xCQ�*Tݕ&<K0�2����<P�X���e[�C���:F��K*�c���W�5�U�YǄ����L~+@%H0Rm`%,����w#J�:���[Ѧ�͞@(��`�Җ~p�	�Ҳz���kY�C�%�0��qk��#��8\�r��ՃQ�5VJ���:��\�{������9���r8g���K���^q㒳#.3].��N��.��I�(���Fs {�A�GQ��_I]��g�"������Wceb�jfƥ���G��Ycq7�b���<�X!�`j�<��6󼠋�?�c�B	��|stW��71�����9�q������ [�&�DI�n����%�\���e�]?���.�B�x�C����t�+�-U�;6+e� 0�81�ȫ*���/k��\���7z��s�;I%�?�tr 2���1� �����9ğưZU12 ��|�q�ؘ�0�b�>5@�.���b��bw����D�ŝ�)��6�?47%�<mc>�Թb���EJA�78�Sj#4߀���4+��:��Ya£�Od�����`���z_�C�Q��}=�`c	��ז7P}QW���?�b�rũ�
���tXtK��l�O+?����0�i$�9�"敽T�>8e�G��	���}�D��;(T�6�)Y~�����@|�]gV(@�RL* ��!^%j wL�*��/����=��M	�r�p�`��z��_��R�x�p�}
�[A�S�s�L�ѧ/��XȆgW��<�Wq�;��;�at���A�y�:���샪�]�軷��ύ^'%O�`ﴔ���*=z��'BCP����F���ln�
�
^�B)A�n��	[�,<��3�T9�~#V�G��J!)Q����O�t%�c��4EX�ޫ�d 4l�s�LN�av�!����W�_u
���l���u�1�4����R��`f�m[��x<�踡���S ��gQA?!AZ�8�ߙ��L�pJe�e��i)�ݚ�>?`Í������o�	�սS����$h��xuEWG�4�om��y.L��O�MC�l�p�at����xˈZ��
	H���g)s?�ED�0�A7o�����Q��$G	�GTà�pѹl̽�5��a���DL��w��1-F�L������q+��[mH-�jm�2ʍ;n��7��)�x���}9���3k�s�t��vr!ۙ���ع���!l��W/^��x��:g�v���s��f;o�Ł�Z�UBH�s�z$�mp�h`["��������<��<$Z�\��#/M6��/OjnQ�$�l�)���wLi	�5W�iޙ�/TW
�~A�n��=�dn�Y¼,t벚�����������6�����TGBI�qԽ�*g�l*��c������5��4�j����z�Y���L�����L� p߾(���=(NG���V0ý�wǖgSsN|��me��0�+a;��9��'Q��:�E�K��y�Eׂ��d!>��\{�����LK�
.�`����g`�*��K_�*D���&[˕�X�p�;|**�>�M4���a {�o'h&I ��'�tn�W:��!�1�B�d��4W�LjϤ��Ù)��a@X.7��~�u�K?�쩁�r Eѧ����� ]�Z�q󧷩I��7	�v�`n��GHs{����<�J֞�$����q�U�[OR�B�.!����C����$���9�b�v�.���
n��z�\��vwh����~O0��Y��kx�K��"	�Lӛ��`(;�)>�~�#2#ηO �vn8Ju��/�bt҃�P>>[�B���1'�ȳ�S�2P�C�ό�p��)�Ե�(?s?�2����톨Lb����up����\6Ư��J�p�t��e�/�bR�	tD�f�`�Ex�i�&�@Ryl���Z�ማ�Y7�Qkn�?4�%��@�|�;<����)��ci�W��P�R���T������k�l��% z\eu���t]|�0X�C_������6�灎܃܀�*�O��h�,�7������Q����N�1�<�0�6N�qqH����>9�Q�hΟ|0l�^��SB߯
���A����q���&vl���o��߸�7�.w����/9�&�bp�ݒ�g��D�� }B��R�w�z����Ͼ�̴S������T�+��v����'�7#��g��dm�s޺2g2�L�J��"`�i��bު_��]�!�?)\ݵvF=�K�k�l�LrOt����g:�fPD�Y7C�̩<,g��Hƥ�U�7�7W`�c���mۛ/�J�/��A�%�UԔom~&+������F�`~�(t��ɏ�_��4�p��[dZ�����͜�������9[l��ʋ?G�4�����v�5K�#i ��~�b�6�!^^sm���,F'������j�K�XW{\?̢��Ci�r�csش��c �0��.�T�ÿI���n�V��b��V����8��e�U	��YN�T���3Q���ػtλju_8^�YX�.bj/DP�Dp�&)Tmn�[^����R�R��ϊ��F��r���	����o�_�D�3�m� �9E�³ⱳ�푸ʣP��ҖD&�j3?DK�����}î&�;����:~�څ�Țɬ��ޚ	��@5!��\��"�~¢�^zi��@\�1�&?Μ]c����vrv�_28�	D�����0҉~_K����o�`W`B�q��v���P��ю~�?��9j�	��^���>t��a�2?���7c�=����	��'�4��K��m��9׻z/�h:�eN�t���G����pl^��W�昐�������v��e��\W� �V;��]�����Wvy�����Wo��kR�S���dX���,���!k�;�kʆ�=��T�o�-��Bs�xG�t��|1i'tB��J�8���p!���:G���5m#9����EA=������L%�iW6����dwJ��߾�͝[M��[�v�S�J���m�dT]1�w��	��g�iQÆLz��[�tZ��s���{e�^�F%��?^��X46X�o�O�N��f�������R��Ѵ>�*��tx�/�:3�m{�!�Y���]\��!� Ӳk�B� ������M;L���7%H��≖Y��.�J���%ki���
ʯ4{�ޙ�A�T���40�ɥ�"�fjI��������>h�D�������9�I���Z�_y�� CwI���4-`&=q��(�P��	�Q�<�r�1���Dە��dm����p����A� �t�d��|�0uQ`N���K��<��=��&��+���Lx�*�[r��("��S�V�fw���>͸��%"��>���i�=�� 3��W��C��&)������Yk|L��}ݼX��G�$�L+%>1Q�M��W[�O%F�j�V�(����wg�[�:9��i�ϟ�A=1���4��)V��x�K�J%�@���$w���Ķ�+������������� =8��H�!?��I��YH�(s�X�?`��T�d�il��k+�\�D6����mi<��U�aB��4��cښ����m�_'Y2k�c�)}�����X�JS����&�t��b��/2��ݱ�A�D�s�XK�!蠆�A�VeqH��Z��^�� @V�~�o�ǖɿW`�]-4C;��R9UFp7Ւ����[��9¦?���V?�Y<'��T�G�(":D�:3� t�JMW
-p�h.� ո�����@��l�mf6D`�+��r���C/�ԑb]��o�W��K�1[�Z%u�ҍ߈�eN�\�yJU6��^��*6qx`+��~��Dܝ{={=��Y�e����?ؤ|�|N ��3{�>4޳��L$��p�YN����WZ����+��i��ݣ��7�>�a��dА?��m7�9��.�\�5���N��Sx5�*��K����@�c(7S��[�F�+�v��Je�mY��������O�KRv湑���j�Dp�7������o合s�%��!2�0f��-X�#)�.
"�I_��z>�^���~��8�\�|�ƿ��� L�6Q=H'ik��e	��̍���|}�>zu0֠ъ�}�{�d^��E�n�t8�jn�?p[D����u��X*T~���Ԫ:��8w���m���_d4�����K���2J��0���Z�羥�UEg�ݠ�V�g�-i�Z�⺏�\9��9}c3�=y�O?Q�ź�]A�˿g���J�Ƚ����_�d��2����p��]?�֧8�#�(����l3NVZn�D�,I.7j�+Q~V��&�>�F}}�-x7� p�.V�?���1�V�����!(yL�O)z8�K/�h��d�=��WG(��w�#t;��ĥZ�������}�Jh0��)���	�""�"�����B�<t�I�֥C0�9���+�F���h`,��pK��=ZO���f|�dK{�@�� ޤ�Sr9�;QX�u�^b:�� F����H�ŲJ�Y�Ֆ@�p���P��>n-��0�K�����nj�j�ݕU�Ѝ��r����B61/Z�!OT�*���Vn�#9GG�L��N/���T��n�`����Ȯ�%�Dm�<��gח�e�w��!B���=�Y-~�=�ٝI^�җEy��#s�i�u"7�<	�����Db�pA�Ed;I^�H3"!�Hp4&�!�ܘ1�a���A
�\�SD��{�h8��"v�-n��aC�cF� �a���b$j�i`r�AY��J�l�y�u�ׁX��ƃF	��tc�V���lu?qL��Lt�sS҃�ڟ~$1IU���4�&�H���O¦���~뵓����i'�w6��#�_��o�/�|����!�a�uY�-@��H2�L�%�`p��1u� &SP����ґ�Ĺf�d'�6�h*~Q�ݒ|~�';NC��ގ��@qA�	06���1�A�^ u��CE$�Z��-o8:}s�T��zz�p�%X������V��=R�صs�-�G�
8@�ؤx�9���z�G�y����KFl;����AT.Q�r4,_ �������W:7��0���b��[��n�� CA/�@��a:���]~*�� ��H�x�� ҥueS]aI��A�����Cy-�_�
^���T��=TA� όa�&%�V���+m�72��'ʘ'��=�6�����.&_��1`�4>Ƹ��J��m�D2�$��RdR��=���u⡸1��q����������"+,������F7
�1?Ȼ!�On��	�ʃ&�Q]���qp��!�y�<[:�'~��?��G���u�;�q٠7a
w
���Po������U���P��L�'a�n[	�܎���/|��k�a�-��p�T�o?�����3�j�~N������D�D��<�1[AI���x�7�p���-��CLj*�X 4�M�C��_q�{��V$�F���ք�W <�Á|�6O���t+��M5M-P/[UOevp�uCD�������=�z�:Y1�� �l�1�^�ݓ�Kq����Ӭ�#��vt�D$r�J�6�^7��3�F,�Op�&����P�4�E �z{F"I}�~֤@�� ���������wulY;v�Ҷ�a�����ک�x���8@.�M9RbX���O����P��ҁSf��.���el�l2�]$q��ݣ5��[�z���F��6�[O���i�ߢ&����PW�ww.9/K;6[[�`����,�N���W�6PL6�9�O�����RփF>1�+���i������8:���Eހ�V��+D1oV�u���,9��V��΄���oʦ �B\���+{���"�6�&D�^/<T0പv+����/wy.����9y��\�Q_���a���T��Հ~U`�N��11l��eScx(z���k�	�>�����8����V�f�����i�r��+������O�ۆ����8���v�\��gw{1��z��c)A����n�JF�P�p命p�6��G�]t�W���t{�|o�0��l3�y��ac�����TY84Fs���^�4����(�y�����.�D���@&[���ec�:�K��]R4`k�"|}�<�W�A�r��XF'��`3��-M����`+˪$E�������˙���jJh��5��њ)�b"���>�oC`�AO]{�UT7Y%`q�JF9�dRZ0 9<�U.��K��y=Y�O���^=�\H���r�W'-wČy���'�#�X�'7�~��[�Pf8����PLj�?�X
�e����`��#*��H���膓�0l��G#=	�fBf:�QF�%�Gf���Ȁx#j��<�v��f��.�[-�/��.�������آf�����'qZ�c�JeM�|����$:!�yU���upPD�a� 8�F�NK�H��&l~�����o���3��=Wa�7�
t+F�]ȉo��SF�����@�c����^�{b�t����g"��F��F��Ð�c�j����*.e������f�O��q�HP~���a]�5pI:E���F]���pZu��3s&T��X��SY�l�X�m��5&%pek��=�9� �	 �Dr������|� �2�C��!�6U~?��<g�D~��(�����(�����p�>7z%�|'�M3e���1^�?��z7�6�Np����qX���:�h/���1���ڑ��,��/�c��8�Q�ڇ��J��\Չ^S��P0�0|	���GRނ�(eҌ��vi�#�}���x���'�[v׷���k{�e����P;/�����p��X���!�#×��x�j~�{
�A?�׿���ݳ9 38�ϤA�_��񟺱�]�f;��\��~��#�>I�/{�+${;4.��/:7�9���h�<*�q�R�P�0��?Y��/)��+J�Q��WHr�@�W�Ȱ��?/���h���5�{�j����ozi4�#���8�iԻ�3;��4��+7%s������v�,M��(D�9�p�gL�~6ȕ��l	,��N��a�\-h�o����e�����\�^H�,�H���r�eAw^ ��l˾�H�X�XٷGn�t��gc�<���{`aw����A�憞v�~2�>gV�ib�����%�R���v��<��{�l�?�V���l���W�x^ao�èn��"O�7hP��J� -C)/.码���)�#X�����;��{;��P���#�2cj��~5إu�����%f��1'���x�c�����OdKi�ũbkɎ�#~�u�5>��H��,�R)E#T(+�[9��2�������jB��?��m�h�N��Y�B���PD�.0m{�����C�H(�<�)�Zx��o�Q�"��&�-Zxe���j}��� v}�X�uŵ��A�9@=Oo���JU���� ���0F��	����S�Pt��Y� ���߯`qi���57�w��)?�:����}G�e+���뽐��MՃ�� 'f�1��YӍ<ܿe���5s� �4������f|���E�!�s*M$q����n�6&�1�����Kd�DkC9.Doߡ���=y�@�;f��XІ�~l�2��P�ĝ(D�A������a���9��y��z#���!9�����h¥�j��a�':qlA��pCi��fsY.Ck�1�_�\�~9��=2�YIr��`
8`�ӂ=ͤޗ[ɻde��PT
���GBl�C����:��8O���ku��R��{f�\��8?!]��9��2�5DE!����i�����:�2�ʟ�,v�6h�@���i�����6������2O���?��\�}H?���$Y�l�ѐ�\Lo��Y?����\_�$|�/ϫN�[����T��M��W�{�I������R��`|�F���
cI@���n)�Z|�d�#FՄ܊S@,����OO�����Y�.��5��
կr~��â�-PW�Td
o̅�r8�,H>���d�xJ胰4��[^0>���	�V������*Z�c�K*h�Yڷ��s�ϼd�-��i�<�"E�w��c�+���O"u��ng����㸩Xw���G�����,z����_�t�No��~T�Ioz���F�Z9ny������d��M����H����xNR���Ĵ��ϣ�������������|�.;[)�w]6)�'�X��t8^RJ��E�(h-hM����]_
�(H�5�J,�\��Pg+Y��h	�J����e��ڀ��A��B�'%/Br�KL ���e�q>4����wХْ�*$Vb�4p���e�rA�j���I�/z!�~Z�/������39p�Mh!�S�<��S����	�ud�����"ݝ;]%x�[�>�7�XSsN��sF��Gǲ��c��E,�X":�W�Cb'3'Y�V�O.e@��Gn���� �D�t,�:�O��)�h�T9T���f͕-�I/+�i�:W"8�j
��?.>��XQ�H���c����e�}��ךmIp��2d�����n��5�g���A��� �FA�ͷ�$�!�y6-[��#tC6�WqC6���9 K��2�X�n�̟��W)3�jغK@#B[�>��R� z���x~������3b��ݜ�nf vj����i>ʅ�+�7�IրO����e�Bs?�5��j@ON�9�Ď��O�� ���IGyn�y�x�B�j�w�g[�;����|YP> �Y��)Dq�oCTYeC�Z��ޒy�;��j#�b�5�4�jƐ��/L�`� �H��
�EC��)z�f�V�1	�w��e�j���ք�	�z�)`T[��H=*� $���G��!ϊ�|^ڸ֔@.K<��e�7"�}*�Z�)�h�0��H���n�V[%�!��D6��*[iFq�p9�a1�E�K6��"�������ۜeI�F��.*��p�Vݠ��[7�D'�ʠ%�2I���O�e��i��W�Vu*�5*�G헓�ؘ�֡��:��Vp�A����w���_2,֐wSp6	�񺛌@
��a�R����V/���L$�=s�;:���Az:�����[:�8�R������B��N�U�@��KHt ��z�dg��:��1i���C: �tAv���16����ͫ������ك���aަz)��5�P�0Ro!�/y�*��?>Q��P�5�>c\=8��m����Gڙtl�jw���wP5[e|���Y~�q�p�I��u��J
r�I�1ٛ�l�Fl,-���u�*�KC�(�.z�lٵ��񴸐���N�F���0�N���X0D�z.�;'��^y�a� @����"� ݛ������XL�`��L�B�n,c�j�Bɵ��	���>����t5Am���'���uӴ����@)=�?, ^yh��C.R��4���v<��Ю.���[�8A��vB����j���`,�ʒ�gǍC�P����tSCA��v̆�����U�-}����AA�����RJ�_�z�YVXF�B��('[��޺竜I״�lQ�t覉t�2�ܵ*�z2�̕��)^�*r��b�E����7�È�PaA�LN�A#L?���qNsi$��\�����P0j�\X��KB�ڴ��"/AC���)S���yWN���ů�&e�`��k3�!���#�r����\��cq"�wض�Z��``�^�9�� s0���`�_�Tf w�	�V�玞��7�Lj��j��|���g^�{��'$$[��J؞��)�M��Qtk�t#�Cy�W{�0�>������_�`+�T�F�o�+�pv��*8��2$�!!#uD0vW��;�B]���y�}���	N�{gN<���yf��\��v�/w��k�6b�՚����g��;q�;r�#�����/O�Z1���<�)��\�s�ADj����Fs�B"��Q>27-�����8d�~��g������t����XEO��U��Hy�Wp>��Ѳ�B�lZϡ'�nG��DXڃ��Sٲ��ON����b�#�G?m�)�N���X�b�Yȱ�I�t�.�J�
���8��Զ���2�����5+���ڌ��ůr�x&1#xWL�K��?#�xd��Jv��9��ޏOGV-���!��kĬ��Uf�C |v�G����?B�H�������\:Y�K�5�����*��R}�:~�����V�0LO���3/���Ԫp��T]^���;��1��nv{��ʭj�@�9yR)fOv���-�Q��/��q~,�����UʀB���yHY�lm<�&��N�e)s�[�Κ����Y�
�EB�x|5����[X.V�*�g�:��Q5��؀e��G�&���'Ƒ�OD3�F`p͗ )y���J�G��3qt�fH)AT��z�?o>��q!�	l#&��2X7I��Eۏ^mW��얋��x��}���)�M�!�(@u����\T�H��g�E��fB�9Ov�G�U�V���@�X�DB���a�U�#œ5��Z*��E,3�촔�%N_�H�
�U�'ϰ%�\<3�ed0{K����MC�00?�^�`�	���T��w�R�N����[��.s?�v�8����z����B̥P����A�z�qX����������Ҁx&?�7E�i��`���o%,6頯	\�gɋC�@�z�տJ%:����p7}�f_���g��CB���	�i��&*�7Ji/a`@�>2������糦�����$��l��r*O�O�"#=�xرѠn���ZM8����X�X�Q@�`eW����_.`�0��e���PÃ�v�n��ȥ�_�Ñn�	hth�V�Y��E�hk�t�R[���C�_[VV-�Xj,yճL�.Wt
zuuNp��X�W+��Y��#�H��V�>��.8�
��n�R��#o�+��
f�a�;ث�O0žg![�d��;M_����Y���v��>�p+VIUӚ�*f�����<�Zd�cԟ�����a �MΪxO��]�k�����_S��Ұ��)7�P��yO�y^��FC"���<�������J�!�ƻ�9��e7�������N��s���z�D���n
�$X{���pA�Q��r/�ڂ�)R�sD�u�͋$iޛn=]����^�:i�s�����]*GjLJ�X|�?�F���'3�=�{i��zM����$e�P�I|q�y�j�u75�����aSL�l�K��hJ�5�A�٘��p�0��_aP:�_I�4�:��3�v#�J���X��P�91 3������X��D�#�� -�T�����/����5h��(86aT�B8|��.��3`�<��Ɣ&���R�bQZ��_�Yh�"�fz�����K*(8�.�-�˱{�6���='��2߶���#
Q�}� {g'�n���(��"�u�泘t��1w�熊��<]���Ҟu}}:�*+�!�����X^���Qd��;��2>�ȭ�P�iCd�p!u#率��$=���N��#L����p}��δdp�1T��ޘ%��0˶\\V�=����-�&.���pԳA�^��v�o?���S#���كi�8�"��-�3/� ����֪��TdWퟨ8R��bTܳ���ޢ(r��,�b�ٺ1~������ƣX�P�^3q�Y��Ƥ��Q��D�D�~�M�}-gK��}b:�H�Y5Y	�٘˞"����>im�_t&f·������,l��g�����,V;�Кq�tP�
��}>3�<�mh�������3�8"7�:B�>NY�w�9�Q�Mŉ��*�����H��ͧ
t��O(��3��|<���]��٠���sj�nO��M�O��u���7�w�eS'�⑔m���ָ����8�;p�~��1{p�I����,��=��������~��H��������f�\L+Ӈ&}zﬣ�^_ܡ/�G�v1'�X K��<A�v?�~�L�
�m�Ʉ�t��tMmc�y���j����1��B�v���=l��Y��w��0X܏0q�,�e��2�t鎦mP�>6u���)��g����ybq|��]�Jy�P}B=��7�/��!
��P��@YRQ@�Yg麽�$9Iy���:��p�z���j��H?�;��*�ͤ���Lf���%�M�u�p��ͨ�� Oj��B��B+�b*0��GX�;��a�ݭ�F@����BA�B�kKId%��*"��"t�¥�����K��L�*Io~�e�Ǻo�KD����4y�/s��_z����I[]!�A<a�$�����}U��ĎO�{������%0���dg|���(��|��VN� ��=�yzzฤ١��m�f��o��:D�|�Q:gq�Fq�F\��1=���X�*�`߇�V�k]A����^�B�����F�R+�@�A�@}� ���5��On$��?GF3�a����[��|���7pX��3���y��u�ߟ4�����]��loǳaYl��?{�������G����Z�V�w���u�ɃL�/l����OL�߈��_��EDvHg��z�G w\F#�J��U��J�}�K�A�`�?.[���i��6��^��t��h��E�Dh�OO��V��t�V�m ��CK�B?����y��hH/���<}���8�Ύ��`g��������V�\��?m-h���Ժ��(1��dm	�j�_3��>�˾f��r��.��r�P��_� ���-)_G���b%% �I��{�E�w�H�鮡�_����؝j���S)�'C��܈ �G2~Is���v}�b�T�_&7ل����&3�����p,�R:/YUN��њ
��	�`j̳�V*i'U]E��S/B����~"�A,X�H����������%���R�W�`N�߳�.t�r����B���N" 1z��C8���5{s�e�lP�c��0q��JJ�T��h�&w8�H(�\K�����6���\�����u�g=y�X&f��׺��cXc#��*����sПtu����oR��:�
q(�#!:�0KL�-�X�%9�8_jO�Z����1D��P�X������r%c�,Ȝ��:� b��p�^ڻ������lk�I���U�W�ʻ̚9�!�O����]W|�Ac^����A!�9�����N q�a����I�=�%��(@w��O2*@{20s}5���r;�>^�T��9k[�ځ(8>�
~j�,��,�}��G^٥7�0#z�r���^�!m/!r��(�Yw@�����0�Q��W]�:���
�f+s�4`���C�"?��h���gw�S��D��p�~��	֜�Y�t[葶�Ś"��a�'��"�)��f#��s`5ܶ�9��
�� ����&N5�˷A�NU�Re&;�����3g4� V�1��$�q�۬&T)�jen�~}�C�C1z"xA�q{��4Z���^Tה�prؔd}-�r<q��]�]��#�wT���Hp��fAZ}̎�KJ9�G-�F�1��Hv(l.��4#�L�!f�`њ�v҆�1b�>$yU�]�\[�bl�m�l��nO趿�Q�7��$�7�-��Ove;z�y4��n��~�0Y�V���W�����y�:�83�\k�vtV�AgYu��f7�D�F
Y���*�Zh��`{�>M�M"��J�׶��#�
�5�c֫�~��āy���3ZX5��*17f#S?N��9�,�8N
4Z�G�`�Yr�Gܲ��(o�MG�J�r���SVI:p�;(@7�P��� ɳ�B��yi�jy��D&�U�ບ{`��a?��sH�⥂� �,�eW��l��th���jw)��,�\��{WB3d B��Q�~<�~��ds�<\���.�h W[�JL�����|�(}��uRFW�2t`&	���7,�rq�*4�Q(�L�H_6u�1_(�L����ձ$�z���C��Q��)�PV�P�I����(�,�M3�_8ݘ�)�������m�|�I�-�a/��'����VWlN[ŕi|�T�	���=As�A���J) ��|��m@���oV�Q��/��V.c�/�?#���sRe"����:i�9�ʹ% ��d�ߏ�(<Q�=M����n��HBI���e�Oe�J�C})u��9�]������"y��G��W'���<K��X��s~
�O�c��n^Du�/��hb�:���K�Lj���}�CQ�;�_ٗ�R�Zه�0z�� o+�ۆ�(�pNsR��eD$��D�aO=���+ ^A����@8>�FT*�mD!� '2��c
�����[�C)>�g�j{���9�>����%s'��w$'�����@@�){΍�u�`I����s Ϳ����߄?�i������>U��]�4:���z�ynߙ���E%�Rr�"�G�&�� ���ܚ��2[��'z
�+��`�T���) rn)H�x:k��ݑ���#R:�W�b��;��:'� ������-E��=����A��c�%TI-5�d�4�+��քW�b	|�h�4�obt��k��ُX�?V��������m��dW���8oR�}�$ې�G_��S��{�;dީ�lB	|Q �`�(^b#��<�`��QVW�s\�)d4��{��O��[�z�Ј$��	�\�	.����V�>�����r�� �~�E�����������7��t (ܯ$�,lq����D���ʻ��r6�wГ�:����S�6��3�߼M�B�҅Hg�-�������m{�i��a
N�;Kn�˒�?�o1/��~�%�z�cJ�İ�������2%�	�V^8�/_e__�A���7����Л�Y*�� �J	W�ǟ�+�';k6�x�]|��|j���&�Q���M,ӮiQ<�x ;Ō
�|���p_u界w,�^]��+�UT��BQ�"�*'h����[���K��b����1��������85�8\��F���r�ݎ%P��F��r�M-���[�#��\����=�q3�ܲ�.�J�QR�k�o{2z�'`�	a���| h��2v�����3��-r�E�������J��~���(#m0�:=��3O� lV7���/�:�pW���T|p����T��D�Ձ�U� �Գ��BC�ZL[��աh%��� ��!r��^miKW�Dlt���k����ŝ/S���$�"h���#B0[���	���%�2յ ������oi�px�J��q=:���i��tt���,��:�xiϖ!�˚���������˸����e�IhB6@dX��gt�P��J�˗U��z|&�=�n��6E\��N���8���jP#5r+5�����d4G�ڵ�W+�m!ߣ�"���n�m��~<��+�|8y�����ܽu���p8�>U��a�v��0!�.mC�û����7��l�_���P��|�-�w�[i=�l�l�o��D�Ǆ,%�	�8�;��;-���;',�CD�
0�w�Ko�,�>'��h%�bd��4hQ��!����j�T��9�&���w��/ρ������2�E����u{i��~%<ד�)��B���j%bg�4��傔��l��իi�����r�I_�c
~��\5c���� �w��ʓ�@f�9kK΃���hLU�b.'J��W�T�����zZl���W6�F����b4�F��0��M&@�r�f����Ҍ+�Ҽ"���eT�	�� _˹N�f�&y�Y,*ϟ-:Œ7�M'��9�+���ܑ�e�3t'˞x���|�������P���al���03���w_�����7f3DO��x!R�B;fg�����箮8��hY�QE�vx�<�`�w��11ʹ8�yCA^��C����wDr��~cL��� �o>�kl^��W���0����
�"�<��i��TZ�ƷR�%`��nr��t�X2\·����{�������Ε,5ߍ��V���%	Ѓ����HR��ݘt�Yv%���D�����NIU�����Ψ�c�6��kp� QOp:2�AV���^_P�X�e��qv���B�B"뎔:8=����-b��r��F�E>�"G��=V��>�e��Y�h����}r��Ol�٬�K����>#��q���K&����/OI��Ʀ)�Y��A-��S�I\�G�N-��g�I/����,��V��&d����k�����.}��"%iA섔}���d��}V%�]?6�w��o�%�����-�|��������7N<^G��l,;Y�i�`�I�{��~���*,�=���q���
�+�X���XCq~m�|�r�� �6��"FJ�dW�9�F�#Y�lV^#��	�V����P�=Ĩc�K7�4L#�i�hU
-W(����Է�6MS)���[� �lV�����<�b��X���ֹ0!����`:���P�m������U�de��~��t��;R��q���d���	`kR��y$K;��ƌf*1���`n��c�-1�FQ���$�«|z��
���+�X�i ���ܼdR�d�l�M��i��ĕ�u�Y�^���I�!�U��͜�0��,;��@d�F>K�^��!�_g� �/@Ҫ�S�I��K�-"_�&���UqIk�er �l�����K{��R5��_��rț�N� ����=k<���}�7��7�aJ'y*Ζ��ҁG�ɽ�[)C������̡f�\�.Lk��oBO�|���/I1=[4XP3`����/�V�N�<��U��ߣ���;,L䶳�l���4sL�䧥g&����1���V��=�P1z��r�/$����-<<$�9`�:^��lǙ�A�Z�e���O�鮯���{�c	���z�,�U������`D'��Z03PH6��@�ަ�%Ј���gB���&b�$�{�՚��9�;?|j��v(�G���gn�U����.�D;�cy\�N��oE��܅'sڨ�
q;����d-4Tk9;���uE��d��:�p9�< O`YW�b�hW�/��%	�ͬ��Ӭ2('�&�{a���=�-��eޮ�������cw�R�H]�NUvm��g�ӈ�����)9�d�ޑ�;�
u���*�/��o�8$��'��|��A ۖzJ�w����g��QJ�F��	���=��w �T"���+��Ȇo?��ٳ|:ߋi�m5������js�������M���t�q�*�<����p�������8���+Ȩ(���b�C�<�k�wOf%�)vu*h�����DY ��G������9N�oq��ر�$q��}��Z�m�d[�&�5%tjc��a�`���jA��)�ޣ0$��\�)�m�����s{�{F���2G��Ŝ&��Z8R��$ĩ�:��z�V�R�L���c�l-*�$������ ,��@�}����W�U(an���|�9F��Q�0ཛ��ݨ��C"#4 �O!��w�߰�(v���l��� /ǻ�[K��]�������"����lf/���@O�������Sa��p :���g?�����6Rzl�T�d`Ar')V`/c��"���-�ez��R�;�)�GNH��@(�ŷi�̯?�a�bc�O�zj��q��:2�����>N�}�	���'<V��$y\���2� �����J5�)��R	����4��;����!�yQ �Z6pܣ��t����8 N
��d��{�����4��N����Wu�L'��t��0��&����ȱs�zK�Y=ok�0��m@��N8t��`���I�˭su2BB�Ԏ�/��-}(���X!fs��K���im��F|�н�q�V�N�ڲ��v�����`���;U\!XM9�|F�G �fΗ�X�$Z�+d
�"f�Ɋ�(����zxz���[5^6�m���.��I��^�b(��^��
�M��F6+�I�ZD"��TbH]�	���sI4 n��|���4pa=�������F�"�)4�1kqTƫΰ{����Ҋq����>Dw����̾/	����gv�<�:M��y@�]�t��1e��B��[�(����t橣��KȌ�1��܏����c�2�� �c��?E��n#�MZ(U�y�d�J�A�����_�	@����#�襓�ݤx��-������ �UO�\�9�N>��a#���-�ܱ�;8��9�8r͚~#�ӭ9�$Ne�8��ֲ
���ڸ���e��g8?��/ ��G�CSL!��T��k-�1L,]��t���F��{�J�
�{�T�_ZJm�@~�k��`�����Y.c��U�i��K��?IH���y,4 ;-�����N��z���0A�F�3y�;4��uj?����Auw8D�(��nT�+I�H���6G�f���fjJͣN˯c����d���>�bKp��J�\XP&��� ��9�z���1@��� �I�	���ݕ�E/�
c�>�?�<Cr�p�G�~y�7�����]sp0�I����'k��1����
;�=��f ���ڧ�nv3Ds��J���}3�޲d����P��,r�婬��_yH<xt�
�k&.�>�D�E�B���L+w¼$��,eͼ��s�L���W+�o�7<�m�x5�� �/|˥��Y�M㈳</3�����U8�J�+WvE�o7�����^L;���V_"f5���tjw��;�r%���*�M��'G#K{�|�����x}� �ؒ����m̜d#���;۽����/u������jG�u9œ��c�c�f��#��+oT�!�i#�%�/��4r�z֮�w�EK��ʃSTܖ^iie�j	'�o�5݅dx��"���UG6E�"�t��ID#xH�`^w��I�9�BoO��Q�*���p[绀}���F�L!��
g �8J��t��|�	 z+L�~�\�b���� ؘΞ���&�4��vg��ւn�Y���2��у�\�n�i�-�^u�`��+�C��S�tM���{��?��0����W�&z_�igb@���=�k�9�RIof<Ya�������1�Ӗ4��"�Q�0��mujQ�3vsJ�}Z�U��g��OJ^(yk�$)�BT�~��]T�I�G��l:j�vF��$����#7���Q�ƙ����?gQW��}�C/�\�tR��6jV�o`��;��
�Ծ�&@m�Qxj�=���h}�r39h��L��d��uYԴO�w�_��.�3����@~o�+�^澤�X���nq��O`�E��U�J�/H�6-�aNI�vF#R��f�5��=�pp8�>#�dDW>������m�	!۲0h�S�.=8]Jq~�LOa%_=�2�/��k+��b������@=5��fʤ�M���S�6���kb�
��V��Ч7�	6��b�e��z�;�탓��i�����g}[eIa�t/T�S}�=� �*��i�&�p�fkQpJj\p1����q����߻X�Lg���p�}j�?H#��<O��x��ۭP�D�ai�s�@��\ԙ፵���$F �Fs���	�h���>t0�;ZC���}��w7��cS�ZCs���aP�X[���D�CP3�":�`��IƵ�T{/��e�> �#H�Ҧ?=�\��a����ԭ��'9�WK�����o�O��pN�ݹOTB����7�e���zhV��q�x�3�|�GH���=�S ��	�����d��Հo��j��]:��<s���u��yaFSf��l�j�[���s����q�ϣͬ�P\5\�f�Ye��0���:��K��U�D�u*g
�I*%�j#��`�?�1ū�c�-��󔏐D�̻9�J���Q~���Ӆ�jl��0C��y���,��^�u�7ݒ�CܸܡP�M^��ķ��\������s'��A9���V =w�xY��"D��D�e��l�_P'��3:�#Yv.Z�&m���#�,?�(j�|ϷJ�֌
W
wk ]�C,�0i@2���U1�̒;�g�o�y4��#�?Y_MW��J��G�s�|`���x�^�� �3�z��25��-â�!�T�B<vY�J�ްu�3# ��I���ZVB�s�D����PUrPQ���:܅腅#5��D�T�2�֌8�0i��Q���[ ���T3�Y��N���L�8�D);�QY\����9�;���(�QQaa�9󟑚�p8�X���:nO�8��b3�l@�>raew����3Q�L�K���D��s��q�ԁc�,9/n�b��2#	:���K.V5������w��=�4Sp�o�f�#��cDٴ>�/�������b֞;1p��8�x ��G�BG�Q'v���C5K'����������zN}�fAV����u��Bx���n)L�k�^'bSk�J��N��,�c�,����W�"1�P�Mꨅr������R0!�ZEe�|�UTQ@�Su�\i�A3H��?Z�qX��?1_��0h�s1����NŦ�a)k����؂78fP~�dgO�}��|�:Ƃ��5���C�W��R��	�\�uBdNگ�7�]���P��&�ϔF�x�{n�������0� ~��^d�#]�)x.����)��{�A�Q��l:J~�b��:K��&�� N���	�)��~�fX����]H�!o��Q�8��_~x�͢'�4J#���H�� �K�WLP���G��$��-��o���>@=e1a�@o}D���kF���Es��TaB���R(0ilc�)v���˪g�3����G{�X[ �[�W�_,��*m"!��#����r?c3���͊��8���t�Xv�w�ԺR�ȤغݛZ7��If�Z�'	�t-��f�]�2Z�P�b������Qs�S�'�[w��M!M���/�)U��a3�"��g3-���~L�J�?�2���S�n�L+1πP�+7k	����:�^�~��S;oz����Q���C��]�����#|S~�W5p�4?�Ln���ݬNQ�H�!g6�y��<���[6�4��tKQg���l����/,`����@aqe���@$�s��s���p���?��{	K@ǡz=�F�/D�gg��ydF��UU8t��B�]��i)~߀����	�����D87�PrPj��Ê���0?ҕ^�v�Ն���;5hb�2WV�灞�~�7�L����s�hP"	����$K�������\���8#�[��T��A78��͋������0���dp��ۇ�v��Ď'�{Z���\ ݯƱ@ՀB���]�u3��\��w�)��Z��t* id9�<����S�V��c�2������^&T=�J3B��<E�.��RU�J���H��)����pxu �7p����#�aE_��Y�Ĭ�'��H�;"J�8�-i$:���� sGf�g����`M+�BӤ�~o в%~WI��0�N���):s	�o�r�o DJ�o��g}%�r�0.cl[礕��@��^1l���,�" �9j��d���T�o��{̀@HS���s�O
	��cr����?����@�d&��^�
8|��&x��d`=3nƘ��+xs,^��M��ѓ�v?;�`�	��A�G��:o�O�;t��ً���W`mm4 �P侀��qv2m�]iv�\+@H�G.�Hw����̅ڰ�Td����u��'�6`��V+��+�[��p�9�шԬ���'I[�~�TR��d�<Z�0VL����+��B�(����\�P������Kr�ړ[k�^u$�}���^��4}�s=��5O�nb�i��f�.P��L����M��f������P�Iu����LIc|�ENN/v��n .?��h��s���n�RZ>�������fޕ��+��fV�w~ʧ�CW�n�sm�^�"~�8�؏=,\�ٙ�⵶����H������q����q���꼛/�!��"f fqWd��	w�l�o�`��i��Itv�o�ƙ�����t��	a��R2]:���Qcvl�n)(&(�Q��Z6��cQ�4eZ�^����2YΛ=�y�O��nC�i��L��HT�m���"-��X��ꗧ^E�t�Wr�|�(���"V<[��I���iY�zʃm�\`��T�d-C.l��ި��snk�q��3@���P'U�rC���Z���cI<Xc9)��|�0.�@��L�����x���³����f���S�2����yˍ2�1��V���1�^ϰ���R_�i�]��_'�F��9�j��>�f�N�yle>�����U3{�*���6r������r� @�f�B@4LN���jg���D��D�h.~����
�b��
OފB'~��H����2e�M7�&w��L�f,���s.�W��i�
�C��	�����P�{����! ��1��u~�R,����
���i�[� ���m����:�Q���,m�|ͤ[�d���6�S�7�G�����5���+�C�\������Q?���zs�$��<�3��o;��~�	��=�r�������_�
ÁK����<mu����Tx7��A�b��#�E0i�Zɇ�V){����2�V�v}��+dƲ�c�RK�lL��U��Cԇ��s���5�}!��l�`%����1��%}��3�i1X�kav7���
��������A�;5![7cȽ�_I���ك�#l�s]�d�˻3�飅�F���c�(��&3�����J���JaC�����,6ݫ}B��3�ƞ;1�mN�M�$�(�i������!�k�b�Js��54��?���̪NA[�:"����4�1�W�����C����\d�k7�^�������!��{79\�in�'(�F�7���@���tn�]gx�e �E�b��8�ZA��_�ͥߗ�>��� 	d}$�^�;��Hr7�t����'�=bJ�W�;o��c�<�+�K�����j�t������뽓~�e��#�}W�}�����%�]^���^�:��a��BZj.������m2_�N�K'�a1�]����>��"��(i���5N��$f��vA�y��VD:?�	h��%��P�A�6�F�-�~��dO2��W�~�%���`0:�H)P:-kp��}v�m�K���evO�+�(��w\Ph��o�z��`�ڨ��v��C����$��Ff&�1S�n(�Rb׫�ѯ��J����A�(>�.Otw�':�i���U�.�y� _����j�=U��.@"9{Vs�g �%1�&-[���_�|%�_l+���Ő]۸^#��[('T98⃶u8r2v���?�_E��3.�E
3![QK���5Nɴ�� ��+1���RR�[lv�B�M�d�T4B%�.nJޘʚ�a�ڽ� �1���?\W�;�*�N6�L�ARJ�I�>ӵt5�*���r�Akk�'��<1�k�F37��isu��K������H`�^��a�f^3��T\���3�W�O@<��E��]�����kQ#���V��.�2���%�BT֌�<�aUh�"ML��M�m���j�>ӻ�c��X�������[[��~,0�)���F<�ґfY0}K��f=�iT�G��`+����笽�W�-��h� �����_3�HC��.JйQ�DF��(�
����C�~�'�6e�&�/8�Y/;H�v�
/�Y�CP���aU��5lӳΟ�+�C�9b�lH�� �	�qS
����l;)�r��*��U�!7͋<����э�0!q��P���ܷ�eyXI��D���A�Bi��0�&pgO��	t�RF��P�.�G��Fe�k�L=۠^ɶ�����A�;`�+�� ����X��~�5�d��Pwdi5մ���'d��v�i�h�Q�q>�⵴$�a��傮�^2�E1'��<��m����)��y��ю��x%D��eUl��{"h�0S$R�B-$hP;� 0��Bkղe�G�&��s��N���#�Z��6����k�GjHٽ϶>2�[���	Q�Ay���98�l	���Z,�*���!�Z���A���<f���ؤc�~@IJ�^�qƢ̽\`��lC�to�_��0�6����ۣ=LgЂ���l����@�v�<@$_���[��m��f�Ḡ9�#��~ c��\D��e-���"�1�x.���603����2̀ۻ�D�mᯂ	�!�g��@���/��F\pjb|��LW���4���g�F�<���g�n7HcT�����3�/���X�����1f��"xLqW��01^6��JQ9��+p�r�$���k���^�k��v�Z����"	ߏ�Dj"�K���i�?�ѭ�C��ۋJG9o´cvg����.�lO��{�j�˄�2S��)^��{
�΅�j���]isT�d�$]'h���ҀuW����qK��[����VMtH�g���_�׎���(��Z_v�!��s�e��X��u��X���(|�X3}�;ǥ�]�5��`H��هH+��#�����ݍ���U������)Ê3�Y�7'޺K��*��s.L7�r��e�6����_�0����� �r�����n���6���ޤ@��t r�,����*t�7�>C��o|*�e���RZ ��cD���@
�锻�!�C���e�q�k�P���ܸ(-�n��>�R���Rq�r�&��o�:�O|�H�Z�}�M8(����l�Ksq��͜�^N���Ceq�a��+���&5�H�α�8G8���"�R���H���F:i�Aq�+Ǒ��r��f^ͣ�<���F
B
�?>Q[,�0d�(P%��mp&������{ߛe��ʏ�޻!R���w= �?�g���U�Y���t�T��ka��q�aNX��?���\'^Y�Ď�5�J���j���WԞp�LcGH{K� �Aq���H��H_���^F.���m��>���ڂ9��Z �����Ǌ�oO��ʕ�Dr�M^���9
���a���vI���"����Ӱ&��`���^���w%6��9�{������CD;�B&���Kw�v�sL9H�n���Κ�����Wd-��A��Q.�{���c�T�2Ks,87��eL����V����E�߯	�gʨ�Κ��{]���LV��w�@GI60��ɱ@�%U�s�4nM��aL�^k*����\��l�a���A�k�K�7�k ��Y4�t���e�C���y��aΎ��{�"ѣ��t@�<.��e���&8p�6��n̢��a��#<C��H[6��P����(����s���>6DX���Z���} ��)�K�0�9�����E�=�6���WAe@���vq�%���`3xA%���N^�+''g.��K�$=��5c��A�(�&$��*�~MB]@�)�*�� t'���D��uF�Ȍ�1��D�dl��4���m�ROO���xMȼ\�t�z�{����0`)�/h��2�^���X�jF��X?�����"yNO~����9���^�Ե�5�`���?1�_�`��g���+̿�Mh�'�A�l_]T!!c��.��(�?B��?M▰^+3�Ʊ=C�[z~7k�x�����"%��a��K���u&�h����U�X��{'BZ}!����:J_N�)
	i"�Ӂ#|�]ꚦ�|S��f=.3 i�H`��΀"sbrS���z���(PX7C��8v�Ti���x�J���zVP={��N8[1������h��	}[�Z�=�XTx���	�{5B�z2a��Y��%W>�,'Y0_{)f(Fִ"㖛C�e�*wv.���ͩ@Mx�A`�@���
�x)�j�[�]���r��|bq��w�%�����uU�=9~���X<�k�~C>��,��?@����ա[%�-������F|��W���~g�I����=oN�O�U@����D�*2��}B6��?�"D���Q��Gv`�UN�w�T͠x=!O����i(��6�^��2�Gi��u/b�%a���w��Ѧgb<c>�a�{� :�P=Q]��F�K).��`c���9��i� =@hnN�(e�;��ĺ~F�� ZR
!Σ���I��^�|�F�'��{��}/�Z�C�f�r��(~Am������_NG#�6����c�g�}��A�r��{iy:�27&`U�2y�+1�&�WR񍻇�V �5�����&6 .�����B��b�;T`�ժ>�a��_s4R���`5vЁ�Z�\���%�i��* �|7g��i�S$�!�̼m��-my��eU��vJ�A�lJ���g����&��_����-hg
�!��'�m��Գ�+E)��;V�y7Rz�L���R�^�~�^� ����� �������0w�":�/� [n��[3�9����T�e$��R�����ܲ��^���֢%��9L��?��6b\��ǣ����2�UэQ�F�:mp�ysj'�,�ݸX�Ҷ*��^��Ht���F�d:�@V��hC勎�|w[��k�B�sǤr?�ӵ��{C�&���*%�OXO�o��pP�����o�Jc�Șvg��О�HM������l�Z[�r.ǧ�js��օ߇����rch���p�O��� Fm5��B|���J���E�k�K�RW��2�H��u[Y�u�s�#W{g�����/[F����~7f�2İb)]q;����н�v�5S`Z����-HOsJ3�Q�*�_���D������v�苬FCU�G��y��^>Q�����jr�TK�U�?j�q�m�z��U��"^DC��ӫj�[����f�L�G��Lt���n�(�m��Y-�@���B����|�_oHL�S��jF�s�>�(����E��
4wx�v>*,l��z�ybA�=}������V�nO@%r�A$k���KN�S�$��3�;=o��d��)	s�X��\������),	C���F@R�Y�O�0���9�f�o��%D�}x�!+�ɫh�W���^����.��klg�no4�-��b�@'J���\ft��૬�E|2g��S�e�g�Z�3���O�پ$���X�8;�$�����-����7c����7���k��-�?8m�h�����AX<�-�墏��f���!������S@�|K���欠5;���^�
��(�X���W�?ùlXk�a�y:��0���z��fF���1f�ĉ��@�R�(`���	�5�'c����==���ǝC(�G"���)��t`��4oq-3[{�zex0��=Е�ս�	�&�`�����q��(-���YxW�kAK3��/6~�,���7WF|%��]t�h������w�}�n�te�\�88�K���os�iQ�^s�t;��k㯇��(��}>"!�W�;���)X_��&��[M���x�#>$3�O���D5�4ajB[? ���lim{��T,��}s�c�bբ�y�	��nh���]f%C��N,�%^E�ׇH��.V@�9�8���^!Y�]te���lx(�͙���y��v^2����^.�����J���.� x��3B�p* 4��A�H��X&�!��&�����*}�q��%l�j����P�!sX�W�V�!A� �����]@f��i���i�*`	qQ�ޙ��1;�\���=��&n�������$��7���Ǧ�݆"�:Ľ�F�Lb��TiR�����/C5nƮ�˲�~��Uu�~⼨��d�y�J�U�Ζ�;<Oz��&��Ze	�v��y���R,�B��ܩv�%��ޅ�-�&���Vhk��_Pv�Κj�}�Ya�*�N�,{]!�ܻ�MT���#F�Nz^�q�T0Œ��,��6�>]+;rC�-���W���M��,�v���XU�aL�p�z>׹\�	sʮUe��.Dg���j]&�E1�BE��^�jrdк��^)ݱ����zJ�B��tXG}������&���[�$���i�+��/L���?|f-��|.�Y@O���"�|��*�ܥd��]Ω�������`� q���,��.����چ�#��?Gr�?�#~����2�PeKzF,�R)��!OZo���ݕ�z~�DW["�V���9>{]9ڇ��^��>�%�m��唦$����ϭ;�\^ft9W��ok�f�h�m����ښl�M�מ�M�i~d��RNf���Z*�
�{�����,�g��G�u뚊7"��l��)��g�1xwQ�1�F2�%�J�\ci�,P?�URR7b.����Pa����k�b�P�M:Ұ��~�������^5��������w�L2�?�����}��������������V�cӑ{��д{M�Q��L3�؝�J ����=�����|u��l���u,����h����z̘�S�
��B^k5P�T��-�k��f&^1��i������x�v :�Ķa����7,���1����ϙF���u��u������p��'ep��i�ʟp�'9x���6��X�Vp�r+��kt�5����H�y��g�`�F�\��i�B�GJ���-�璭���g3�*����A�՗�W��֔�i+of_��I�K�BW.kB=о0�9@���e���fn_���z�R�[�k�9	%�����8A�d�r�~��#���IIMp���HV|���Zɬ�Qf;����Jh.Z_>k��:Ӝ-°E�Z��.�_<x�5y��>	!�N��'��:o1[[���藣�K�Et�@7���s���V���7�ZY cQ���pZs�Ehm}�z���LRN�Ss��ً+u�/TQ���JP��/F|�Y7^D8>Wi.�\fa9�U[D%'!sqpUd:?+L�Q�P�<��)` ���1Ke�Z"�M[�q(JNt�g�tL:P�Ys�<g�}�����%�G��� a�9#�8��1��4�ZK	|E��%a��t���VS��5��X7[f>p=w}L;��M��C-S�<t2�2@��1�\�5��]�IH�i�*[ڵ�Fc��yb��k�4f
�@D �����%&P��+��A�ؚlb�r,&w��.�d�l�~zb�	%#��11�Q���)������6���-+2/c�͗mQT�|�cL�_>;�[�x����K3&�P��Ey?os޷��[���8��{�S y][+����녟�DD�lb%�S���D;҃P
v����iavk�c���ٞt?��\c�����%�rO���y�̵Uo̄h\�p ��r��?<3K(���ܽ'����^��}'T��ߴs���|��	��@k�������B=E���H,.C�Y�������
���V��j��g���w��%!^��Dу�<A.��3H��B�4Ze�1�=�5�Ok��.%��Q�'oP1<�"���z7Q�[(�Gw��п/���1��#|QVعW�R��1�x�8�x�|ߌrv��Elm!̦�})&��~������԰�p�3M��x��H~�f\��\�21vJD�(]��ѱ�lX����Y�	0�A�pkMy*���,gVm��Ј^��c���8�t�7�h���3��^�ӥ�-T��@��Vq~������F�>�w��͹��۠��N[WL>��&&Ѵ����,y�:
����>�F�1��R��*i���X��H�𔷖���j��w�s�bz$��{7bHy�z�����t(5H�B*�B/��u6-�'칪�k���ͅy�wRp��X�Y/u�N�<��_�M5};�%pS#I�"-���5Sjȑ���Y�X�^X��~ݳ�����BY\�Oe'`���v�?�Z�j�Y$psa
r��C7.�~�Cw����3��@��꘹y�,�,��&tTy7�j|��	��%i����}0���J�uƏ��΅��ZSWc��<�<���R{pV]8��H�kR!�࿡I�@�n��Ħ�LӢp��og���68�y_:�
OX���)�(OY�v�m)k��VO02sĶ!H�t�Q��	�S�7�1u~�����ed����I(h'"�H�� 6ǰw�P�����B%Bݱ�5�n#U�n���Z���/�p������� �H��#�V�>�o��P[���'�~�Rs�5�>�E���`���0琵�jW;�c�FO�@V�:�Rb,�*-d��$(��'����Vq2u��^!��V�9�F�Ɔ�B2rMo��L��t�J�-�{�݇Tg1Q�$����^2�МڬFh)��責�{����۾e���+���ES�8?���?Y��T�K8� x�[�~��ͨ�\��~q�&�^�C]��eV
�_Q��=�Vz/2 �v����9v)�da1���� �~�2��p�vȩ�E�%�� f��%:7��_��h��2C͏@My�9�� P�(�<���]#'I�N��8�����M����D�h��Y5O��p�Q	'��:e��_��f���9RLy��J}�v�Y�Hu�3m�lׯi���Ϊ;�m2�P���@׮P���u$O
Js@���:��U���ڔ
�ȗ��s4�@�?Ħ!d�&�n������+�~��x?��\9����� �ZV�6?���u��]�����#wy��_��}��<��ve��e��q�ùZ?�6�'����_�Fs_`��@v^��^id^�C���ˀ����|���y\��֩��L,t/���;��h�嶱3�o���P�c>$}��P��%|OD�X���8=W��&�ۙ�X
;�΅cW�<�e��'7����P"����Qi��KհcصB�u�n�Px�,�/�"�<��1��F�Xk��x&g�b5��_�ej}�þa+�ýY�U`�eh�d�51Ռ%T��z0*G��A�!�zi�@��D�Rr��23��)Dv��uA�2y���|����
��fp��i�
�_[��e/ؖM��=e���<������A���`�K�����{Sp��C�\,�\Ԫd�x8�G%�� ��l�yY ��جF_����5��"� � &�B�?eq����y�����v��IJs�w0�i��������,�mGm���;�P�P���y��':��Rn��e��$���7�}�
�3���M�T/8+����7�I+T ��v>�+�Xx�>I0�ղ!Җ���Z�g�Ѧ�&Ը����X�ؗH���F�+O$TQ

ү�QQ�W<A݈A7l�q1K�tw�@���~������>�S1�[�^?���26[ Y��z�i��z��Xl{���\��܉���� ���.vpb�=�3��kK�=��q �a�Ҭ�:cP�@+�D,�g�����v����&Z����p+�q)� (Ϗ3fMK	�.xrC:@/BV5�t���m��Νۍ-����Sf	ܘ�/�������s�g!��F��='e��`��m ���FL�W���%I8JO\;���\��޵��ڷ�,���'�_��,ܫ	bY47�G���N�\7�8�����0BF�8��kO�>��x��dmy
������_�\�S>�o�#��E(K��P{�L�3s'h���ſ\+�ߪ[�Z�԰lR�9��Ds���)�a]a^�m����D����Vor4b:�w��� ������%b|ĶV��(����^�̋������&t_}O���.�X�7�ad���i�xw����������Ɖ���3�bP�kȊ؁�f�Mu�|dVS�P��J�	ث����yϸ�Ѡ��"��rf�<�g�>�&�B�i'�1�?�O�+ J~��K�ß��s	����̐;��	��s�V��ӷs�_h��:��u�d�aF0���I���(�l��|��-�nM���6���z~L�ȶ�jmYyU�C4a:a��/���]q�G�a���-���ʼZ�ӒX�O}l%s!9��
�����y^�N4�ŸPWH�Gy�j��n��ȓ_����s��Y��9���a
��秋GKAU%���ˊ��A"%f|�i{�}�����Q7E�����0A��+JH�OX��������
⭛��L&W��uu��|��2c�&@G�E��NKr�ɛt�Am4���L��da�$���E�мK��Y��mJK���T�f�ОȠ?����E$������kV�oC�W Pp�����"^��>����A��A�ݦ}��E`ҷ��U�_/�9C�ݰ���n�Ԇ4�u�[���Zr���wb }ba Q8(N�^�(������b��]����BC7� ��y�����g�A˄�����6z��L����{��V���S+BM�@<�63@L�w��h ���Œ|XUv.{d%�T4�4"g�Į��%Cu=��EnT\��obV�`.#��5���G:,���{z)��ol�S��.��oB�C_`,������h��dv�7�~�]^�F~6��~lz��}�Ě�&ȦI~\��5��M��d�Z뫩�m��5����lU�Y#�I���
g�#�b;ۜ����#��~Z�<$@b���:SA{j��U*e�~�� ������&y;H��'�O��]���/d[4����=@�N`��%�j�o�B.>}w;���kσ��!a�q?>��*$��޴V��m�I���X�# ��Fk�\[�Ϣ�S%E!���i �NI�����JBM2A����ͣ�N�����%
ξ�����2�\ږ*�p�?ay?�h{0!#4�eQ��Q�N�<�m���x�Ndާ��+����mm���a�����aYuMZ���iy�+s��U�n�;n}���Z#L�8D�k�2�*OQ}���V��P*] ϐC!����D��G#fʴ�I�;�D�X�%��ő�@�&WU���K��ҥt՗��h�0F����	ё�O�s��W��C��y�Rt>����!OD�ƃݹ!d^�c^��t��v�X��S���kE3q�������D3�H̝x1(����G�z�'��� G�7�p�U�E��4����4�V��A�i��D�hf�+&��ԉӷ]�i�W��F�Q������I��,�q���?����`��N0�\�^�^>T�h7���(�ƛ����S�y��~�As�Z{=n���N%: ����r9�?�񤄉u�a-�{�)�A��>H[�1��f��'V��7f֊��+��Z=|5�zB`P��̛�a���l4�Z:�v�Q';RC��|��!��<��/8n�}���<�Xۧ��LJ��9�+8���t��
�W�!�����S(���Ѷ�ٮuZ
���DM�����G��i�+�0a�Й����������>�x$}���1"Bp%��v�-MD����
����J8y/ނ��"-�)lpw+���hޕkI�yH��j��k�n��n�x7��� #}�ִi�,{8�a?V#�2�df��CD\9�M�lC~E�Ik�mȀ��|����#}/!�m_V���S��$c�JJ�5���>N5����c6K�����!���%���cP����h�J���~��E��T7�����ZI�I�ʣ3b��{6��)(/�S9y�P0k+����7�z��<�k��_��9�pz��=뮷W�H��2c�tC�V4Ws^���h�Lv3�P���x�f�֖�=i��^0�Z�n	��v�ڝ���)E�n�W5��g��QhE|9�����5�S�.���YC@�����r�,T���׈�!���;�"`�JRp������jŎ]j*�=9�H��⋇����'�#=�J�2hܷ.�x��#Z���ٺ��]E�N8tLxjӨ���F��ś��d =�H������p*V�=���pl�������f�BŹ�H�/�l�������zi�+��0�����/jݚa����J��������9�7p� I�O*s�6T9D�&�ڔ�e	����A����$��Ŀ6�u�Yq���f��>7�m���O��s��R3�룇�'�tu�u/��V��<�NY8!|���P��fC-��"���̐���aF'1���-ZQZ-T[$����otV�!@����^<�^(��]�w�x=Dd�x��E�o�M�VF���*Iۺ������}�.>�9�}ˍ��&�8�p�x�.�`���}6��U���{}C���f�
�g�ҢG g�t�+�\}l$��0������rpf[s�k�Z�����Y�����sNক���� rj�2Ew7�l}���ҳ�Z�{�p�H����/W"���A
��a��w Ql�eDs��bm"�zr������h�ȫ�w��xG��͋L2F6��Eϙ�b��V�']/�	�Cl���ٳN�o���ï��H�8�R5�S�Š�i�6���c�f[qC��LEu*?�s%j/8*���X��_��SG~�nR-����U�8�z�+X��M'#V�娱',��R(߾[�u�WF6�߫W_D$��f�!�5L��Lo ���	Af��.�~���0����i�(�����q+H��n~)��{�����^�C����D��N^�j�I���">
l��E���\�D�H8$�N����x��ދT����w'1�悃�@�Ř"h��kH�ٗW5�eG�Y�����P�G)E�i����[�?Œ��`w{�)*�r�k_Ny@���lo0�N�Q@d��s9�������AC�$4 OT����qꊄ�zHp�~���x�%Y����̖��&��#�;ža.����{��Ll���J�`	�ҵH�PZ�x�T�a��L9��p.C H�@���:]@(��fCeuOH	 h�3H3�l�6���#Td#u8-��xb4��y�3��@%0����K�f������(��7���eK�BJ��/vLl�Tk)=�`+��NZaz� 8yw=��p��0���q�^�X�䉤(<�g~�?�_�� =���G!`ЕBD=��zL���LO�������AC�,�=&ǣ���I|��U�vv3���o>[�gC1�l��ȾAhW�݌\&鉉ty���#�æ�c�7Q�h�7-i�O���n��dT�O�Ϝ��p�T�/�V5u�A�|��Q0���M���d�ܖ&��F�������MCɆ�Lh�=�������>N�Ok���_����_	���n��,<�sm��:o)��F^J4���Y"�鸛zxV�*4�&��$��'�+7�cR n=.�n�#��k�����v �E�% h ��c�?h<@�6�&����$KSw��m=�5}1�)���`�x���D�XBO�uR�����=���z�A���.�j�"8׵r��>����8�_%����7�1���Q����N�{Q��È�/�\1�*�L�J_+����"(*� }�+�����`j�п��)���t�j��gY,�7G7ޥ��[�<�jX-Q���ږ��ES� ���R܄K�f�����c���#I� "NAlm�$[!���.�F��?I|)�A��r���5CT0���*�F#vw���4Lщ:)�n�$~ӎr*��؁�)�׎v�����?�K>�Zצ�#sіz�~���`a 1���3��1OD'����V�U����ځ�M�e�;ϨcTN�#F9JS����Bt��<.��[q]�a��A�iK�����ʛ�����t�Ю#�s��Y�t���t��-�[b��Q�m�̍_��2%��~P��3Wa�zFߑb���*�nk{���e��+�-��G�0�^���][��Ŷm�����B��Q<��rP�nފ�$���=��>Yc|�fD��ƹao��+��oi�����r�	��J�	W�t�2�]Ŵ����:���<��-9��ȋ-s�% �]B[C_8f4�H5V�P�y�L���.�>�FI/�ܵ�\��F֞>�S�7L�xp�-�����͗��ӂ�8��vJv�CY!&2a�����c�9`OԼt�;��E��D]isWa��i@�::�e	���%5P]�j�X<h�|�BqrD�JA���m�+'��ICot����A:{}�m3����� ���!�{Y�\m��Q�'	ͬ���\�T����)Re�Z��9 �/��e���F�e�9!�q��W��D���w~5�Z��:A="�^���*K V�do��A�rnD�L����ʤ����������.�S$�(i�������gZ���c>�겼Q*�)�F�>���d,���G��*ʂ���1�&�Ȣ��9��,!�v��b�{�c�)��A�l�:ά�65b_�w)�+�L�ܣ��A�m}&~9�s�Aá��5�(tc��c�%��k�N��JL/Q�S˦epp�"��J]����\?�N���
Vw���ד�An;m�r���rJg�p�a�Y�nz3�K���p-R����X�N�U�Z�a�W1��l�uD�w���l�R�k�C@ZRPF�b�!n��m�A��D�s��o�b��c����rŜˎ��U��3�/N�-��?�er�m��[��W�%�1/Hn��acS� J�����03��2����}uk2��"�o��19ل��	��29n^��z*[#�F7e��O�i@_�%�������{��j |onaxh�Vǉ/�@Ȯ����_tD������=K������
(q7��<\�%vĠ~�T)j$�{���]�j�2CQ�1��M����R��"�'�i5J; 4{���¦`'A`�a�/�K�����Ԅ�^�9ŶR9I�B�CHB'u����OB�b�-=��T ����[
��W�m½����~�t]ҵ㵦�G?�J�D%]]�f��=����0gT����"�������߀�4W�i#ߺ�q�!��3���c.Y/u����^vP1l<��~'�����@���ȣ��*"���&.i���޻O���?���s��ƿT���$7򀝨����_�>��`*<Lmδ�h�Lx���f���Cjg�g�3��ȫ�8Lɳ�T�:��h7sğ����ρ��sY��F��N�pI��xa��l�Ǝ�I-�T2�o�,"K�������i���r |���f�(~.2z��=�7�Ccn��IVi&�:��ܱG���$�L��*r��^U9+$��4C���0��u��6n+� x'�C���Yۂ��%�� ?>�܋��b�+8{�hz&7Z�H�+m(��D�����{s'Pxpt�3� 9�WW�V�AӀ��n��{�y|Ǧ��=ND���Q�
�/%�gi&��Š�Bx����W�`���&�l��q�Q+x�R���.��.m��< ���µONI���$978Ғ8��S���w�i!Ɩ�*!���2�ٕ(�{VT#���CL)K&�|5�r�Ѫ 3�x �1*�ՔWq�I;�PWo���8u�P���(0�E��?*��zq1�$d�.����9�*�P.O�<�2����=�
I&��!N�p֜�v7�	���>={�v�����,mE� �/�k���~�u�EAR՘BӈÜ2�d�A ̢<�6i��B�ŵM&�Z)�;ɏ��o���t����<�e��'+����w0E��A'%*����J����ʠ]�2��b�߫���[wc���y�!�
���i���9�l<vwv�fL���Ԋ��ZډC/7��5Κ��}Dk0��G���}~0+x�J!��r�rc�g�z7zR:fb���xDd��<$ʛobbc�V��U������ݚQ�|�RtH����8Q���RSa3�[�"/ո(��8�X���'ɭ}�C�a�FϗU�Pp�F�Ĩ��+O����@\$��V<�7��w'�=d�u��y����ns�^����՗�
��q��V 0%TzC�U�t�1��_F��'b��E6�E����jB��9�ې$j4]ؗ�n�`v~��������V������	��.(ȧ
�\�(z6���]e�� �M�X^q��fr�����Ν��m�5:�����x�/u|�,.tL�M.D����J@���Hme�K��ju��'�����ʳ��4���Q��+�ف���*D�'q a�� O6Ù���#����b:�&��av)EQ�l�S�/�Z�� Q���0�(��Ke2�t8i���>��솦~�Ѥm�e��
)��VoH�al-
;���%�3j�Y�g�/�⼵���-���F��(��$�=dIW�<��e�ٿZΊ����O_��H���p�,��V��i���1[�mo�f���#qR����`_����DS8�э���z���`��`֋Gj]%H�p�`	�:VU��(MM�Z�w��������e�g�j��)���2��닥�Ogm�ڮ���{���򦳸U8�bF�n@�	�G0��!�p޷�7��^QY���1̮�A��t�����g�ǥ�TC9������圥x�$gR,jM}���4���g��!*p�H3�̈�Bu3^��h�E�u��6�#etuQ��Kٗ~�:�q��rN閹
��q�k�TL�;n���l�>�Ν@�ނ��L|��t�'�w�~7����ǏE��������)p�Ƣ�������ƾ��嬗�vr�\
�5I=��������*"C:B�:	���?�Ԉ�PfW����H�3�T�k�ND��E�p 8H�� 9�vo:hfi�2�_�m@#��綰9��"�&[~-臎I��ʐ���HL��>��0Aސ�_��q���q�����Ls��x�Ԛ�����S8�h�P�쓊�k���vLF��8����Q�5�-ㅖ����f4M}m�/=s��*�W�u��K��9F�E�r��\�Q�0���F�4�:��S�u�:xv`ZgŢ���0�Oe��5d Q@*�T~?A��� xb�>Y5�/�>.�ݴIt]�充��o�~���#��b�u����n"�w�F&��i��~+�#�}��ƅ���R������t4�B��+�Wef};�˓G�6�&��؝t���xQ��)�F���#N�S-�鰹�O5��e��a�(=�:U=�r.h�ϟ�fnu�!,����oa[`g�@��\��M=�e{[DÙ�����%I� ��jJu�a�ڢ�g�$�
��NZ�i�����|��O��fu����|�)�]B��Es�g�R�A��G\��H^RW�`a�7п�u�L
�d����G
-��6!/P����s�tLK�+nZZ�T��&�1�`QJ�6%)��	�S��h�%�_�}���di���y1(��-��9��
-��}�:� ��ݡ�9�!�f>�R�Enm�i`��%,�(�4oKyź��3�|���j�����w:�����Z&�80���Z�n�4�l%�[]�WZ?���H���H2<V0����8��h�m�'Wk�Rb�b���-Z�h)��;E2%��Ucj�{������̞F���S<��2�%QÆ�2���M٥����7Qݍw՛��-r@'\S��� -'�i�R����:��ɐ��^{���Y�k)U�<�1�R_�d�>�,�f���q��Ki�(�������[>��9U�?^Ͱꫭ۪��=��V���?��y�sJ-4�ȷl�%�Jg��)Zƻ��V���d2�f����A՗5S )6@�L�r�3��>�~��q1c܇Σ����qq����I�S��CV�[�1��/��䆚�7�t�R�z��zi3�i��2gEӍ���&�]���k����	�p�s����:%i�H^?�Q�w�*e=����T�'/���u���G�bS<"b,eӗ��W���o������ҾtU�5�ļ�w�wY�`�I�F��,O�����}5�M�d��1�4w\�5S'2.�k%1�E�5b�����Ttй���XD�\Y����&Ï����@\��f��J3���1ykωE9��:Q�pt�,��GMe�kmbU���=����(�U������Ζ�3��O�]��vo{�x%�0L%s������S�a���^{η���Ծ�mz��:J�}��e�Z���Y�g��]�(�ǿP���" ��-'0^��ј���n9E��x�@�x>�MEH�Z�r�Y�OτΣ�����:g�-@t���L�e�R��	�7rhT��� >�%��$g�9�����u(�!��d�{+�eK�aLhQ�Z`�m(.^�/���0P����
`�6�;�w6SA�b-~�<�yXچ��%�kaKn������K���UE4^�4���Ru����\_q���<�,a,�b
d�w������N�y��5�#��P��i{����K����#ڏOFMǙ��J�3Ahϳw��qp4�p�jI@��"����R��7�n`x�e7�Wqν�����A�@��=X�L�gf�x��$t�g�_����Ov�j69�芡����Fn]޼Tg��Q� � �*Ԧ�Ee	I=|�?t�_mG�������Ћ��4_��ƉH�lDc��P�AX�8��x�'��kI�S���E�yD+�jxf��TsT+ y���}�g���7H��*9�jZ�2�^�p�q�����kn�5aʈх2�U5�B���($T�D���Y�9�VHmI�GF�@�SC��i�"�c���MY2�)�-:t;b�46YEQK�K�V�#�����t%�����N��+�|��T�>�K�s��*��Z��b�X�k�K�&�Ɵ�����b��x�H��{6J�u��򒇱��?;�;�(��ɋRgo ����=Jp�c��%v�k�Z�G�������|�B@Q�r,g�TF�q;t�����1� �b�:����l4}F��-��-w�������]m���w���$�T��	�m����d�=���Hy��'/�f���=�iذm�	�'9Vuw� Bn<�)��k?�P�#���.��S����o�x<@_�(lF� �*���[�^��͕�����_�T\�i�-�A��9��t��k�9�$a.�0x#�(.,��P�v(���}̂�7�iR*��B[��F���w��R�������K��V������謼r/�yI4���C�.�r�"��f�u'���Zh�Rj�n��j�� ��箉V>�E��6{caD��w���`�u)��ڪ��c�*6ha�KqƤ�ޝ��A���:-��?����2�1��H�sX{�0 Ye�eAZNh�I� ��~f3{�Ehs�4���EL��/�c*�׼ܕ��#ԅp-��"#��aMc's���4'$��Q����2�-9?0Y$�6��qWld�n��Ԅ�Z%���~ehǈ�ZnS�{�|w쮇	�li��[��ΚW�8�mP��p�r���6��Al�������R�h�q%1�7\�!��zd�x��d�*�>�:��t�>Ѻ䱹�B=@���\4o�)���]�G�T���-����7��_[��.q��4�)�,���B#��=�J��2���f���xG�*T^��+��<�?B3�SϕBȕ�A��Q�=aB�� ����U���6f�dr+��4�Jz?�BĚ��TT��h2�\��|�.F�����a
-�	�+��b�n��[��!��4Shf*X�~ވ ���x!�NAgc\~���P)��y�e'[�{b+R�ijx�,�{t����������d��^C���R\#E�z�C2���*���_��:3��/=��E��0j�.�m9j�E?;��ƹ��o��:�L:�1��Zm+)��D�AH"��T�{l?Vm���|LR�"�d�+�}��K�_Ṱ�� �3�ۦ$u8" /�|�)7�"�/H���ҭ��0��ic��p�C]P�\�h]��
ͱ/��$ޙ-��IA�)�)^��8W���E�]>]���M��q��%PN0<�9{[���k0��|�+�����3�|IE�0���;���v�&]�ׂ0�ң݆�\ieV |�["[]�	cqp:���F�$!�}�����i!ƈ4R0Pf����N�/�V�YXyEY�>�i��>W�G1?� Q�,%&nI��	<o���S����۝�\�T�����@$$�_{AV8;dDleU�D�ŝ���m��\�U���q�7N�b�|��0�U���巪��&�0�暌-�wx�_��14��UA�CfTA�F�_�
��!��R��4���1�{��t�� ������1��e:�� v����������n�[�Y�&�~���KeRS�q��B�`�2,,��4�y��D�W�J�R�#�5j�wDx���>-����l�Ҧ����Wʖ*�ӫj��킳���r���_�/�rnl;O�̭<�h�_��M�\���)�v��.@53�KN$�����Q���&6,�+2�͌�E{�d0V���k�1f���nʰ˱�KNz��Ѕ8�'8o��βF��m5؟~4�W�<>��Gb���B�h�gf"�rܜ���rA[���9D�i�'޺�(LE�Y�P�s��z�9�O�9/C�K�|"�GrE��������-*~�22��Վ�ڄ�v����T`1��8O񶢙�ҟz��X�n��a��j�h��M���÷���C�!����O}�OMf?U��� @�ax�c�I�i��)s�ܩ�y���������Ǽ�j�B981"�
����FpH�Q�nz���_]���|-����p���@Δf�=܃�	���e�qe�hA̷ExS�g<?<�֋xGj9$�5��B1�-k;_�H�#�J��mpꝦC��;��ӹ��g`���|2���9�9e�/9:��*6��c�OFD���Z�|����K��	�}ۇ��!�Z�m��R^2�k3����Cd2ų��$����f������P��XZʞ�Ԣ�����2a>�����P���TÉ�]�:8 �I������5�|d��@��5S�p�(��rn�4�!��Zi�Edcع���y��ī�����s�z[+qܒ�������G�CM��b�w��7��!�F��W�l��BٸI�޳9�)vB����qV�j��uڛ�wY-�:���թ�����b|u\Qx�&��y��ժ����>�N-^�4�|���C�(����s����.*�͏|��޼�z�_��e7՞so�0x�Q��T��$u�X���F��km�r��25&'�N'��e����>�udQG ��������~�-h��� T����
�
�D��J%5�Ň͓���M�m�� 5���u���t�a�k�z�Ӭ:�0d���~ӫ�Fa�ӽN)�:�\n�Tm0k� શ]��G�����W�C�[&ZѨ��	,�J��	!��sCɉo9�<�<�i:����^��)�(��H{���8@���[N�>L�̕�&� �]kq8����%�E1N��&������0pBC��Hv�R_�, �*`p `﨡A�N��{���O��%��˽��O����F����JD�q{K�q(K�k��)�r�L�_�c�Hb��4�i�z�C����b���ql�1����Tqg3��0��1B�B�c�T�$���Y����k$Or����^87Y,��A¤����'D���4iih�X�#�]5��Q��7I�8o�������X�cH,`�J^9�9���5���V&Ը�� n����t�4V<~����_���oE:::.O���D-�;'Re��Y� ƼUN���tr��ic��*]��/�o�!{̣��׋0X���I�Q�k����M�S�ܬy&�BYV�f�%(�פ�,_".Y��պ{M��S����ғ-�I�8��a�^��:�w��想<��#J�0�t�����u�|�������ɑ�0�JR�'�^�-3ޖ�קD��< <&}��L
�n
��w����=�@�%�'�ϧ^����@�Ѹ���l�|���5J{u�P*@o�ی���^�jq
�[�l��V�Hk��I�uN�Vx��FE:W��Dӑ�����>�/�*b5���U,�ӂCA��%�H
�a�0�����=M~EƧ:�� 08�� ��ֈX���4ȣ-��5�7�w�Ʀd��6�q��$����\���
[dr�=��K�*oe���4aw㜄����J�$�Z)ܰ^�H��|Ʉ�(�n7}c�%�Ec��C����ƴ�.ڡ%�&��'W���"˩	.H�p
�HF�1X�X���O�y��#q�X\�_�d�|�1hT���`><ZsX�Cm�$�/���wt��q��u���v��S`(��p]�ur�F�I[��:�����.�]va�e�91,�&�x`���4Mi�Zj�Zf7�k�K���~C9�$h��CP�y�;ߟ��ɉ�d�C�*�|���q�3\;�B��{5&�%������
9/6h����q��c�9�_�`9��]�Ez\qܝ�t���o��Ҵ��)>�b�]3�������goE�t�R�B�01����)ogc���A	s=*>x£<�D�<?��l��F�����~��5S�C���`z�+$�@���Ʀ�@�jO�ڭ'���4�ɢk�I���0��7�D ���z$�$1C=*L��cF����\TU�jL�MО{&MN�ȸW�L�f�&�,��#�^pCK�����M|eۢ��f��$�m���>�v��рV�c�ք��YI��^S����j���kЦs�E-��'j�F�nP�����mY��ֵ#͘�{�nN���䏹
d��^��;,��X�����(���nKP�16����s<��$�n{���$gQk�Ю�n{�<s�|x$ޓK�,������?��p��o]�u��yOZ ��X�F	CS=��G���
d�5>`^�L�ￔ�þ�г��Es��{�O?�V���|ݑ��הο��ؙ�ft�)@��u#\�Azך�B-\ߔ1����s��":;�-�� W�Y�t�Fu��s��n�3`5�oX�p�9d�)��$�}D�ʸ�f�Q���N�	7��EC(��4�f/�F!D���x��X�?��5γf��H~ޙ�F'�A�f����\�J��Y\Y���tl6-OH��dg��K�Bs)���[�������G�\��XCDtp ��K��8�kB�{��c�3�f6d���ښ�����͵�Ux��[RCPPQ�M0����,�Z	�H��`�Q���p�wSңv���tl����7ҩ�p�������g���-�����r��qe�4��HtJC��v<sr3A{�Ih����J�x�IΑ�T��ƕE��٬�4��@�;8��C,��[qU 5?���]�{Zh�q�d�s�H��&���v����eJ�.��8�j]u�B����&�,�י3����(�Eޡm%��W�Ly7�eq�(��ܧ�c2��c'�h)�N��.Z���� q~燲v�0�g�}"e���D���Åa��~�At��Q��z���Q�FE�ym����J�&NK+Fh��z2��a���别o'�X�Y��%_Do=�\�����@���b���ͣЊ�C��G�̥``&��V��R9��L��
Y�I&�P���%an��Sr�KGkB��NP��ջzh��c�p`Ki�Lk�Z7�ޣzg|z~���ô��8���;�\ƟF��W�)I ��K�Ⰴ)n��Ѡp�#mB����+>�C�(�}8�&����6ǌ��Q��/8Ѿ،��`n`�Ew]�ܕj8�������(�r�B�Zg���qT02��J����������8������\er-�_�^g��>�i'�l_�x��-�Q00f�Ŏ)9��9`��wv$�9ؘb��>/y�o,�_�+�O���܈k�vJ������\	E�f=m��Y~'� �TY�O��\����
�ƸvPä�4��`�^C`s��Q7�tȆ�rBwo*`Րڱ�-�{X�;5h�F�/@��Oq��`��3TU�2Xz�E=G,�$�C�+v�PWL&���;*ÿS$�����R��榋c��t$Qϟ�@p�g�dŁi�d���Udf>�� ����=�%�o�j���I{1(�W���~������[��HD�&�I���`U)�Ӛ;AϸÈ��n��oL�4��2���w�Ķ�%읂��K��|��*�D4�1�1+Y��P	n޷^��h���MpK!�9���[0h��aV����÷��:Z0�b"�p��z4�l%�	��ؽ�[|�'T����;�R���ǆ���xJ�8�g�}��fl�	���l�@��,x���0W�?�!HQ� j12�Q�|�0U|FtSM��X�Mh��'�V�4����U�Ƶ4��3�m#z2?�cY�P��k+%��0�Y���w�j!��Y���ZG�����.�h�M�x~���+���3N�K�ޚ���S�4MC%b�"h��ƭQCM	!?b(���g�e9$L63�O�o��k"ў	<���'T��V�<��<���JN;S49��"��#����ѹK�\� �c���
p��UuJk'�i�sO���v�C=��V%,�hE6Yj뜞Y:��	5Ζ��)����	�,NK�����D��}�w��o�B��9QOG�P.�p#*!��)��{�_3�0*���S���Q���/~v[<�!u1`'�����|���S�F!�mz �4�l���b��N\x�)��kl�T����n��pT>�qtyq�8>�N�C���e~�R�lzkH�r���l��.K����{_5���I�0R���K�h�$��e��h��%�7�1��!
�ui�s1*l�!�7���:�\��������w���H���w�m�u����R��:7&_8��e��ј��J
�iX�m��Ȣ��0��6\f\i��7��m�R��E�$P�."�o-�i���<әZĵ1iI�2%�����wVJkb�$�ɱ�����t�>��%V����rD\Ѝ�Nɾn"��l�V^W �Z��1񜇇���+C)�)3]֠	w7S�&P1�uA2�y9=/(�ՙ��N��[I)�U�&'o��]-x�\��f�<�y|_�,3	�(���u�d"�b�2�����sĈ qWk)�O��ڏ��xj[��f��.�v�7�py$\���G�����#�C=�/��1���&���2��lS ���fA�<�7쯘���D���%u�1�ω����Z�ʔZ��,��#�W���B�ӢH��RCT��,C�7������Q7��O����
�����M]t�2OwŁSV�FN�&� ��.X//�jm��Dy[{|�b��M���^}템�Z��>�B�u��A�����"����DP!��T�ɪ��Zm�F�@�x�CR�R���-V������!�#��g�� �z�9R�6����}�\���l�(^�H��=���E#ޥ���|�.w5�Lp�H6�NH�ǟ&5�ͣMj��Ŀ�+|�;�_#w�W(.��ˢ�ƈ���&Ie43�� ��R��LW��[ɭ����G
�ƍ1��G:.ksT���R�q��ո�|�0}97���a>��'7��=z,��\V&���I�$��
w���=���vF��%%� N���b���}㺓 �غo�}��R`n?]�Az�I��ϿCy�
N&��eo�K��Y��䠒�6���zv�JM��a��GI!�,k�crqz!���&�����C�e/���N"yY_���)e���)Ư��R�� n`��kJ,v SY��I?���tU.C>���ze<����l�
�&���U�/s�S�Mj�����Ϭ�l���ɧCb�`�#է��ʂ�W��LkQ�%,�4��H�����s�Z��iIJf��@k��"%BW�瑯��S�X�D2��{�\j0s�&D��LUQ��o1:�.7vc�y�]
m�`��m�y��l��^��"��i�WC���57�Be����,��g\�}��te>�Ѽ�9�$S�P��a۲����F�����S�x�?�nX�7�2լI�����s7'; }"��,@a�����i���lj88W��'�,ȋ>'l��� �n��{��;��5Aiz��]�Vt�>2�4��a�Wn,ri^?qO[����f����ث����d��nu8�КS3����{6j�uv�Q��1�r���X5�;)��`�23D����Vi��2]O)�G@��� �pWZ� "9."Z8�(<�ڸF|���n���l$��g��Lo�#�ɖI�~4�f�x��fzr�pΡ���jf��k ��O_cd�Ƙ�I:jA�8�[`�����όMhb	`='��C���Ր�����ڨ��mj|��g� <�
���D�U �ɒ���8����Ҙ2� �t�\2��`�Θ������W�=d��y���8�;���v�T;;�H�^�����
���&����(P�==_��H�#��a����f��6��\V[�Glm�)�+�ޏ��PHHC&���q����D���o��[a�v�`�uM�����՜C]J� �C��t
C@eW��5'uV�jcU�7�kH�y4�х"�ܓ�����k��"&�PQǒ�u�~�z�6��`-���tQ��!�-Qp ��'UKEPz�*��U����@W�q�����M=.P���!����E�̹�pZ����<�Α;M����6���<F�:%#���j�Σ.%��\�Vиg�U�{�
��>m�I�����pw�r� ڤ�ުd�L>��i0�4Oa��Uɴ�/D��1�^g�<�^c����&�0)�Q[ً)�s�q���Fz�e̦���1^r�������5K�K֮o�L�*Dnmׄ� ;�+ǜ�	� �)��]&��rL��-��hLOb��[ynŉ�e�F�!xWm$���ә	?�=�]D�}�?��焷���(�����% adO�c�!0��b���
Ts̬ρoT[�OT�<�_�����B�lr�|��}�׺�I�Ya*e�_�>���uF�w&����:5������p���5�L���w�ޯ}�6�<ҴZ����Cz��_W
J[�C�ڳE�d��ߨ3/�֜⬒�"5��N
<�]���(���Ҕd(㣋�L�6�&�8pW��B�N(~"U��}�fM�蠀/�F�S,
��V����^T����`Q�79i��~�v�
or��`�����ӫo�x��h5�2�"_�\������Cz{RK?M�94�A�"6�+��!�w.Iɾ�+�7����ɹlM�)l�L_�D3��A�̽����k=0�R��b���Pf��8���OedB"9b0�	|����`M8$�!�LYB���ˇ	F��E旑N���9T ���s���<��p�`�\C��O�R0��j�x�z�㋒	0&-OG9���N�O���ί�<�p���8��/SO��a���$������{��Y�&�6V��~f�S0�������D�Y&�`���E@!�2
 /��b�V��[���?b��i���YT��\}�(��F��
6��Z�p�������H.M�$�38n�	�y�r�M�g�{��3����E�"���,��㴥�>>��S�����]����Êyn;*r�aDC�pɳp�b.�p/Z�q��>�A�xM�i1)�t����$x��;��-_ѯ����`Kt2Q�dp=Ր��u��0ĈV.��*�~�G��S38�^�#��w)쎅+�$�ae.ϢbQ����s|OG�� H�-$&2���H��,�E���� ��<�f\��{�A<��$g�o�(����zો]~n6s7W3�L�8jF�y���!a�	�e��B�KH�G��<��$!�(m�9��i6{��~�ļI�i���(��5����Em��/��e����Ȩ����˔
�E��ݹ{� �F�D,�c���w@9A�ji�/��*A�9T3��L�Q�:;����mύ#o��0Ml�,�)�w�L�M��ǖ�+b�J^Z�<����l��S��x̺�C|My���N�"��;�IcL��V|}D�YK���W3���<C��4�\���$�>���O�P�ٿR2�Z"1���BT�@|�=&��Ǐ�Tz,����m��0U��D���\wg���g��O!0xЊ6�-5UF�D�
�_Fյ���G�KgƄ8v��`��lg��YM��)z�N��*�ߋӊ6����eG�h�J0-��I�\�x:ra�I!�����	,��e�}�{�i���0�����dP��M��栉�y�4q
�:�e�V@ػ7�
Ե$���4`rf��(Dݐ�Z.�zW�{��t�vDB��N��C�N�p���͌H�G��j�S�d��߸0�U��W�|�\�קz�~����J.k�j)��<�VH�\�����f��o����,j�Z�AH����ᷞR�����*1����b1�5;��%پ�0j5��<rB�KԴ/T���u+@��P!��6�}q�n����iw�_Z]j�Q{r���*���%�(�)�I��:��#%%Y[9����'��Oe�+P�x����x.�j)vbG-!1��f���K���}bׁ#@xf,�?����Afz]�3*�A��}��Z���F�ϫyX� Ȼ8E�ɋ4�S$��m�g}���"�p��!�yb���&�&SiV��V&�9�w��L��B��"��uəR�b���gF�se�?�������$1��3���}�_�evi���tyH�P���\]�^>��oM�6g�U��m{�%�sq�n�I?���q�7[��eX����2-�z
�dY��-��)�\�m��
�i�O�m���n�-Wؕ0A}��%��SJ4�u/X4��7?��Ĳ��k�R(95�:���v/��v-zIt���fva'�� �R�M):�,�:�Մ�)�
{�<���%�������������~��:������5� �!�_yv(./l�i��_���o���Z=�jg;n'��� �G�
j��Htn�.�q�U�f�68X�*���M*�JWWwm�����P���uf����-��8݌}��0mR�M!DF�]�B�X|��0�|�
����"
�jH��݆��QY�iЬ[l�VG�.��0g,I�}���S��p=����76:���_�%����~EDYA&N�S�>�,5N�!Ls\�w�
�y�;��Ŏ�^wv�{y�n)���i�F"��6Ո�Ǔ[H4Ur��>��V���j�j�C<�G���U.v�������Ao��Ƽ0��Qda���^��L��򱡽��Q����,mT��i)�&�SL��LI�'�IL�b����t�43H4�(z�$�[�����N�L���Y��
y�K۷@��(��-�a�\dk�H:��uY°�-d��,Yؠ�=J�$0�@TfI6� ��c,{䣟��P�𒌕p����N��
�U����S���6lEQ�V@��U<�������X�R�e�sA���ӏ�M���]SQ���G9yd�,������n�����VK3�a��p��+�X�8��J��>()��&�>`ڪ���-�a]�u5Or���S��SzH�2ѓ�5����6C��Χ��	;�n�MvI�V��ܧ%;�����w�,BLD-ĬG����ɑ��O��Hq��pt.������:�}?/�I�D5<oJ�I&��7����$�"�q�zz_7юp ��^?FyTq&��*�NX�Y"?vڝ;#�@H��9U�s���ڮf꼓W��+e��M&���L��g���$���J����Jbj�p����	�l��9h (cW[� .wJ�n��v��x��Q�;�zf���yۇ$�b�3}�-����b��FZ��XD�&Kw[ó.
����� z�K��i3
ʱ���!�b��W	����Ev�2���~��0�f�%m-��%	,A��X�չ��&����G=�U�l�PX���K�='������a���^ٚ|�pv��r�rQ��.��k|N��]� V$�.�ΩWj�L׳�f���_>�.��m:AN����-/$	}��p�XhF5����7���֑����7��@�%e�]����VP@^���>PH�Q�.B����&:��Ve�h��r�j���dO���w��Y74���+�B�r5G�|ث_�����F�G�2^�6����n*N� �XM,�rY�#s��z�u��Ն��Z����臏੩�����$�s��X>͐S�z�A�*����pa��?�i��2L������*۷Y�߁&��`0/�p���[��I�u5�{�hh_���v�p w)��9"Ē���+�v�F,����k`d �"�bD;,�tmx*��}���*!,Y=T�._6�)��2����Y�RB+a�ø��q�[~�-��>��G孥����.w�6hCl�}��G�V.��k�V?_��p�~���
�3�S�r�Lk>2D@]��Oo��tm�u�!�Q�Ҙ������*5��j���t6)yV�&-�����?"�27�ӯg�3,���B*�z�`ĺ��Cp���%��@`t���l7��%笾/���3�����Ec[)9�^��+ Tە�Ġ�w�� �1d4�:`�8�
RX�J;�Y?hU��C� �om�*�.� �Ȭ�b��e{w�*���!ֲL�5(�y��=�J��HɩDLަ��D��l�8�v��6a�B�K�A�C"��^[���F�<�x#<��������Zq����N�A�I��<��P?�AT��*�-��nFDNaAM͉��W�A�&��;q��#�q�<9`>��l�S��p��4$�������.v��,�[�Ϣh��g٣�py�h�@��5�mK�������.;.�*�WR���a6�P?�fO=>X��hN�1�� ג�Q���P��sW8��1� �PO�.�x� UTF��O��tc�}�z�r��jM��%���d��7L���L�d��?a��F���'s��M�ydbVz,
�����v7�Jl���QGF�]WxR�h���N��"�x?�l�;}��~$�[��ۢ;N<����&1cR�>PG�r��,�	�4�]"ä�;�5�	Ce��	��ݹ���S�*E8d��ꐆba��4gQI���2����l��ax���[���/�:3�t�yն����3�A�Ωm�GP[�����	k��_�B͠��u�rw s}���TA)7��_R��V�F=��lD���~-����B8�(��ҏ�Ή�v&QN�j���T�S&M�l�	���/4<9@�D��%�*(�tO��G��9��!�h�K̮ʞi��EŲx���\�̱Ü���)m�[�z�C�GB�p�-�H�V3$�ç��NR�T����^@�H�[}64� <�g5Y�����i���oS�}~�R�Ĉ��vrJ��O�N�<�:�>���-.�e�UD��W
��d�2��L�\_߆��[��BsHZ4��XM�s���j�m	����, �2H�����X;�Å3ɋ�J�o$v�Ȗ�3�X��V��|�uq�{}�:�nߘ�|
�q�_Te;i2�sǿ�߼�1_��N��N5d�5���iI� y|�-�S��ޜ�6� <69�i:R��� �Hؗp�1AT��c�M���a6;.t���P���*��+�/�iJMbN%�[�l6&���j��S	�8Q���jh�N��S��Wr/�]�|��JMSM9�|ҫ5ۺK��m���M�+&{��ja�D�W�a��a�ǎ.����9t(��]b��d}�qo=�k^][��m�eB��6��	d-��Vy%����kg�:]��bǁYo�v�yG���H�ek�>/oڼl��rx�y��< �:�6E�������s;0䛛����`���/j&���]�7綋�E^c�D�h�������oQ�A�?���2�G���+d+A�8I^/x���k%�Ɨ��T�H��7D��<��C���7�(!+x�ml"b��t�HB�Z�Z8ͥ���f�lm���ѱ�E��yH��(��T)�9���S��Z�c8`�T�-����RP�Y�"P�9�b�|�e�t�F��7�*��Z��Q��+�Kg��%�ǉ��'�O�J�7@�јj��2[�B J{~�PU+�"��zݬ�'��5�.§{��PE�U�O4�un�X�j�&m���>r�1+��_��9D��Tr��W�눵��Jև�3��o�W����7OҔ�T6B"뼔�=���-t��BR�_���������hߎ�a�e?�%T�F���?Pp7�'Y�GYѧ!�3[�0x�Io�����.��@�ţ��&���b�|mt�YkAU�V����!)��16*��t��.�R{[�f�2.*��( �k�X�#l�^Q�#����X�.��ڰ~Jk*���{�Q=�D�eyR����}��<�nb{�����-l`E���8sEE	����P�ǡ�'83��'!p9��Jk����V��Uf��>L���i!�+Z���ce�8+������D=w�y31��=�ê� �
t%�eU��2	��=m�>�.�N�(��f4�.�x��[_�s�Q���M�<%n��uD�`��\=qnKD9�W?���TA���4<v��&�S�gޜ_� �U��9��y�^2ږ��y�H��o���d�^{�.�֔��!�f��	�x�\��l�����R�\����B���A�.� BG�����o�j���P�6���`M�L'd�?tml�� 5�kJ�Xnf�A*x)�Z�=@�W;�Fu�U/�W��H�{<�Q{�����D�Q	�V!�|8�N�ܕ����=�2j�ן�Sœh.E��jPz�m���"@����%��U>y��q�*����a��"��c���v�GO]@�x.V�X=�
�`B�I{	�ܘ�$��@_*e�\�����+�+��v;����k�g��iU&'n������
����MU�wNc�4���q���ǇP
�1�f*� �����?��(Nd�+�!��VH��|�o�߼�A��u|d�[�4S�[�V��z��;q˿N�3�DG����u���'P(���t�p��ŔbH�j�h���t�6� }�t�#�	����E9r��'C�����<?3m�fP����D�x N�z�龝q��5�]S������v7R���K>�B��|-O'�Tsڪ���=$�7"�����t��X)NG�댻���Z��Tn�5( �>�{'��E��w�z �b#�����)���`�mt�_��^�|{<]�8��{�����ƦҼ�@���aU�m����sp�R�X����N���j�c_���a<>7h�מ�7������X���?@}t��@����N�$/"�K�d�_9�5_��=B�N�U&���Կ��IO��B�<��~�2�^bcz>�EO<K�wU7�'�4�]f�����cv��+�n&��y��|��������ޙ-4[�Tl��6#�;��2�ZH��/}a-�W$(�)U辵f'��E���� ��4�G����2��c=CdyH�8ѱ���	�-c�`�#�i�97W4�9��%���S�t V�(��]Z+��K���P�ޏ�(��� x��j��Z��5���f-�����z=
�
-�RqaKuY9hQ���m
Hcʰ���vV�#q�R"kP}@�w�Y��<���Z���^j��k(Q�"@��n_W��6p͆�r���AΉl���"_�ˉv&O�4�7�����4Q�p����@���0���s�͚��ӮI�F����7x ?R���Jm���"��$?���z�BBm'�j��[�^��p~.�%��m�&�Q��J��;��I���*�xd'�g��QC��bҜ$���ZoE��e�V�Y�'" 
��B�y) Z�y\�*�r�d@Jv@d����/�vG�HBh�fe�*��X��޴<7W���DrY�?��y���ˮ#=�"`̷���I�ӝ�l���UډxGԧx�S=ҥ���U4Uj��k(�5��2R���JӨ���o�����
�V��Ѵ8� ��^�x�_�3w���k��o�U�"�~�\�7��"�0��W���ʶ��)<�[�#��G��J��X�H#�f��jl���@x�O9v�e�a�q��1�C5u�X�ml�Y�/2�Q�}�ٙ��&C\U�����w�}�E��PG\�Lx4����z_�y�J����[�G	ڪ�uC%ä8���=�im>���*@�) ��$$��n�t���/���9��3�K�9'g�I����<������n��rY�8�`p
w��Nk�wƮ��ݷ��aإ��p��V��ö:�V8������� qS��¥E�\���(Y���H��]h���&��K���bߍ�7Eُ�&��$T�ǳ�0`���ǘB���	<T,����A9�uE%4��``J���݉�32�q��Fs#���"�3�-a��{b��~�����v���V1�l3*,��yѱ}�&:WhF|Q��Ҁ�ݨG��:��Wq�ճ�^�I'�x�f�efq�#��H��I�ol�A����`���'�����yA����
�[I=BG ��^f��v�-���~K!!����G)��O
!u��<��?��Ov��7�mh�ѿ3�s��%W�~�X7��Q���#��7�zo^�G~U���Կ?{��yO�](���\��T8к\��J������!�@�b].���>�9��2bcH! RP�y)�,����NnQ&�� J��R[ Y����c�!H+�N"_+�S���|��[��y�t;����xuv_���su��8h'�@��r��G��1��s�x�na��������o��&��T&��
�3��	Ŵ��c�6�,�X43E��4Hۈ+~�eZ]���AC� �·�u����謬�*��vg杮^�E����-�PZu��e���ߝ�F�W� ^�7���@�lX��A�����)�SB�~2��>��e#T<���L��WOU�r��-��sѐ��keH� �� ��6��?I�n���f��xG�����7�@�+QRr{9rp���B�xI�qdc�D{�Y)�+�s�8�GĔ�5��J��R�S�T�7�^��2�#��u�,�F�C�T�,��%,�KqPk�vEEx�b�3=�IL:���9�4�$};��,ܔ{>�c�ؔQ}" C7M��lL X�tFIbn�A.�^s!�R�ٚ9��|%(O�cX��s�0d�xL@�(Rf�LU�O�G�GW�g��I[�.,�)'U�Y��o�{�ك�m�����\�숩*C���f�}n�E�yk�%��x�|y��X��|�If�Pi�V�U>`�+���|ʺ�v�@��:�(�p���pg5 ;��O�-t�cI��|�����;n��� ��d���/39���o'�RcV�5�FB&�.��Hj��՜k,vv�+�� �:x1T�M1˽W;�]�o���`$y�1ɒQ�w˷�ǫ��s��K\�y��eM��K�ֿ��i����e�>�m��%e塺�p�8�_���UO;L�HbW]ճF�טo�j�T�H[�k?���ř�8�ֳE;[����;�����Xtb�B����s^c�(E$n�!��t!;J+ ky�@����-e:����=�މ��o����d2����m(����Tc����7��C_^k�j����TwE��AiP�g9�a<�c;����SDf����ۑ��} KEw^��z,u͙-�y(��Eu���v#����݁b��)�����|{ �+�Am�И?����H�g�Fš'���MMv�:��6��eH��\ �b��:�1=���F�eS�K�H��:6�/��xA�՟�
I�G���6z�M�l<�Dثm�^�yJ���\xkﻕX�	��?��*P)ab/X���XIG��1�3B��Ppz�	y�U_�"&�1�؉b����>��Z`U.m����%�SϕFΤ���O���t���rQ�^�����$�h�A�2Ld��^��t�)���y3���cdQ���\��KUZn&'���� �%��
�I�'�@����]��E�R�ge�Z�E5ʏ;݃����#nT��c�r��t�PL�p�D���;��*���l�@rR�}�g<����[��{�}A��m�����#r4gokC�S=odUA�< �m�� f���r�m��/�G���"�>��Ĳ�]e�n��X�y��.��`6�7�7�x��P�ę��&���� G%a�_zy��-J�
#�D=yu��٥�iƮӗ��͵�7�$R$fh/��%U����Uc��Ē?ӭ2_��k�8.ce$Tg�D �����·X��ԒpH����aj@!��.^�8p̲k��d>�"��j��.^���'��<��ӷ��KV�Q�
�e�A
��(�E�N���^�t��%B��}�8.�/P .Ъ&U�Z�0��N�X���)�L�O��3�U%C~���`�S+�8�\2��zr���0���8v�����Z����wJ��o��F3��+֍���J�W�M{��(�T
�B�L��6!��hGf�����ʠEk-���-s����hzvØ����� H&y��4�G�$�J: ?Ŀ��GK��� 넥7BY���
��V�#,3�9��?�k�3�M^�Y�V{fp���l��S`�FYCT���^*��=',t�K���k�Z�(�����ʆ�%ҝ�M�z��S
�axv���^	Z���G@os��8PK�Ki���M�3-��!̋ˏNO�����C��HƤjd�!�w�!p���]JJk�\�=�l<�:��ᱼ�J\^�_Oy$�^�#vE��$7AY�L-ӑ�>���,0�����6-�M۴�Q��I�y��U; ���JJ�ҩ�5\A���c�L��ү �\3��AO�4�}�˿�"�ŧ�1��ՠ������,�G�'a�Gú�K.�eTm=�`�̛�U�DZ�[\�!62U����;�q0��� �#�Ɓq]�V���y��R�y'���!��n�v���qEf�w��`�j�!��d�S}O|/���'�E-}�kWT�m[?�w�8o�+�*NT�H���V��u��x���Kg���N��s1�Ew$�"�4Tg����Xjܴm�۽�5Y�d�{)���i�^��ϧ���K���&���Q�P����ql��*2�"�����=�1 �Zظ打���	n���r[,�L�����5x�����*��Y�ە���<F2d)�)�$Չ��E��Z�хn7��ׯ���>B$��=
�ln��U�F?����8���E���
,�87E|A�r�둥�hb[�k�O���P���{^�,��Ax��=5{_�M����u��Ԧ5(n��9fW{|�6����S����Ƹ�+��?�r�V�fte��Ɠ��P؇�<⪹nz��-�3H�-ɀR)�|GX�@'
��HN�v��UK���1�����������Ik�:�_��'�Q��l�o"o���� )��oe����k	)�	�lmP���(߹f�jf���p��m>��V�v�'�"�L�G�{�\�MXE��a�Z�n� ��L�#�s�H�wL4b�m̶��z������o�
��#xћ��:�{�����X����j߀��f.��������1b��^�M��F�k����\����8'�j��M���%p�M%���3��1uI�L�k��uW8�pJEE[�!������f�s��B��{��4op�Q�jbg
L�Fk����[iR�p��6
*��`���}&�BL4&��<���l��m���I)�x��f����0���?�{C�z�Anأ����v��E8&��k@&C��r�*NФN���
�t�7�����[�@�A�Z����,k�\]A����~#6�J�H�WV\�l�?�u���"���/�t`nAb/�1q@� n_s�j$���D䁐=�Ԡ�{�l�2چ}�To�>-_��j_JpA�1����qDy�?�D�������G��7d�����"?Yz%��� '��R�ONd)��.�S����|���9o�b����3�W��ʢ].��~`���1�kTd��Cx��f�^��뷍M�9�9a��3��O�0ml��zd8��[[W�Nb�WV��ѓv5DT봏�tN�0n��rh��XR��e��X�o�x/��M�S������p�v�c�"��K�j���U�M��RP���Ϸ/����j���~N҅�����z�NJcN����? #v_���`B>j��*��ݷT�۵8�:�0�	�ܶ�<��v7�Tt^G�sp~M��m��~W���r�Չ9��=ǂ��t� ��՞<9W��!�ݧ���v�CO�)%�-��ˈ�O�Ι�몴�L)h��;��-���d�P�@��G^[��P	#��.񐍁��gY�*��=\ɧC~�F�NG4���NFL�P��ƯqPB��P��&_ZW懻��q��Ks��o�I-�Z1�S�J��T��o�k�	�	 ��u�X�'j�	-Uk��Z[��8�SH���eyd1*%J="��P��fcؑdsק6]f/��t��}�q,K��a��,x.(��+Ow������Y��9�)�����T�%w����'�*��U -�������/QH+0��|h+�D�K�D�����WZs��~U����l��!*���