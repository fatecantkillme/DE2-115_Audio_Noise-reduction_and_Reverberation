��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<JÕ���<g�䑲����|J���K�/���7�����5�'�\Cm��оk������v��RGd�A�e�)�#�2���*���66GhM�/���fQڵ� �;�]I��=� �(P�[��=�T�e�6U�N�2��X��鮱���lp[z&PK�$T��
}o�����h��)w��#;e`鼅��2�^�ls�7�ݗ\�7���A"��,����Z�#ޕ w���F��s�ǫ�9q��-)��m�(��$z�}�V�Lu�W�+�S�
"�܊���#D�[J6������(�q��%x��.�1h˶�f��<Q�MQ	�x%$��ܺ���_B0�?n*�3�UB�O{B;�̸g�,x4 ����\F�E�������Z9��'��B���U��J���.l��3��s�	��Q�prmN]�J�5�`��sjpn&?K����|WW��T��f�܈�Z��lA�_���O������O�%�O�����(�@UFG�g&�4�u��B�x�*ZH�'VAҴk�aֆ��@�b��N9V'E�s�	 3�.YQ����ŵW�g��%��A`��jh���>�"�>���B���+�h��*�o�zp4�n
��(��ۃr�g'.ӥ1YC \&j�⦀���u7H��C�G
�\R)�>�ځT��FD�w~��$��}�^�62�1f��&���1���k�a�,v�k�|��c��-WB�޽E
�2(�J��$�I�-՛h���+W�ʻB{+%'p�vs�,��G�ϭB��u���m�� `tS��7���h���)5�A�e���Ǌ��e9f�l�����TME�q����~~vס�-�|�*� Q�^��.�>����T���	7eʭ��>���n�![�n��n�J�k��m�Fm{mG���dBo����C�C�%1��۵"��Z?��w.!*�Jv9��Fḩ��SӦ�d��%�Ui ���xp�Ӭlt��F�tN���C���n.\�f��2v�߿H�qtL�u���p����ZV���y��DW&���P�Ӯz����՗���q�g�>����:�T����bZ���J�>�!d�Z�u��}WC$������	}���>��g~ni�x.@�3�ܝ&zA||���e5Y-O��%�Vh��?�tO*l�Qb�Yp�[5f�t�"�F�,(�5L�z�Z�ϱ����Ir-<��}���¢����!���4�$0a[�(H�h��V��k^q��~S����c��2���ލ������ya�)�w�o��4�e�	4�N��3{xTcDi+�$� ��0��pA��2���\T���zC<J �F}W5i�8��b�4���6�5}�;i�����>P	�M/�l�x�ѤmY�D}A��E�8T��z���}�c�.#f������k"�z%u^�`�*��*��@�mDuAU������L%F�:�皷:�Kt���+��y�����LE�畑�4ҟ9A��$��
�h�5�l��v��~�m��"��lI�rZ�� ͼ'b��8���a�3�s��\��k��񅞻�����P��]|W+��:����$�r�[~�n��+�)�i^ wK[��''N�n������)��Z�ĵܽ�	��h,�U9jvf(�/9cU�ߜ�u�����<0�W
+�Dҡ50.�W����j��[>def�Nޭ���j�*^�Xc͎Yռ���i/w�6�O%�\�^&Y��.i�W��W��%���0�l�Y�q@|-��O���[���]f���
�ꜩ�� YAj�VKZ_գ��^Qpj��I��1]y�#�kpk�su>���n���?EzI�(�-k&�w��v!�����eY�Q��4��tc �3��V54�~`\yqi'��L�N@ 1wj�;:-���!AB[�H�yJ���x"�n��Y�1��vi�)���ӸՕ��A��Qi�K��o#����yZ$���NYʏ�b8:��^��Υ9�q�l�_��ڍ�&��!�J��D���ا=�55W:�}
�n��gA�1տf!ZGr�UC�ʉ�t�^t�����/-�__�<�D�|�Ĳ*\�x�L"��`�ߴ��B���iw:j������:1��44~t��N(�=
8~}\%�$�b��_�Ѩj\�QPU��u���u���]L�*�bh&°T��C���᷻.�� �;�	L�T/�-tĴ�
H��BQۊ������J/�w��U|Um㖒��M�hd-2��k��S(��"JqQ�->��2��B�r(���M�,*g�h�5�P���-�F	�֤�[[`B��Ir��_HTY
2�^��E�*���u����f���y�`@]�cM�2XDH0�\g_���U��Ȇ��-��~|HKp���p.�(���������S�D� !��狿HPN��hz��>����l�\�Ą�[�^�  V���L�
j�2J����r�n'�h��,�;39k�T�
����@mM�����p�i��ρ_�
�R����7��q��4�v��2�����zf:5+}��Fr�SdB���&���
�}듿�բ�Bx���A�4"QT|t��E�..�u�Rc"��@��#)/m�JhCU4���W]��ˤFk\�}i�ɍ��(�z>�|6����р����W�ڏ���/#�P����IOm���(%޶�-���gf~��tps��f�8��]@� ���)͌�}�Y����T柃&D�3�=c����5�W���w��إc��li�j�>��)ZɄ�`d�#LH��F�I��͈2�I1��u�xq#��ه���;���K�-�� ��b���B7���*'��ʖ����$G2���lst"�i�I�>�L��;���E�/�#*���|����;�\~(���#g��3�J��8��#5����{�}�*�J.��O�ѧ٤U1�an7��"'�S��}��vc����Χ�Q��ɟ͚~V�p4��Q�ߔ�/�n�]7��[p����ڨ �t9�;_W�{�:�-�	���L�C��g��q��;;�#��~Oi�R��Y�Z�;�'K��x��EE5{�/n�@�	�c�c�����ݱ����	�@���s�t���ջ5�#O;p�`��\wH�M���k^J�`��a�g+�:��z��yɠǋh���-Y�&0Zm�78��Y�:uq�Djcc�d�����2W���%�]�6Fu��	%Jx\���T��e����WP����Yȹ��V��)�4Kw�~)Ycc�V_��&P����@��H��r�lk�j��wOA��'�֢}�0SYXc{�<Zi�Q����N���v8P�V��E�j�o��0e(M[���H��M�cN��R�hc�:$�k��/�Dפ\�8ԧ��.��<�`o� ��sa�?�>�]#�P3���r,��kV�)o!�����̀��\���7G�#��~��,0��} q�_�Q��R��V25$A�J������]���r8�HE=����!<��-9�����b�$J�(��C7R	�����$�Yꮸe*���p��-[�1�}^�+��ˣ�(����mYJA����y�:<I���M��T��9�=3��Nrd�ަX#��t�*"čhVL�~�Y��^ð}��:龲�SLl?�����~�\p�%���;�(~�Cy����7�{�j�ˎ���������z������sK,M$��bA�/H�ސM"2�O�.8��#<��-^����/�%n���d˔l��4��w�	���;�F3���tG��޻�^������*
�h�g6�e ��I/�R�j��u��'�g�6�0�!�1�V�.��s�-rՀz�*yl�h|�D�\� ����+i,>��I9-q�����=��.Wtw%�B8�����5�sOZ|�u��� ln�d����cm8�C�����Ȍ�6�N�8*8YZWJ�fka�(=A�B���_l1�����Ki5��ȹ�4�&�*��ۈs����Li���}}dĀ7�H�2���fH�n����m��ճ�Ze1�D�����G�ŦcAf�"�����f_�;�s!�b�sw��m�kzc'�:3p��J�T�$ַYr�T�9�Z�Ǿ����J�"�&g�D���$An<�8��8���2g	f3��{̸�?����z���\�,���r
���qX��S���:�r�t��}�;��h¹�m��h1:%��$�ƱQT0;�s��a�`0A�GKs��_t͟m����>�B���bɭRb�<Nθ�Jx�#�z�0[�.�>
��v�����z�zkρ�:��4�DU{g�K��=Fv�=���#]\�F�=k�̒�������x̖H���'���8cKl\�[�s��$V<1t_�͖��뉯GI�����ٷ2���^\K����!�%3K��|�Ż�-�DJ_G�L�o��&�ߜ��I��-N�F8H��h���&��F��؜ª��Z�.��Y|�i�x~�i#���o�x�E6OJi�� l��\���S�>0v�ϳ��/؆���Y��*��ȸb����Nk�B9q��D{c�>�\2FOV��@���ɏ��y��H]=9���*%t�9I���f˞�v׬��ô��i��
���_���a �3�����v��2g��|���M�a�)�VM�	����l�o
��I{L�!�����G0Oop�/_�~Y��,�Ș�@�-���A����"���ߠ��Ӎ'��k�B[[����ͻ='mS61���fH�	��z'��b��K�Z۾l�����X$��/l�=e�3��*��Xu8���e�o�\Nj&6Yŝ�غ��.i-B�(��:��i�Z���ɏa����s �ZZ��Zo1��y�/�UMR:'2S�[���S���C��ES��R�^���2�N&���k�E隂-`��^\�]	6fI�`u�$��Bx7�P@E�{@�lw5U ڂ��B3G���Oh|�����$*������H����S���v�]���|����:"?��r���лe�r>�j4��G�?�6AC��O�JL3�B�zR~�l%�d���Ԏ�W}��t11zkx������`�{��>8Уr$���.2�ƴ�5�ʐ(��0k��Gp'�l,��J:P�����m���[^EdD�ژ���8���2�Ln$��B�&}�I�.�CZx{?�YB���0��s�$*v��P�T���I.�d� �T��M9�5{���^�X[<v*(�9΂:p��0�����)]�Ō	Z3LrG��<L�<�H>��hE��[.��>����6��r<�Q��ٔ����G�]n
ي3�����9ҁ�M.��G�f���� c��<p���X�#���G�L�G�f5�������m!��./�����SJ&X�o?�����h�T���u���s+5�F4@Y�"�ɘug1��t����Ge�φ����d��R�$h0-�*�k�����i�����Htg�{���bc�y��|Fj������E~���}Lf��Vgi�o��>�� #N�_����bx^��lܾ�/���"0'� Jn-���V���'��?w)M#?}�R�����o�P�X�ڏQ�$����O �Q����T��� � ����zU���,UNoiN��1����`�7��I*m���4�2eٝ��Ȓ&_�u�T�|OM'�W��8�9�$�z1�M�V���0�����w �$��!�s}�]�yJ�\�=�&:�{�;��B��}48����F�"��a�?or�1g���`�fK��m���'`�(�w������)�&�D��R\R0��^.]��������k5�ڤ���h'��P��\W��r�q�uw<��r�J�.���է
�ptJ+h�|����	�4�^0��r�Y��*L�z��u��Ldȼ�d�;Kb���2<4�㕠-�`��Y�lsT��m9��|���㽍�M�ޯ[[�OؖvZT��6���qN�sD���"�\Ee4p�R�dmǉ�@j��7�^�G
��b���Fކ�Zd�/H�����w��"zE��C���ѫm��gY�A��y[y��-�����5Һ��B�+]��6�L�4�y�UJ����Rf�2-'��9�S��b��ڌ[�4+Z�"�����Uc�Z��}�����+�(;U���,,�#ц[T?�
��t]@I
���O���V�c��4��hKKJ���lq��ʭ >EV1I����Nc�upUܺ�h9A}��xk���Ӳ .�k�}+u�nn#�l~��*}0u����C��e�8����Ǒ�QF�cU���/�y���~����f���6��6������}�����R�n���k $W2�߈���<�bz:V�?cÖ�>��`ojx9 �Y5���J6���jG@�,P�����N��� Tga��/ܴ���S�6-Ac�"{?m;@�%ܥHs�)��ϥ&:����\H��#m� I�0��o�h��)J.k�����Ƣ+�����lfҚ���D����"*SS�@n��U^��@tƪ"\�'{aF*x�Σ
o�o�NjH׽���PFv�� �z,Нx���-S�����Pg�I^�R[�[%/'5�y��6�*	dME���3�O�8y�Ώ��ax�]lS�f�Z����u Y��_F�-W,�)��n���C���q�Ʊdl.��k��`������-��ȏ����γ��!xU Tj\,�Ch�7��jw K�~Żh+=�J���<r����c)d��yg.1/'�ꡯ���W�*�ѽ���u}��.�ot��o�{^������*�D���H(�[O%G����*����A-7 ���A9j#+B·t�u`��ϰO/+�{��Gtk���,�2Wc�,zb/NVu�;��g��4��+���!~�N?%	��V�t�Ws�`XR�k��f�?�;V�P��6c���V�m��W/B�Y���~�+W��c3Z���)�_/Ȑ�zǺH�$7�j�[v�.�|;Gj��I��nXKb�\��}���8�LlAN�cfZC��y�L��^*0�P��ap��h�����Y��/�,�i]�\�h�#'� ���:9�:��k��k ��?|%o�Y/��0���}�L��F���Y׼֨�m[�'�z�+:R�dGgQٞ5���ԟ]�Ǯ���f���������S
ÿH�aM�.Ê
N��-��8���z~�/� �q�f*�:)o<Ϲk����p��>��C4,_aV�@�b3�i���G������r,:l����pEg�D��4����-}w��kl�re�0�vu ��r�x�Mϻ�B���i�P	s!`k��i a^���(�z�o��Y�8��k��&�U�R��������ÅW|�&2���}�e��e���`�6#1��t���q:�LR�;C���=�8k<Pn~�A�����9	���Z=�ײϓP�$�҇��H���l1)���æ���Ef���0���j�ެ~µ��������I�KBi���'���\��G�6R�2�L[��+ݥ����} ���O��02kO��t�"��b_��ӕ�������޺�`~G��Ѡ��E�;:��?BY�λ��;r
zIE��P�&�>*A�]��Sc�L\�M�-r"�!v@�?9+�]�lm��<cx\᧲c�m�"إKǚ����T_�����j�9�"L���Wjf8�C�mL�{0;���::��t�)���o�Vܟ#����^3��O[���<����H�L�$3�o�Q���(���^B��u�_��oܨ,V������B)�5FPj���+G�3�e�i`�B_@�ʦ���[\�d�e �/��F��O<�6x�xTfZ,$�ўr��t��/�=,��T��h��v�!D.��}�U	ڪn��lnmv��� ����]��*��آ���Է��cKѐ�����k�o�yV��HS�S�#Kӈ!.?<=�4�<���Q?毌��61�dÉAKg����Vd��=�M�@R��l;�C$�ѼW<P4����[XʓQ�x�1\���:v%(x���՛�

=*0���C���P:"՟��vA����'`���%�A*�f��;�i�-��@�l��}��.���srK�R��{�f�޼�$��g�,�)0fp5��������U?�/�d�l���P
$t��Cz��z����'*�B�5)���8V�s<�	��� �����QcIȧY�~��g��a���Y��?����\�v~�.f�ti")��njf�(zpj�+��H�l�>�{瘋���%n�o:٬Os��e �z��g$Z�p�.��1����mo�,�#b�j~w8�䑔 �gg?��)�R�^�߀$��$קr�Mˌ�K=h�
�<�kuԛ��T�������đ�h���!���^���Vo�s�KjR���,tG6[��7f/��	�Y���;αo*�C��*�p
���NV� � � �@�+��\������V�~�;�������y&�0�|WA/h2Q����6�A���#'��mGH�1V���y"e���TR�:&���V��?R����-�aV�@@%�+�'��Z}��$��+�V)؄��:�<�vE�*��ĩ&S����ߞ��y����)���O��A�i��p��,��$>BD:$Ƅ�!���]d]N���ti)��Ċ��*Q���-l����W��.sR'xxU�O����#�x�|����Yu� ����)4{��#ґO�_��ׇu+��j&���?TN`uZn���gN	v���^��9�;����u�rV�r/z~lA��\Y����