��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��!���w�9���*�*�)�T��Ym/�3Ɯ��@���<�w��Bk��0C�aYm��\�4��!��y&7�V��=����^���^	�\H��[�s��k�)���l4u�ѐ��u5p�n��Yvn������d����� .�z)�d,��C��n0V/�M��I�)�nl��M��"�³Qg�R�EA�|���!f��l�F]i�ޝܺ.h�w��=AY�R��јQ�[��&2�� �0#Q�T,Ek�>�M��Ϛ�B���q����):��2�S'�{W��l�ժ&%#,BWd�x���t��f��4���w���l�x�j���	O�z��g����������!��L�IB8N�>d)��@Z�B����z������,}j�a�M��]�|��(�z�[w*(k�3n�I�`�z�l[��B�H(�I$���p*	+��ġ՟��-C+�^�(�"�Hގ�]�=��ߒ�ݑ���c"dq;���<)F��/���������vN�Z�G|��!�f���CxU_���jF�őG�n���a��X�06����Z?�m�=��!D|	�J�L�i/��V�����"���7��>y��x/alV�h�?��/�,7����ltd��C��|���_�]b�Mv"͕���23d�K9�9���fjJ?���nWI�����j�nY�\�a�XA�OE�x�b�_�zG`���K��4Y�`�Ӛ-S���mƆ��6	е��j�i�>^��n��L4tD�����='�$���Ꮝ�PL�>�E4"�9���	�a�62�Ui��^���.�Sk�]���/�Ѿ�&잎��F<�9�N�u	��rH�0�콾��Dm���/�%��F.:^L�޹�E �fNo��DJo�䲣eS{ȿ`�9K�~�ax����D)A�+���EL�li�u5�:(I�� �c��e��>^���<_߃t6�l��E��L9��֪�6�����ȱr��o�N��:y6g2{���6�x��7P��{���̧�8z�Pf[�)���0@�O��2F뤪^���t����&�c�F���x���URn3h��������Q�U�{�sP{���(ST <�|�xh�C%���h�����N@N% ����{O������ӫ���i�C��} �-�a��}yeg�	H�(}	XDfA �L�sH�ٓ'\��d������!�x��6�0|¦{y �S�x��yLJ�g\�\���	�{�$�%)A��δ=���Ӹ�'F[sr��R�t��PISP���4�e)������,w/]띾F�H���J%E�+]��SЇv��̽���(�b��=x�pRW���E�$�R��{RT�z����3d*���C���D�,�T����^�u�.������-1>��:"_���'�>�ni��g�դ��>��w������X��}C���F$מ��/�t!�=����J֖�6��J/����-���뜫�/p��P��a��.ㆱ���n�-H�O���V�,or�<�z�6p�t.o�\���@��-��N��Tc� ���G^���LHR�s9���D����յi'��RvS�+��))��d�SG]�)}��OR���,��Eg#�CG��U��3c()� �~[��(8*�������*峁�7H�N�&��KSi*�Fݟ��[8�0k��
�v,ȇO,5���6�����`�V��f�ʏ�
�%茳��B���anγq�^Z-�%�p=л��,JFX�W�ʅ�s���12�垳��.��V���9?�B��ls�r��5��+c9Nhk���PD@H÷��O�JI���~R�@z�����k���o��,�"v�����. 
m��T�z!�B���C�=?��P��Q���!���|2��c�Dh�Z��vy YC��t�Fٟ�'<���C�8�-i��d��24�"���P�ZM�#r��%���/^���7�1��n7��iP/U���Wyx`':a�,X|)�'��<w���e<7e
�.[-�sH�̄�d�<�Mc�E�x�s$����\ �K�~@�j��~�S�'�����]=��g�&[�Tec}>�V`46�����`���>5��^������k:9'J�e��o��^�1�j9�G*�#�{�`v�-��+�d��,�|$�f�"�"7�+ӑ�П�m�b��P���lyW^���N\�ߔh?`i����ݛ���z�O�xҞ.�qrml�k�)�����˸����+<�	e��[o'm �K�X)����e'�����w�B��];'Sn�\����F�M�GCE��;����cB_/w������3t��r��M��R�<����������`���<�I�ǅ�����z��Mq�b|�M����_0�T�X<��`�,���Mx�1g�T�g!����֏����b�I?�>���EīyM��_=Ik`I�3�����^��F����t��Nԭ�k�q]ֳ3�D��ԁ����tC<����Y��'���G��L����6
x��Gf�P賦�q���)��fiR!Ydپ�N*�j� ��[�F25��	�A��J/�^���J����_�gY�*����ʕ~أD�V��B@Cb�l\����^�=WD�u���ˉ� kE,�\�-�����p(�5R*����������hwq��!!]
0��v�����b7�ۈz�$Ta\e�.'>�a�-������6a��W*��փvˡ.����v�n��Z�����D��@��>-٧�B;+���V��0�X��QW���Ề�7V/?�|8�j'�������s���_!�wm?���rmq&�#�I�UP�m�@鍞w���E�:��cSVZg��NT�c
�.S(��s�VN?{�͒�$����f���P�j�C����Zp��;������kƾP�o͋'DyDT��k];�ĔQ��@cM	Y}�� K��ԷsWY�&��ޒ���)� >!mJ�~%{��׼6�^���'��.	=S�B/A%��}
�i9W1�C���X�W�m���0=<c��HY���LtD��k��8�+νX��u�$�����t/Y�v�@e�g�ZVK,��2�Qy�	'�=_����+BI��[�B��1���2��i=X��_A�h='�j��zuM��hbd��,7^�o&≀z_0�[q��gW[#Z�r"?Vى�ɨ�%��g�;��y��~��NE=�|����e rM6�ɼ8t�K)�҃��M�����hj灰�*�ĭ<v1El*ZkJ Ø�F���F�}��/�W^LA���o���x:ۡ�l�M�8����	1⽄^��sl�I?������%��g��Z"ʄ�p7���`�,��؟���ډJx�˥�w���WZ�x�v	x�o�OS�ˌn"�M�r���%�}(��Մ�	&�y: $@Y=LD��f��BJO�|=��n��,�d,E���D�����e���%aǬ���s�-��9<�1�w�Wc������)�&D�u� q?_�PI�k�������Q2��y�K<���USy�LO��[�_Y}�>��ֻ
4n����ʹx��)#���p�̤a�r�X(Ol��Ǖ�à=rг�/B�)0�`
@�7��C����f\>�p�j��Yƅ�hܕ������R\���ٗr OM}+P椷@����(*L�q=�DD�|�!�?r��d��<�1TP��Jg^����?�>���)��\��e«��g�R	s��)`��)Z5xJ�}'I�������*3��y��B7+����"�}�se�:�ƺ���IHo5!��>�9^���%fYCsFnE�f8���5��*y����*���2��e�?Q�����$+�~R��Im����U1���GD�*���b�c�"��#�g�pStx�.��a5���mR�Eآ�#~�Bn�1-D������Z�R�����=�3�:@��&?m��Պ�łł�z/qL�'�k�}���ZC�I"*k�|`t�����oÎK�)�R���I�GG��!p��bJ[�:aҁ�f��fTT��A��ҥ=[mY��&�g/_p��m(sh���U��J-H��;����6�ᝄe3��{m��m�]=��:���Νѕ㑩`5D��0`"-Zu���k5~�q��W���i �zc)Y1l0��{,ݷ�������N$͞��
ֶQ��"�Az��H�c����/s�,$���L�R�q�^7}c5�s�����E궋��z�����^��ۨ��Gr���N�&7)��;k�h������3T��?~T`�kZL��iL2sG�/���ni����<{��矩N����AJ�c��g;4}�"�"y?�LA��'�d*��
�1�a ��r�M�-:�S��<=>�x��G�����˯�d�5�_��Y۶�?._:���-u��@�3�{��\�@k�[�Ǉ)V���-��ԱC,G(�T(�]����JnF�3�g���C��<?G�9�2���;���kL�c�;��/w=L�WM�<�b�&�V��������U��<�o�[`눪W��xm�4=ךب3f1n��LKa�ݦ���wqd
x�������\^�H��C<�;=!�j��"@�v���0w>�5�L(�